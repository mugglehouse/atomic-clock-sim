`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
K9oij6iwk0LonhuF7twf0DuGp+L76FmBC/9C7UhUU+N2r7qm7XFl5m/EC0no7XJPQ/87chhQgjbA
0MGuITxpdQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
HYHioU+pbCrxBDypSA9lW7mrUzWxqvW+sgPR3ujd7VIzQsC5yLYQOutxj191ZKIZVIVlEog/bcZZ
ZbKmBBAvGuS91HPukREQZQezJWAYmg1fggEpFn/0t6ZkcIb39EvccuY2cbsYpOF9fyjlwOMxapKC
SqG0qVKzMZ9WEeLsfw8=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
DyBqzQCDgW+5d+U/pNLGnrPlSQvHQITzM0Y6XI7dQP5X06XNaNWpw3TNJkHF8zyv1iockFW7F2kZ
sfVj0JKR71G6EV7xnZHgxPVV19P+WQQXE+khm4luILFOSxuWwmURf4ZQDzPSZu4R67sTNJ5dVPsL
zw0dxUl4bjZ7qSb0IBE=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z0JSLRkuGgT/ih3a+Yn1sAcBn9Vsez+NlSRFUTTfF2RyepPNDMbSHqNZDv2ESn6+Z457EcOLxq5w
ey7DCdXbxzxPbfxuDcCo0p4iyH7NQL/lTZJpOHari1uYSaJwuLyb6A0SQ5lAAJuMC3EX6WgwhYvh
pMtdot1uTY+3OlkrAYUeAW3x9DhlAUAn6vFEnbZtEK9Gkzd0CVQBFJWGNG24WATtBZRYfqrkdaz6
+t4Rrj2IfxwNBk40g0H1uufcICMXAO+hU3MK7jd1b1o+xLHLzXOhA0mTUwR3KZ+FoaaZPglxokhG
TdNu+JzCf9bSeJvw4hDUe56GnKNQYiNUAa8rqQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Llisuf5pultSHOlycrxYZ6dDEkvfKWSWP++9jqDRdjSN9hmv6RC7jMVwdCZB7TIpsrbuxA0hA+jY
ZgmevTkKMipYtgtHLEntBDRNhJX5tCj634mxJJ0qC+y07mqJMCCsTXbEVys+iAX84CcPvgaJo9Jm
I1iSHeseW155F/QluLM9l8MXO8iVSA/MsZ/kuYq8rQ7AJIh/c0I0UhMgtporD2CY3wX1T6XCYLNp
cD/FTbCeg9lxykLA05IUaSkjDLKdOz/MXO88IvKVyGYalcZXj/lKz7ppWHM78hpNXXQq15WHQbq1
BoFHsA2N0jX9FThrXDs+5Hbq18/JmCcwBbOs0g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TjiasDLWZXRYL3PLLY7HqSRMZ0BlL9b5qZ8zWV6R3sTXjuDClcd6JY+GOhwLQxRMpF5KRWx+FaWH
BJfxpeHuDG8Ktu9ZAfdmakHVtAXEUl/xcilK7cY/Vsa5p1q1f0Dp/GAxrTwVw7UvYJb3c7Bi9JA8
RRsJ/1f/xwLi6QMs1lvUKGXkj/2J1HwNHbyGGUUpTys6y7wk+6Hbi+gPkqdJaOak0Mh4/8JixE4L
WNQtcZnhwK5RN8mFlbZhaCXUPs2rf5dhV2YfwJ+uADOAQIkL1+nh6grVWdqlP7RN2bjuQqBRbpVL
HF2CDQAgdKGkucFrPzMrzsh8BUsLg8ugZhp4Ug==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1558368)
`protect data_block
ImY/brvlwVm/eMpmGJ+FlXLYFnuhJVxbMlXtwfmWCYtQbthWroUWAe1xGmC9xSljjfuCFUey/WC3
O6NDTk/Q2TbWhbP4fI86Mo/26szPGGf4HDGdJhtSWlj0nTZVCBMS2hV4bp3bHEaLdz8g5Vny1NXN
6uQwUqbk8q2c/vmFKbkLOUBFBRSYFNr80uGgPWJqnRMNTCnDRawbKC9PJZhAjmgOlYy9ICN+5RCi
vAIAcIJjhRWTWWDXbI9vY/rFaugX4JJTAduqRmUucfe5EztuBvDXwRfFxf++GrSGvvc1i9qBoPFN
YQ3zx/oz39f0/lvkGIRHWQTCPaD80F6nsynSvzcGjPhhqXNnq2UdECiyOvFx8JtywDOThYu+IYQj
7yW44EylQA62iEXAGeHCdBqhe7nA83NUlf8El4EkIe6J6M6765NCPuWzDIk7dj4Qz5DOrGbqb7Zg
kOhC9AdjEbvPAjTByzfgk6v+XPE+GUw/zE8/Y47hQGZMPhC403iudflLxBQezwPB1TDzQydQe1si
gl59LSNu4DT6tXFJw0NsCsBGtjIfJw+L6/aUhM0VjgGn1XtNZ1OX1JPq9jkT8hxE3tpeY5GpiE0w
/qa/t+NrqyH9gBqADeIrnGjQyQumKdtSs2bp29fwint4EC/+suzsbM0juRIHW90dogYqY/2zYmVm
vgXeQtayQU2W3f3dIxyEn0jynUupyb17mdU99vHQgGuXdnFmO8jTOoRJsPhUP5/aGZ5/Zmjr8EDv
Dpn10GeSc+0o4Z8mTX3/uoCVORYxF8UyOghX4NX58YxEw+t9xmIyQpEjb/dUcWNf1huAynt+8bjf
0HThV96EpQK/Zt4shAU6Rg77xXdccdOAetjiA1A3ms90dYq0pR5jPV0lMCnDJm4fGXEBboIvsQ8y
3UpFPntNOYL/MAP/NvHNSRXj6ESBvl22v0VCDK2Lgnu/17Hw7FUZ+VxEVZLxVxhZKF1kQTGyTTXa
wAGGtyS63qYbYhVzoo6BFtm7KwgoKyUxpJwXFtgHvH4ChzesBPbfz524iJshNHWBi9JkpKjcUkPZ
crNrgSx+wGR4S1N8Ys+ueJqxQKSFkdgp0p9WdCIsrQG/00+8xGi0kIHOmN/GZ6EfNFIq8Prh+Fzx
hX7gMiau+fyMtuQIyD54jp0o3J7jBDGoNNdMAN/eEthSQ4JobSk0vGU9fUCuZxo17QmnQBeir07A
Mn8o40nFxHzUz0caqKLlON+jVLfsXnMkpzw82kKKY9QbN1MUM1+8LG/7Ikb5df8Kwmx4RoQ7GuZX
q9fXa5Lkr6rmrcYnQzKnlIRJEadQ+Hh4GWw3Az7ps/2xriTMZfyyh0YcQKfhdtIm/eAF+lLVUYag
uE38iTcRuzDNHPNO+K3eeNzRWoLOmXD1ovoFhsrRNo422/Anf0icWmh3SHFpdn0eL4ZCYyYXOfMg
BrgPRVIHKj/jb4HY3lpNig6X6i0qUjfb7QXo+6Zn+7UBSgV03+FJXn/x5qqzbvbs5o+MxClinAOq
1bXPEXeTkNiQOqbpd95nOpL903jaC4cAL6oE0dEPMB96U7QgCA/v/Tdz4pZp+LkTXXmkvMQdr7rp
+Ar7H2bKBBFkiW1WFa1kg+BsirhFstC33J4KuJ6j2RTLvJ0URd3BPDck64VxjaDk3wxNLqaK4ASW
E8PhZC6zBcyrMMruF1Hr8qe0Vtih4jtfnRZwMY4urvIO6hFwnACCHFqVnHsfkEPc4Zx5OGm7pIoi
kjyzGJOeexgda1tlTbaaOX9xBtvewot7FR8F3XU/8b6a8CYxLjEID1pFP43m0SovBVlnSTqtabkv
05vH2Tej79VuRgGXCLt4RNGaBPPXeBbjeoep2AG7guWPtqaJv20wqUX9mbSOF7NoP9mmgmTSk5th
vMI2zaP8iIbyvd3g0NJFerahcitgJI95i9t1sAq1XZ6Q+ssHohVybJWEw8fB6fS7aNzQG2wzi6hw
I2aeDMsvlfZvvd9uKgNzPgxlbR7MAO8yVdQ8BfYFzUiibp8e0dfvLzrWVXLWOhrDMI880PdP1UiB
mbdHKC59OEAuMyMMEtYr8WLvyBPxjlFVVlEaOYdHIlrofLr6Ds476pIDJXbs98K//+gztlJGqtF8
tF6+4Fwat7EmD8XMCELaG3DEb9CxeMxwVEqQUKPLbH/LM67IISSSEtr+JHV9AiDXQKaGAvadQ57z
vyEBnOeSq03Dt11PVpvTXNJzw4FbaTTpRE0xBoTUBxua2jq3GZiybANtQcSFQLpd0ES/U+kEJRJ9
eToalo9aW42UdXX2VcSkrU+yMNreKhC4HR3fbCeNAIYe2VgmfNsD2NYNIDHjPw1V94XZpBx7VmRM
HtxA2gvSFmH9z3658fHinnUjpaLkFk7PCGDzXDNg7CwdZDi+EJEz23d8Zhkg1EtyDSLOjn/yGi+V
qXPGIKv7eHFVc+dH8CaRIWa/yHMJ6TaVLzIgQKaq9KTMFuEqAqXsQjUN8Ng4BvFiFL6/J27lhnex
Jfe3ICeWaH7Ujz+g4663nPP/tijI1fwB8eLmF/QS2UCsIEvCKhfDMi5MJAQeQM0XgLs9tOqBzID5
Ct3B0iOsSCNw7oltb+tWP/F0PySNH1lY1retPvRTng0HykwnrMWPDxo10dtDmjf1eDtZi9eP2krG
xlYf6ESUuUIZ2KSfX/zX+B1c0bxobs8JxAvTlFXIrS+zAPJCbDc+WL9Fk8UY/Fv1KkyQk69Bg5U+
dBOt8J+sSTP9CyJTb2xPt6AqEuUwbfiGKA2H7o/GL7HA0RDmi0i5ieEzqGbYfPC6Fdpf4MlZA2DF
WbAD9caGhBnuOaSEtYzn/fE+mQIgTCrdHVEB9gPi1GemYy19WvY4gJlQYdFYcItkaeK8vCt2uqeA
e0eU56aM+TT8HTrdpv9gviaXtEUQ65P9ogqp4BLsT/DUKHapJpvRAsfF/YLCz0pT5QlGGzsPxBy4
1SLr55zIt0oaO2PL/mtz6Hlg2uGGQbrSbDg3HJPEdPmHvsfLYBKcP46ZkpDq2ZfrOmN0x/FQ1mMu
UvYro+i7xY2TFjAtAKNeyfXSJDtgXZSegI33eyVaJurIVVqP1qRBMeXOFSROypncM+R85hh1d/9j
JBVBdtqK/YjzGxBSWRad7Uv96yoTb9EX5nMY1zDN287kszysSkOHJySxjKb5vdr/6YVISwWGZVwP
sVWYUm0OgvUtObwl4B0mZxacFdkN1HJ4sI/BCTuxpn3y0H/6ZZVVoQ66Zf8QEo9DUazPbWYvKRzq
0VzCTq9TZZuhcGfOglp7btJkREdajzczB5xj8zDtEznaLCcCPbv8J8VdkdJwsd7A4P5IEF9lINXb
x3+hSerbuRozKQ86OSWEAKmtW/+MR8xsndDWcqbtC39Y92dqgpD+1Uwh6iZLVLrs7K5q8H0FwuhZ
FunCAC4donGI1vEEMKAwq5pQMwQionFre8vHgYorzlvpPPb6AgjoIyuaMhcwgKZbnwhbqw3DeqNZ
UUP74fWtmU22jgJsnzS3bR4OSEXg9a6QoF+odK0Baw1wyF5ahf/RiPD4dfLSxXLrIkOrQOHyGBfn
5FUZm+RYkM4Uei1jMcpb9/I5cJ0D7AyWNz43XsWagAXHweWi5umdIlXwyX8Efx/TP/Vm5JOu04AN
9E3An0i7ThU+7sCfwdAILzcZdZkyMQODH4ZjDp+d8yG0Ps0G1fKxQ09blbW74NwRxjt8GjwH1Ejy
fdwyJHZaxF+Jdeu5T3NoraMHNM5Dk7Dgppk57Wx/SfT02AbFtisx3kNUfOxsMSaml7YLzjYhMj0v
GkWtTydBv/LDN7kzU1hEVJiaGtPvUGl0HVGchSsEOvQxciavRrUlA/IDrivL2kzfRg/E1EEHQ/jl
JAKe4/HIeHYNKIsPkkgVo3iLp6/RtllC0ET7Rwmy4fstUzdRblDCT29K4qQmFFc26K4mZ2KtiwGH
Ugk4FmTkDVQSDmPnXYOnMiHoLIf8QoZUTna3SOQFzcmIV764k9aXb24feBLMvj1zLEQyCohxn0MF
T/gNMU0Ye3n5Tn3WhCvB6PsuSvB3Skr/fm53etLV3hRKxKP8Vrr3f7mWzK8cGKioUN3Iug9XdU5p
Bd/1LYIpEvOxJJiS7rtZHmi38lytJMbHOCLSExJ20WWZ7rZxKrujvPsuBecGEnAk3bqfDcvTVoXq
eXRTv2eItnlaXUvpLSNJ7stV88PDsjPHIfPZnABQiQwssFaZ6u9R1XItxeqwQBuemduOMZCeuqKQ
zMu8uTgVGs2wBHdKdQ32Ygbw6zu4C2poWEQ2v3Oh5OiqauiOs6K9HWmdpiaD9xEWUZyfBzFJ+qUB
Q6evjluWuuj0O7TzeroAINgXusQEu9GddiDm2sWuvNXiUNEKwfurWCRb3vYO3Z9xNaD5iasiolrA
Uc13uN9fWvF8q4waq5GJdFpWQGY7fFu1vgpL0hOuyaOBw3H+E/QWNdMudu+gtZoCoxHizQdmP0TR
iVY+GIdYxrHDjcSyr25oj4pFfWIVmQVHk7eD0dJrmD4UWQpvObJz+GQY08CKolcpNewmU0Emi1FA
lDGluZSaoY0Lu8ZuBFQIXpPnJswbw9CZkmCpIhpSclXbTIuzQyFcC18Kzqz9DXItuD+fiMOa6NDf
P01euoA7A2g97plOx+9HJbCRCfkQkhLlRgytb5aVF++URb60qi/uR672Zo1hpgGSh777PqE0i4r5
60oghljNkXr/KSUEIHsxZkC8iG7EfVtOSnm8sgBEg8Ul66ZiDetbjCCE4MyudqQjWjpyXc+hvoCw
oWMso+EdDXG6cAU1a54gIbmpJ5wTwXeieYY8U1JLBncyiNwz7ScFlMWXouuAWHmhI0qW4cJIgJ+k
XLvHYAHOB0ju+w1YOqZ0+ljkjuitSE1YSIZe6V9Gl65JPyRWKpKhvGo48JyeaHOu0m4SL3IXS7dq
vvwvSbieEKORYHSEF7DC9l1OYN19p7uD+dolEDOEfEMJoQlHqQC1RFMbmScPBCKdNXKoAdSuCldM
tsZBrldqfN4Hq5m30UlpcmpNvl22zWEypOHGADxrqaHdvdHtA7II4SnBpnOIB0xZJIscwh9AdRvQ
Yw+DKpXSviOZSXZY7yqjLm2dh3MN43YznqMM7w1UemyOq/GvKHUZCTBaPVT9MmhyC8+9qJXHUxm2
RTa2xhH0ZjjcPhXgIvPjxxKTIQffrdIVOW38SKDz8V7lpywICs1/MgTdHY3Nmwe6BO0lKHc2r+c3
hipGuv438YJJnBZ4nLrJy01cB79zxhsyJKJm60EFr0qV3RMTEibJFoTYQmcLgy3Ie2iT/J9/kqXT
4+4lrtzrktD6BMVAvXnvndK8pFVHMtcP/Ho3bpz3IIztQe0ZaiO24QKKefTII0LCyOzpAe+h0kmy
OoayOwn6FoCd2JGYIq31VB7odp8S7waWTtCKGJ5rXaSjdxiljz66YsYr10cu8gFegcsjXEJAcNdM
lYxdsrLg5YcUGzemeodS0wklx35nVq0wRPh8koUspBC5uOcHyk2S55xVHOkVndQk+dL2qMwV63KL
lS8dF23NE0+Sk+PHrnf5Tl/NBqsvYzib7nHAUCYh39lSRpN3CJUTgv4t6uOqhxsTgsLozRmmBnzh
qwWFR3MFA51cn0z2JPQV+8mhTfW6VmmwHpEOZ5fAMgcUZFvSrpqy5adqB+UrVRbyqIK/HX2NyvE8
zS/V2aNKHZMzlwyqK1I45tqSm7NrFbyma6Jxy0JwO/pEhT1lnkVdSD6rbRbNCP5CCKX0RMP4Hng5
d8cSY7LF2bhYvtjNOXQOjBnxIoixT6UC3YAOaXOsMNm/MaF8J69LFQOPs06RmKrugwbzaJSSM9S5
tGiL0xFAGRJIaPrWIUHEb+6D4Ww6QNdDVP58NxZ7YRV+QJSicjDza+sgkDPFa7c7b6TqnSymtOLA
6DsuwbJVdN+znv0ZvVhun9vRZT/zlRM76uiYE8W6B88kF6iTmg8/oBEqJZK4AGbsmJdE18csxzG4
lpuwCDW294x9pOHItrmrvKkL9e4wH1PlZ8paEwhuW5oxAJ6CFMtczMxj0rCiHkESQFgHSJDWp4M6
90bqj+sBqyjPBHm+1x1ytuiW/WYLsS6y3WSqpZgmVNJBjf4hb8hqyjvMhrJrHFbIAhAo6rKWtSge
zXGPvcdD6scanNwfo481USeEJUi5k2k876dQWFTGqChr6z0e2eWbMKCpxIX7525xzArC39tlKODF
W2qap86hKW+1E5u8x82OJrz0En8pFBSGHPnnp1/ihtoE7p1IF03A9AEpnVXE90CjQ0f9+MOv6kZw
b9FSgxZXMmuwk9zamFBvpr3eVTV4sfh+ACJg2Veob1DqqIrfZ4WroNN7qLYy0jWbXrQOOPiExPsb
X9yDMxtp5RjqmVzOCWZzrgFPj7uaxkwUuppfcm5R5Rmb2TTDHRWBzUAXBm6r4oovtJuARuNrtB4W
ibL85Fq+/rQBFs2+jDYIPlzEZX4Vs57Ra4YiprBfD5lw3z1K76FrF3Jmfr56bh3i9gfE5lOYtkF4
tQUFhLVZSEevW0R7dJ8itwisSlWyv+9TfO2H08s+o8QUEpWwfVSDl621wSbBX8rO4AjIiMuzvnLH
GzLkOjhcVKj5qXJxgT/FzVH6+Zy8TRUB/VVGmDjuFxrlgoWQJXZnbEqICutRKzIk/ftrOtexavhG
qlUWii67vQMsqFrEyTDuhQXncsr3FvaZKMxMA+WsapKnscaYWevryyUe6k1xqvwtFGitONdhGQb/
otb+ic6JipGd4nz0RfKLiTFgiI1NmL5ajbRAd3ypHMHTLbNkvlSeeMnl+HnJPWOKBCTQdUKEu6Ct
I8ni7wohjKKyGNUiulu6VlJ8VrUkJPRIGxv8523ZS4seB9XHRsn0exWOtriao9i5xQQRQHnj1Z4v
tT/mkgU6pcKFO/5x6KPN3BPCpghC1UumdUKuMyEFeh9ndlr4xzwuX7Bcs0nurrBq6ipuE/xNka3A
u9AjNCjqMfIjPvgFOydgetnTWZSpD+j6xk62N+/FO1Mcuxg46rQVIkdvbpMjkykMqd6RHPlekBs+
y3RUbXBB0tSQDSOKVUAvvTj9ogD5TGVfy4Qoz+LLFyxWfOlbJav11kutepIziffRrSwws/I+fOQJ
LQ9CGWdwa0gU9SqnZt2GfXcZB+ca2uwHb2U6u4VDBdGX9+FYnIykyIYQHC/H1uAJf/OY3UUNzO4W
ILEZoDwqYMBEqTPi0b8SOrXidKXqDFJ8275x2wF4fjkN7aaNk2Q4pKxw5W5Ry/XgW/zOKAWyWOG7
ywnF1vXEEaKD5MOEwx0iT26YQO25y2TYPY4p5RDxGh6S13W1aMCi4zif3ERpbaUiCUvlizXYXeko
iE58FBz7pOR0ztrpmjO5LTxVv5ScSdFmj3w/wvixO6lkRPNe7KyuxqKczWBrbrJ/l2f6xFT2Vl1k
RKZSPNZhEqMULAUpo0LF/6RHTtQTMpTewdnZDXcmb9fzo0zUp+qFS9sCDepfdmtRGF7BN58iS5DH
zNHxl6jni9EHUTv6nSWjB9orTJvxq1//PF9rKb2F+Txjun6MGqg1GiE3fI0dKssJKpImWDsJ4K3M
2KQdVT3ZVqM4LjlhsvcM1mf0MEAWtRZ+2GpmsLL2CTEhmfkn9roeRzscxaiXLyV2nPYjpZWvJbVy
mPwIAQQCnk2OUuvmwD4q2BJM/5UzLqLLLSWCj0JglAr3EDym5mC/bKjD1qVZu3SznMxTDaLd770t
JeOSx/B8f49qxXQbbF3Eu0Qeh9OqeabBG+sliw8k5xkw/E8xTulVCZJEfI+Jf6GCo8GL/P0bgjfa
YxTi4Gk3FypkkjuBIjH/sHyOCDmwFwPjBGGYsLHLHgnrgN1WHhO+cXqBofdSXlEso5LhLA0oCiOU
FyN953gYwzy1+GpU1LzQMCLLYZ7cxUFVseousvLvPllR0oKbFOEHwH9sJQKLOMXVS3om8lKmJqX7
+UdH3p4CxhrtRqzeKsvVh85feIx7OC8nf8o0rh9Pm4EUdTSMZNfdlXcCSOzlIdkB3+OHJWv1Y+za
9lIc/J+3L0w1svoPf5yW/MzT7IodUF8toWq1UKS2V9B4S230Y98IqI0B0m8GZDnyxT+lbLIyzcMh
wcIY3OHQGl4nr3Kc9gfpLI6D7zGplYiVTfVSrV/IjopXnsZcTDdkYnJ75GmaLI0Cl9NBNyMSuCo2
SpDEtBs7+MetAaOe7SLzTG3N3NRDF2YllPu5Sx6uCAWueJdMdNN3y+/eAp9ni7mRCvBdOy//aU6c
OGtzUhhiOTWIkGZcwMLXw90f9hTgJEdLOxEf5zsDUb60j78bR0s/dzKGg0Dfwscisc588Ct0PuB+
rfaPTfcerO/G/BVd8Fuc8JSpHGi/RPkvyVRt2ItlvWbdOBNW9LZg8dNHkR0xmLRgtdsjmew+Jsdc
wyoo5PT6tNzsJ0oP7T1quKUdbFr3qiE6gX1Ncr9kpaDhRJLlJbPbO2ApheP7Uj+ZSHCGpsfCNPL7
JcifYxWzH+Uyt7l/MX6GscWYagcjFQLgslaitvgOKaBeU4rHrNBEKvGQEMF3bx2DsExNwSlOZPZz
qrGdJ4DV3weCRndRu8g8G9Yv7T+25taZHh175PUgRpbAI1no0pH0mXMgY9s5pm4Fknkzdm3/PZ1e
ySLo/wYvTPiOvv2kK9LfNgq1tB7AlrvMlZvGGd+KVxI3LssnOa7BybjaPLXx9xztNL9YANgbHAaG
EaCElBUa/aB23w/MugkFrP1wzCxilGh1MQdx4AD/fFLx7sOjarqfNgCzifW8fdLURCBld/e7ZSRS
JdkJxjhRxY6619dVI8dlS/2icV4n5EAg/9xHtlATBLWz4V+16eIocg4AGd1ynv9tcgZXvzQClCyS
MDqKItF5JDOAc3KruBQjly3ilsm3gqIn64SYrqRAvfMVneyEsNalTB6SB8IVgbvv4oK7/51e1xAP
vt6LU692GmNonFQJbfA7V8WkPVSsTTjYqAqqVoqQaaFMDkCo7EzFUtdofVSFfegSNm+QPKmFdmgK
B/cJpCCzo88ieLOSRkyhF0PF+zBZYSh5svoi7GRgFyvd9MK9ZlYi7h1Ws/UIEjEXDdzWmtyujPXo
hlIrQZb+yWoaFLPPAh/GxZlYMV+/KM9MhdSc9HEczgUFnR0F2pb0VG6U+6Qqh+y149GoQAPE7V7O
OSD0+qNKXkgsOC+CHgMsQ2PIOm6x3dX4t+DQk5YXWwLtBt+5g8Jb5Z480C155rm+HSjsTbNU21WH
JibcuEQhxX9tui2HOsVW3frRUpkamgUhF0s+3XYJdRDjF4JQzKVNrz0skE6leXcYCwUr+WQCmrDA
anrXlw3rixwMiUMuceVl/h7WbYmuwWz/FqsT7eWbBaSIxND+cGEkaPwy0R+ISuVg2Yssp16JWmAG
EGQddvMjnao84BoFwltKwOlmkPw73+gkwN9D1sktj2tyhgaPol4VnXNTyzU0+zNShDLulhU1IXoC
TK7i2tXufNiNV1BJX39s6kcILCqFGNpG+9zAyBAT+pqSnAz9bQ4p14iLjpp/vq1V4TZOLOt6u9/u
/Jq1Qb9yW+BU74we5JIIa1BzZu8KBHraadHInktOenprIs3ang+OW7lUXuTvfdKhIsj2YF8p2VF9
3I8qulPdM8pu5OBWeOL7J9KvUOOssSkGvjUznnbmXZs3y6OQZEjJJ1LmTmtNqY05oGLulCD7J7EJ
qaTqExJDJLuPidcbASBcDalXe8cBO19GZvWcpOf1WgKSuu5N7eKe5gFIIIWtsgpfjyDwKFPhX6Sc
rDCcMi3ZRCdIoJCG5PSw033S+OZVVnQQ0ezomdqiqGKc4v8VWCo5FJl8KYQtMwEng6fGE71OiDgK
jCd68ls62MV+AMPVTrfHJppb2iPiCsNbbq/dH3kkr7D1ZKotPQ0I//Eo8d6VWag19OwuMFZI37f6
ExjdOnPhQ90ph0GCSdVIITWah9FBDkrAFqfM10idVE1iPDSMicu2GJ7k74iVfI67ByrWdR2pmggN
YXk/JOLT5bS7x8UAWaM4YUfCytL9NS+RDS3N+f+QdhnistCC4dKzvgNie7N6PomDO7qBin/RBAXG
F/npdltMf/6DALuRAGmstlwn2HgBETLAZ7couc7msUwNgFJQqAt+aUfx9E7kg5KX1BeSXX18bZZK
LEEvQAgnLcnlxMsU5cQlviFeL/uwXobo1sHkWbQ2q/96MJiNUnVulcdtl83EwImyntTl2TrTgnN5
9i7IhDq5MZebMthmQXab2dmykQmMu6TCJCgY4g4sF00BS6TmLXH86QrIygn1b4r4sAvBNkJBpz8i
s2w6nbfumHBN/BaEtw6oEn5blYa4r5an4YjWxieAc7TUa+FqrCYIEKReZfrXqYt3vTkxmwSB2ByO
QA2wXYvbqMOZNLoo15w5PjCftj5f5ZfzBjUWLb085Drj+Mc76EcqxyX2+3AFjHkn5z3uKbUx1DmD
sF+LFbCJKFze/befxr7n9t13n8f+VWvNiVmCLjfIwd2ssdDKmKM3Th8pJRoxo3bGEY80CKBMi4R/
2/7A3RClwrPEtrDjeINHLdABzv+YFMYX14b62Fj/hFoyocbkOVnF5C4FoLOnNlguo7FbQCje1dXn
UoGOqnKcLVKR1cwcE6DC4RYkVoChLKS3i/gYdQMXscOv78IJ2WsaQIx694uk+B+m5AdeDNpBwaus
zM0HP01kH5SC2cHKNAvbB3N4g5baszq7uzsK1B5NiVI+inBqwidjUMvK1ovVXAobPWj+bgIfkTg8
3Q0FtWsTaziVsVrj2AGCTCxhUA1VLQ5l7ouCczypthFPR3hXynxRkNBq927IykmVqX9IlVmiGkGD
BCMddlkZu2eAQ+OVSqLscGoJF4wEozT3k4mxx4bZIrNSBUDPo9+04XxSMEId36gd4EyOYVvB3Eui
6ShS6qRXXhE4cvfo58A4klhk5veYKgD8LJK8PBUphDUF2N1ZdsQwuNsMfdP4OCA205ldGfCrlxJp
hFm7W3Tho00tWJRSC9bn6uGO4l+BoSi1Rx5b3QD988BdfQdclGSlwp1xrQq1qXfQnDKFDQ2mcpIg
PGdaPg3jCysq2zB7bmyjwc23RWf8t0KYe/rPbRaqfwGBXLh8l45an3qd3X8SJrhsTuxaptNmAkMe
EWLA/R0ciZjy2xlYl/ILSnne8x6TtxuGEB6/5V1hIOgviTtKWzJrEGs75/ZAq85bKdY12J0OMGoN
EW17F57O2pfIgoBi/U16mNGvJup3f/KZ8WczPPYsf4Pu4LovBKBWx16GEg9rZ4cGmtwtw1RJJmci
RIOsrIgJREE5zUmo+tZfMutBnY46/bW5qpaFNmQUqkjhBHT41IGsvvSajYmbBGxV8GHRgciqKyxc
DCSKqSqPq+kzeWyNVX9hLtoYBnqJNxDCV999vW7Ss+ZJLeR0MnT24iUPBsK3VLmtO+hNhby/yvA9
p/C6YiayXsMApl0inMrIbcTSzqUTe+HHmHf4sD5B0/fDcFcaGcl9uZ5+Vk6RgHLbas9mlPUVvlSW
VD+t6+cQ2W0TKKupaTViUbc39al1lWmIdhil6pQ1EVBA5AUUiSLNO4AzXZT004L6nbjkQaUCQ/k9
brId75oUDI2QLdKoic3ol4isTWcwHfFtrIButl7KH31vdZXYDHq6zieh30ZwfwVBM+PJJAX036qY
L7z7IvhCs9kO844u61SO0Zf7N7wdYRCt0/AmmRpkmsbFIIxNvw7PrK53cCoECGvWexiy9xuCQWTR
5mKgyRTcYdKnx91YwZAId+iMWnOWyxc+KA4kU3Wa9Tfv5deW+lifdCYRzYZFCuLR1B2upQ0TKEKW
y6MtmmlArIgIouuAr0L9V2LkbNzSzBK1y6rUzqPbb75IcSuokDtX9McViPciK4Q3J7V4HD4mEYHm
0oGsYqZRBvwIQMdi3IMUqtT56SvlF04pbpnONSMFqNM3bZs9uWm1pm5rsgXggedy6fXxCuw9QW8+
Fk3rBB/R9clQXxiErg7tEiQm/Xj84V2IoXV0VBI8s3fIXWsAydqT7jWXOVMg4wFGQmYTEeL0h7gH
L0hjzuwOS2dH84qfL0SpPwqE5IHyS2CrNDUG6V1JlINB7Alo3Q/SQW89AdyltiWtBLT1jgF9l6Fu
OpIAN8CVLSf+3r86vycsmUeeUzKzdyB6Pl6ZKWEZI+rtGw+UcIhgsbG6r+PrctOyvdbXV/oKv3lp
3714ozryOhkvCD7jIDr57ICMEXeXGLEN7onOJPPHn3eCCy9jtnKNHHVz5TTWp7y8jdGnMukBXMbe
HaiKdSdrkIpwI3+GBprpiIYKsz3Vvmo4jJ+t1g2zxIpfuqfm+0ux3InGbY7FVUirxbLm5vsRA07S
Rs27w8isk0/rNmV8z7BKwEWk4HLkDEFwODnQLT4MnrG1SI3erXQXgZEFewTg1EiqSMz1c95Lq//q
j9RgVT8WQqFIgySzVnXFfdXmSea+ZcPTUL7cl6LSGNuEAM6EeZqktQXT78+bTFpY40RJ+b/GdQm1
A/k1nVeB3mqiie3lF3UUmEcMNLgZTLYUjCD4JhXF+b//L7VwUpKHOQTSOiXvDO1sXdoaEeIHPJA9
TqzlRoJvlfhN/sKpx0UnpT5OlPXYyVd2s1U3JBwKoOUStNrNrzB5QnM4vpfaXyvubs9Q7ON7NNQB
DFnMPgMdG+XTcdi5Huy9eGumoc3YCB+BSqWHL8/fQQpTXUsBLlUl/236YgzVHT1efFHChX8iaQNo
/TOSH+lyO4uPmB8Ay1Jd+IXGkV1Gt3+zmszrkGSmSqRD4bNCciM2yBBIR5uD8huBTeBTQGCpkuBR
6Fo3/VUrdK65Wpwxon0krZhT/lmpv5CwgR5SC/7a3gEVPavuiovJ2iQTAlt6yhmNTa19BAryCy5C
IXtNGedMkEbWs8Agb1JKcaZnqSzvJNR/uv4s2cIPCyaq9rcWYEVspQX3jpqWuJKs1nruHrVVa/os
FWqxvILO3A5ZBvXtaSrJ41egnlWFbDfGKJvzEKYtZKO0M2P9rtcjIAZAMKXjOn8gpQmhUIZBlbFy
f/jDywsngx+5CzRdmo/v7reoEaAsLLaP3ureSt1wlk9mbNW/Ro73tVOgPtsExDiKwZM8fHM5N89o
vkM99LZkewfojc2iH3HYAqhXB/vAsidz60X3totlAmP/bTJd+hJT7uNwBFDsmAlZwRMGTvdI19Sc
qEwrI4NKdv6sqV9Ied8SfnNQgOclRZTR7Yje8cUX/Dx9KPpvOSZ9ZpTA7+bGVc64UO3hkFjqifgB
/EMeySNpRByhU0DhSksZHpKe5PLO3fd9qNGT9r+VFYhRekUSgFKqq2yQ1GvdCYDXBj5z13Ck13pD
Xnz1zy04qp5/8ZqLCywse2+LVnuoYlU7AaW1xxiRqQObyzShUNIQeS0YsawItuzCTHsXxneWyIuY
Gl/HgcN5phs+V7Pye48fEod19TZzq8joW2UiIPZjSR6/a7cEJ+mNGEEdJToutVpf19MXVwLLgY8/
h1nqK4lsgkPxaWF44QF/ZYAzJ46xXnLGgHWN3mIHFmRHDGw3fHLrD87/uvrYRNOsqRTd1IHSH+9O
+w9kLsTEqjwB8C5BmQEXsyoSdSOBdVPp7rwxs4OcSO/iHcBOIcfbg6TLc/6fw+9Px+jZyjszkufo
rbdVlM6SS0JdqBKsRb3aN9W3RjODAA+j2plBg3oruXuJTKoV+M2r8GpFSblt8jgw7DssdcUb9Yeq
YMkofAE/V2qh/5FQoT+EsXwm0GyXSfQ7r4WlCc5TSWE85UpX5Clw6Djq2iWhjH8xjhHOAj6ZJmov
MHv3YttQtw+86L4NVmuCzB25n91rC0wLCQtjVm6qZ7rIwOBaJ6y0P3vcZZcYKwP2TI7pJm3bf8ex
r5PVdAMVHOw/zyQSZQl60kDZn4zmKXrX+dEgWmaBpOn4jdJeV5qfuyz9Dl2USS8VldVIN6QBsQuF
9SdxMvEO/Y1pZP2kfjzRcI+pSmvL10ZKp31dvOu/8cjzwHRkvgXVqrEz5Ch6zu1+hVdtZPIQikwy
5LiQYEzCSCN4p2Jcp7hjsjGuJlXkBZ3lFSC+ArSzK3lZDpAK9wybcyopqgSyKzL980Vo7fX8jn4U
qFKdQNAPPVqhFAJvM1tBm2updtMSNHYYBSE38oJIVBk90zPMkyFcCfJ4gt0ITkjAw+zxFh1pOL71
fbGP0p/DxCor2K7QqYm7rDusM4SdeGESRzumG/Qq0J3lG0ad6aNxcLfZ2xKkgZ+brLr1CWZOVKi0
s/zO6nYnBYaI9IgLl+0JgsP/KSkXwR7blQtkJCGlcH2nUOFpwv+ljcX6tIdR+p8oPOB2PnW9H8m0
v0b2iG430TZcRdQoAZUAhVd04Ar+CnEMJzaEX4CyU1vxQSiTgHJcpEycQg2d8kWxBSwMJ5QAcJEr
wMrLqBu0o8DoEpGEO6UuQhjxLe0OcsPcMutpx+yBvMoNgr7TUnfH5lLkMCcrjJy2XuvRonVhyzgG
Xk+3bAMDPK++NuVZPt9Abr58WElaGroG4a4bgDvyKLtQ5yQN/oIvpE9SNBUnfBSfxXl8lrkq6g30
5e5QEBEBIrdXnQARwg6br+MZITwdsneilS3ieIunse+joHmmOx35npRTGtYhbShQ9nIABO1T14Ks
P3HmP3QWuWIDtss0Kp+JjZImG07nkhAR0gy+0BXxx0LhUzrtbk+i0lav6ElCID+mhWSjNWfqvIxP
5tlM1CqZOLpTD/5YOz3vBg2aaJFnOJ2bRaNsM8Vay0m1Lmut3cce9fr9c1KCiZP5Pv+SaP+YIG1b
+yuUGEJXvdLtTzeYnhU+zby/1h4Z87wJ/ukEBg2ng8oZHsmyFg9LW2ndSLka9ce0BYj/ruA+A5PE
my1fIfYFw+21KYQLDJurov40WvSIaEdOKnnvOUO2/axxtBSzT7SOzVbueiZljqvEuq66YXQOIi/O
imSzd9A21E41h1xETStQ//9zaEFQsmF59UGWQGyxJROL6QP6VYNBb3Zy3LmKRMRDe1uR/cKDMZ/h
JKS4/GptJE2YvLjPAGLOqWEy5XxPfFqzoHTrJ1wLA6z2CjD4p0L8LhXpQiA+/cVT7Cw9hw+HAVQI
7boecbHTf5LEX2dmJ4MHQwYtNY47qFpvvUYBRVteC1a4ihub0b+TXlm39CJ80g1VO6YSQi2WoZfe
JeiMMegX86HP1eb6VK58JwXx1YvP+jQ3SOXh/nGNzlNcVWb1vFfrwVDFEN5fhWDCik2p8DNyp/TF
yOJZDH4Rn5cvFbbuHI/rdp7Lc2LIcZN37jGWHZ/MmEN3mzgOyeZPSuoLLEankDlnHwyD9iQc5kb2
I2Ex8U+dDByFyiAAeeXS1PYU0+2O66za7tzr2bmsSW0PHIE6lvESI2VbAyNXMpcBSkgftiDH2x1w
ac4rMFQUTZ4PTbQJkpbgof3fHzjGBBm0kKVtB+W8sxoHyjZESYVPdfbEqMYJueiNnp5dRoA53buI
thq2/zSmL+ZEpGno4Xf4IDunOHHVvvB5Td6cDV8HEuhqbJMDLPriBsuLKlXahPWsdyIgzP/syibE
pgozYhg6RwGdMntoku9hqhJUz67YYB4QTGWsMwDqsvqAEle+EI519Q5YfqpPO1VZYsEzNCNhVaf0
hE6J2nLq2UhxlH2B+R7DHfUSSiY5aWJFhX9t8X9HIhdKcNeYSk9JtWxLAWVmekut5wpsNiGiDgcZ
qZrHZd1PROEPbg52g/ouez1O1hToQ85OfMrQc67YXm3QS4Uda7DI+FxjSXG5ihvn8D8Ptrzqalyy
nwK/xvvoh+NCJqvzbOHbUNw7kcxxxfT4MZjBAUAx6LrzA0rlGc69ye2Amrv74gy8//GeYXINDNor
MVpu4+PQc5dxo/6nw0GILiM3tuMqeQM2sWk/9xyIWTl3CFnjjx+wE5MYNGPYvSYVqm4hO9TyHJDH
laMgFHHn8TsTcREhcWDsIM/oe8QHZiTKPdt81VbFuEUZ9tjUC0bTtsRrsP5Gu168/+lRKJRSg/Ss
E4yqFDdzehUbqWW+Bbk8Wgd+eyTAOoBwtJAYeuT+efu/3OpZ49B6Co+6F0auhBU9xa1NgZFnvE2I
zsvTAqWk/JlmRwC5vpT/m+iw+p/yVTbCJUlxXodbJDzMC1xBh+pavWAW27vrz/YaWcksx/6tGCtc
1NSOgJsXp6BErdTtuSi9AO+HQpQt9m7BI8F76vQ2u+lmguFSD3RU5u2hEgx9Au/DqvpLxsNWtHkW
yeJdtk5DcuEAyqFV2IdJUmMFp73JXE7Qn4WEdyzBSOpXAWeptoJgcIPdCwvHkvL3TPo/roPzbCwB
bFtthQR5FhovOZThDYsp5OfSNHWiQkMnbmp3EhROcBDsd11es7c9ikvdpF2KXGfcyuQIzV/2dVo2
Gxmgz9afUB+VtUevlcv7hhtZcYa/WOJOElwYTYuMOJPqhG10PqWR7zI/NMbM++krvJEO/lFQlWc7
D9QhY43sjRtmvMvgItlP85woirA28Cbuol9h/tAWD1/SY3MIxENpOtowvIajlC2B7XkmfXeTrjm8
MYiYDU7LSYeujYFSpTOMnKdfuKd1sRhzdKdi0SR00MQDUsTCG52+QbVvNF9PWtwnbbB+SREGbcED
zobcfQkVRrEwq3miZY69dbmjFCl16w2JwIxI/P2si9vJzo5z8D+JqcRaYDA1xvkXxkzcDbLldZLD
poIA+g6CYHbxu0y1Zv969j1o/lB4kcXf5/wMj6vjUQSCflXXmDz6sdAIh0KXCtyCeRZeYj+jnU78
hq3qjiTFSIXmscgg3G5/+2zPrp4xOA6voolXTLyLJkPYM9/B9QKkXyOXmHJy7rxDp9uzrdDQfDHw
+t6lW4kAjeo0QsuQU0gfurWJTXdVacLQ19TcxVBXXRZQcBzEnxEmTNJTQgYwAuUvsghGEshIB3KP
peDlctPcDmuDSSFSnfbX/RwONxQjRkW/WRK+WLa6CVrji/fo2csqvHELKE79szkYveq8mNdN8m+l
vI8ELel1GZWoip/2E8LO+jSgsNIvHklqc6nG6bsR7Nc2BX+l6BlLuKx1wtmR+GNQkThp5siYW11I
4g7YMA2jJa2xfuFxBwDfKAnRkbSH8sr5DGGwWYP6/s0WyU6MMa71Kvv70FZhPqRcq3rZCdawgNl3
GexctM9irPq0pKlKiUe5BWpa00cPam/P1vGOrlVhcmX4ki7LUp7cICxg6bksYtbkCfXbVKGrTIo5
bv/nPSmWVaMaclVNvye4ThcnONOp0/4tEMP+pf67CLkzQAS0f0NBSFCQD+xVL8mWfTDLuJrFVzZU
+52jAZdK0wYC0GhDfGXmailKO/aXTYczOfhoNRlYuxZZogx3mxKY9aDwdZTtyQiCt39A3E092pHN
ApH18bqD8l6TZB/QBanGcTYeQ3B60v6n8GxRYk995vovtAFk7nj6BTzfRqY9VPukO0UqnEkfuNMN
KiWfQltcMMP0T64OBo7aaWBfUO1oSJXjK7co0b4QiYEJTUqyX+tuBJ/O9LlaCsyxVuUcM3yHwLHY
7DTlnm/orDu6a3NZgM9YPsHTuf7YRXpYEq/wDv7cmf8ypFmakrFGMzZc4Gn7sIqpNoap43NKUmq9
h7VNxeX8Xwl3vgc5fkI656QmGkAfKwRyiz4KENKOrNClWcta1rgW/thdugSE1oPY8ZcU3pnFxkrH
/2Fw26VvF/QajuXtRwAVufJahXQf9dNjzhzaItAiwdDCTjx35HympbM7oEntNEcnaeQGLqVUfZfi
JoN6X3lXBn43tyZMZjisofw5ijviEAlKTPblQ9/xc/C+Z5ZQ+bBawups3skCuZkzdRiG2P25McFX
eVrsKtHXokhXYTN5Uv7KZDZP73l6AVp1j4RDu9DPdqk1Ymnw30F+21OabZTHiAsI3LF+yG9ADM3n
K0R1aqKxjXVYuGU+I0L8reORfC9kDhV7GmCCApmKQOwigYo2fLJ4PpYROheZhmk/dz1CM8OGpn4M
toSCVyWgKFTauf3fZkZoNknd2YxNfqgqOb9QR/IIYTJ8Y5FIRYEsOsSTSBAnh9ZNzx+1APE28ehJ
eZryuOb8TBFoH5oLxTXz7t9Uz30up24FUPtGhmj4CFjxWHBGQQh+DooHuS8Kpmr+0DUm6Kdk/Z7G
Ve+8w/OmddChDmzNx5trSR4cPWF/VPDBFUb9Aa+6w5jHZSq4DnRVq3boWcYjABJ+vLA7k93crcGi
cw/iHHyxfp4nf8KwAf5DXFxZko5GtXPxjOc7PCPHX6WetHzUqiGdB85guKyNCowjyOgenmwBb4S9
7fVlpnS+Aa9jTH8zEnTIw6GEmZkcwmICv/IyFIfUdhhJDsQxoblUqZTsBfJFUGKXhnt8Liq+E4zr
oRjK5C3PW/44GRZhVWFNr3xVBorBhQ5Cq8XKEmLMRzkgXpXfrWJcsmLoJXrZuMASuXnCDXSzOQdw
zEVMZh0JxYStEjci4CG1YjJimyB24J+ChKQiAombZrZnVHwijV6b2JCSRM+05ouY1LrWpVvHDT+K
1IuSLCPmwGqjqjl3ohPv5LgA+PUaJno5gE7CYQ0xKvIVK+P531NOYGalCWNH1/0nKrZgNuQFWRnf
FEjbMeC7gxIoJkeTCz00cHyq2QUI+rCtvMo/68V8HnQiDMCqe0h4H0y06wpUEqeCA+8/37dhHWLB
2gWSrNEA6daYsxrlbVRDAxB3lsL5mPdkIIkVUu+Smfvy0X9nqUMG+JLaL5dQanGrZ2EiA3mJJM+p
1fR6xSgLFOJp+yiuPxGp663s574V5hVk5qkldGFNQ3xqIxjIgEnXBlyCmyg46ym+sw+ybBgvCn5A
PLFzGH4ixSDY8CNlI63OjBaD+vfSqMC5nZLQxJ/v0jQMcf9j2ifmlj3qFecL4lhbEbyKm7gdq1kB
FxXMLkricNkFplPB97u+kh3ZS3R6Dy++ZIY0wXfZhAOprPddtxF/MWjIAnW1j/6ROdalooiMJav6
PrtLwjMxPW9CPBYJLOytabgDIxaiW7VhEZ9pdTfdJXdE8B1EONBq2SZScPxMpnQZ1L37hdE4+TLg
vwOUuETzPO5YLE2xr5CI2AQXZvUpFho57A7G49mysgQ8gd1OvAFssM4q4leJzr3IMhR+2mEpSL+T
RV8dsEyFZIjKUbSs5KJ1wgQJQXxlxIyQ4OVwtiEZAnl/OI0n9RGowuUz+N4Bl7X7C1CZQkUqt1//
XaUkLJrFX7+Wng3VTKpji3jUinbQbzMgSzkK83TgjvyaT0iVQlJJZ2B38t9wdpGVEvKBgN3KooWw
cXeCDqLUr1o25Z4ecdjoigEr9OSLmLFuM6DANPWWiFj8vhhm3hm43SXzKPQZWs9zH8iYZ3PZk+Fq
BrNwM60aBWttLDp1ruQbO4fwR2nMk3/IKnX8LDU01GWDetaiWfSp8HMDnPYm8K+kiAukfKUEH0x8
+qvwf/pwfopTwb9J4xXXaJdO4YdE0eP1+Vb1fF5PMGfoaycQzhAUnDokFdg+Nx8d7yWB0iRnFZu1
WKFUTcHxL/pKQ9ffKmVxkltd2RnqAp0/d6MrxqZyq5RaJrT/GOaWoD8KSbO0UVxEX5fHz0mg0JWI
OZ4KI3L7fdqiE6w1S9VIsIMmiWTn9A/qhYZorYmHpXfEckcVVcGZo3kJraZpAzMh+qDAMgzitUgg
nyGwV/G77I8w0KPtwiPxgvUSDgMdsIhGlOTJXCf7yBW3MvWEQqVBiKs0hDXqhoodXlFNXg7IeJNN
01o2za5IXINOcTyCGqX7QI7AI4mkJiSyEG7sadxhJSBuEZW/DLMChRafZzaIWta+v6A4DAGMUgLQ
aIlLfJwO+ERGl2C8CjA+p6rKf1iRcGXKe3pGI97GZ+OKaTqRfhuClBJpku88k2vWKC46qNUv/XNI
3avdtifdbgDMNlHV3XCzFl58gGOVIsk4j/HetE43OOWCbvW4fWBWS3rwpfnpRX2BekMZSQ6G6SRc
OvUVnZx2Izt3wU/SkLqHEWMMdsltyCt1Wbwc3ZiZlhjVpFLl5Ed9NWmjzD02OBmXQN6bBfw4H/oK
+5Y74JI2tLBGhT5ZZh0tZ5k7BF08Ocy2C+EYdAP7Ig0NwJr8mLDROuk7B7699Vm4WG1j+q57kzbu
LVusT32f2VMc24gHbOxg7xjg2Iq6IzDiaSQNHsY8yHkepSEP+55gwz9CO1TWNjwuPydl426XG1VS
WjwlE35zSwqT18NVknlW46qWMl62/w50JpG/8wCWr53LUVNUgiNvQ/YUj7bY+ove1YVxL3+Ty9Am
300iSshs5dV7HJ1JRn3Hh4lAHuGBbkMkyqx8yAa4Grvp5Ih/SZMvPs2l00WFSHvkZXuHV6ayy4ZQ
7QeayU/8kJ+b9qtup2sGPEBUx1MBRr5N3VRwJK6dSr2kC58K6p0hvNCa2lDELvIE76di+EYi+scF
IZE/l7+7h8iNGnZJteqvIneW0GPum096IUyrsS+8BhJIVlrBu646eak/votrVWl04kCDr6wH7szJ
N6XATbFx9cQavNDV3aJnZxy7PDktChREhKZ1Iyiyin5kKzgk0Y1her3WQrZ3BSVLiLh+dSIaRXh1
+3z8YufIEJtKHXvdv1qxFU7CCAB3IUF0Bz19TuiefsnTnLKOoERfA1+H77wdem9DNpYrdplCLIH6
8EmkjqaCcPmQg1pp5GLqvn2zxyqVNL33QgnRQxiVNQDosS+XImWQB6mgd1iZ5E/9U9p7o7uGi12+
22crBM87TlejQSKXXt2Yare9Keb6QuFTkNVPxNYnRs21eHTuROlbjj241bA2dFKLYzjY8EEjjjkS
TKVpwfdw68elCKxAYVzGb9BmAXml1QdGXO4S+0QtzxF+VSvywygJl/RtoXvFM+gBfiT5lEN8sULU
GBkAzH6iVTQba8FWkeyIDAvMeYTl+elRql49iNcsylG56HjYhDysGsfmfvdOuvr2yxw6/sSEU1L/
BXjGqaa+TK2MK5PuhoPniJSH/UcGRh2VT+nwb4JmLWXRBDLmJOND0Ielb+W51dg37qiHri3PBAKp
BrDoaB1dw2+UohUfunHz1TN9gjDSHeeSFfxcCrTYJZUDhh/Q2aeHKUh0d3I2E2ZixcT2QbzmbFuW
54wVgRWzHSs02mty04RWsfQN7d/d9KzuR37Gp8b8U1jbb36otI7z1XgVZczTloa4D4kLsaHnRpdK
UDIT1+WLq6C9FviZeaK2Mhn0BNf4EnuASRyBPsQclbKEa7Uf8AVqEs7xibhBmmWSd5g0BCZ0ztm2
ti7s3V6NfUMAwll9NW9cEJQ8bSBwWZL1dT+nciaaYs3p1eiso51A3Ilnrsx4sRbSE8dApDte5X2m
N4b9c3QBN9UukHli/TL77Ar28f93NcZ1uMwEPJ9eouDsWeQoyvgRKMUw/IebjqzdU1xFupA5ueKS
7K81gKIY0IWqpwCZmPfyBcaqT2mwnQ4or4FaLZvaNk57N0we24jrUh0lKJvvcKJ3pHGEmydKc0ge
RLBWQxOu0FLT/9WiFUdClrvvsYJGU7gMEOcLBbtd2owPlyen/OGaT/0aU9uZLrDlqf2rZ4vO2WPK
IwgmwsfJHPQ3LV9u8FTaVnFTxCP//J2f4UOQVPGgwps7drBOO3HHhbG+8tbkcqOIMamEs32kCE93
a593I+kDkVmQy87SrIeeDPaKwLAyPxaiCWd8mm/KXvD1XMhfxJ08SMU67x66RnfhYx8g9dLLAo0K
Kuw7IXOs4VljMy3vVAMERRvyzHE6DlbjGfnrwKMfbxN/2q5dhPXvZIc5YFh4AlKUIB8NNxb/HGua
pvjab+9LmTOD23MQkWhTAzdqaLWlrPfmVz80bo3GkGUjpGX4ShcHeddWtai9u5F8JBS2/Gk38o4u
bIMOSQLFzzhnpEP4yYan0vp51Vo6ShUbRdHsny8srUL9C6hIlHH+C4Q3Wr8xjvuSeRtueMvcBCvV
CZi1VE69nCCDJThmiS8LwDdGP57uBYj3GFxLq48NrwmdNhqKc9j1nJFPqd0mGAljJ8+K4cSPbnDx
bVeZr2SGVVQbH4pl1gjg6lC2L1VP+8mrhETWxREXh7fIYg/80PyNAImVXMYXEb6mFlJ2+ian0Dn1
OTU+y1eic5PoXa0vAFIpfADh+txH6GJboPV2YZWNu5qRsRP++jz2CUVAbyLiFUtSdANyfOVnrAyt
xOLy0SKbTvYCN0/mAeZ0kJTYfFxZ1ynVCAlfm+DRQbteOHS23JKS/bVW33YHkuG2Hurntg75VbaC
BguT6PlXRIESwXJOxicmmK26CaDA/sw5wlqZfaWk3ujexHunkw9L2ZqFlENsRXfWsh+5RF9ai6UX
33fisnUOOoF+9gdd8LJlpymUcSqtYtbPaB0v+nADPW3Xtjf9kgmiEh9xhXVli2OC4RiYotIJINvV
Zv2aGD1iqTG5WHxixqo1zqP235CH0zuxgZqo7Ip6Vi78j9Z0e2qWQ3Ya3LcF6W+wtDLaGaNUFGgD
WItQyiIxKHUSFbznwvSSPrIU8ElMjgrPl2gakb4MNPymv7vEx/MW7LIf/EmU5gIZEJhS7D30GH92
PT/iggCiNy54Erp/+BX0D26q0iiW/MOn9E3cP4QmWh0g03ZjsLmVzeiO6s+F/0KvlExbCHkNDqTt
aT6AnvCDsRN5pm+SAQsO8XCljw8RA+3CuGNOAjZBCRu0yQTtzKkZen4wR8/KXaeggoqQQwgHCvyV
Cj43FSEDEYOBDa9nIAgtBgdbxat9+of+UrUZo3gbnhE6b5pif9k35Fa0sGPFgswP3MyCTPhgSc5M
yAy35uS17mqnoSqiT6eTir7lzA54te6QRJNx7mR0pL2cV/0cKyuwvPs5Vglowvvl5RiCOOkMbmZN
QUdlPC+89MSisxtGyjIf9D4xp7edi+8xMI/DLsmBkLqpxOe5mTzhJJeOBgj9R58tda1EU65NgSn0
axyEWJNGk0j9i0hMk7NGeahtRVgUtEqwc1WMV7DSVpaIzfQrfv0NLTeGQmvsv5kbNLWKJXksPJMg
OJ4Vpe3uuuatt4gAO5jCR+51S7VItMqFk62lK0YWh6a60+udjMP98UqQpW/sOhowVcrDHh7Q0JIk
M2nyG6riDXF2xFoNRuCrbfQX4XOWzfu+yyngrKhdCggykU8y4zg7jLlZmmIuPfjNoRRBFnCKEqRp
5HRTAp1UAaARfSMR5Qc76UW1uZOWDtopnH0pO0JC4GvwJe3pWZb52sSMvBD6SBqn/WmNpZkXFSQl
+Di/53HhzJ+k+IGfYlgNNdRjL6yajgiucJCn8qKomgy/u0112FIMdTES2+CoQnNgglHSjhknvHN1
RYuFF3ou1waAplcs1AUegmvhhCrbIdNKq/7DUpVqUI3DLgHnA3q9ULmRfqmKOIYU+S6c4YiuMinK
6J9YEeWdOAYtk+vroeZM5fn5OaMum1CbFmMrOon827MydKenHJ4JZqjeXaCQfzOEMK2Ch3Ly+PJ+
FrI58cJ1pqeLQk8nqCvR6OaxDNMUXIZonfAerwD0ZSnax9+Mu3yROLWH/fCHMZ5IQN4FZ2pNhNF3
BIbPa8ZTSseAuKxF7suqvge+x398JuRYJeKWEIHH+2jKiq5Zuvp++gNufQEvk03kU/HCyNXmKMc5
GwNlgQFTWGR2ENk4GrbMdmOtDKzDGzvSD/+2BuWUohr6LyZKcTTK8lrhleSls7cxlKeSPC+dVSL1
Dj9PZi9kKmLzpPUbkVUQNTsnc88XuUxFM7BpI8YqVw8E9ELvpkoiEm9zkZyst2b8nqdKIkN2C3Vf
dOukFvnkDyK2+y1P6JeVrhK3Usj2qazdSfA8Q2hOQasqY3J3R+fHVsSlbb/fEsZ8TWuZCa8OCseh
Rn3+9r+G0GIq3DnnJrmB7MyDkLf2LaUSXqml0LHATsCHBvSpVWKMgGbcwlr87soKYDISFJbfNhtb
t3F7S2XDz/7lQ8eMs1PzyQFyUkn/UJ0LDblqRu8EdoIj/UfWeK3XCKeHs3oHggKeL3haxOG7l+XD
NNuF1NuFENhZs8fnTSinkhLog68MbGS0a49bqMwuWWkmQV9+TgaBmqjPsE7Z6TgVs2tGoD7dr2eQ
Ka+4SSS4401dD0Qsi8Fe+1h13dgSH+xETGbBdas5KOZ/inUa4TkgZfNGtr0Zpof7zB4H4QYCZO2h
Bh0Og2d4/t4i25LwdL6XtTD2NYMLcHPlc6EM7B3te2+z6641diOZg7yARjb1V/idepYW2AY25SO/
K3aB2Kc8ulqReVmK2XXloA9y6/7CalIjyyRkLGtFvFMEBMjQ69VkWhxkpAlKOMVLlcW4+4V+H9yd
kreOrSlnAHynwVHNu1/5EgXo7Km2iDwiQQ0Ee36y6wbdUSzJM/fLQolUNzyIeVWcmAlEU4AS6v8Z
iRDM3opg/V2+lWC0sp1vq4jgTgc7TiBHmATb9bwfcyL2nJhSomwixJOhtRZFjaurxDAUWtsO4677
VBYhQrM/yD0I/dkkHCWWvyxxlVlp3aNsLvHnyxPtCjibzo3OgMOStTKry/o96f8g0bzSd4JoyLgg
/hAQo7fVXyvqMjp/9om8TGeWgM7qcE0JV5taC8PXgJHswc1/WgOV696vXGMk3/TGYIjFUZRNRkVg
XX0azuUDnmfheEokY1G5KVtN80msIyULRNzMNF/1lCFB+731/4YH1hTq/kkYF+WKWrMmkY6mwf1Z
+lKAMZsDig8I8KuM+hYTcOQlIuXILTKbZdwCKij5SLIsI1GqxN8lRl9a4PGOAQgBWzT+bj7cWlh3
cbfia2ahoHUE56DjP37x8AHENeC9EbRIs3KUMI4SLTUs1SpWQUCjdDRq1aABD9g/xsIlEbdYfiFj
zRMrAwADUzBRpEKkIK90eujTikNmMHAaPWqjL9xTH52fi3bJB0z/NcBnk2acZseLJyb8kBK6Effi
093Jk7GXpPyldUuolVC+huN4NurBVlJ8jMK1q+5LGua2cd8/WFtQdGboDO+LQEeYH9Prh4dni/GS
pAfmME0+HeVFg8VZhlIJDOzan5y9CxvwW058G4DdOjta3jI6Um1zfMLuew0PGSg7W8h3Sx/jeU/h
w49zhAv5yb0PQfNul8QqF15kQBmS3BQym0GaNfo3wIX9FWyr0j7JkAZ0F9I1VNiu9LL1ysNdxz0p
tJwvXT5IRw4TiSVPYq58tNEfHF1rEe4KEyjcw/rEhv4ZS+sHzXrnIipeI2ccvOSRQ1fGXfw3e9Xr
Wc9EtB9NB3R1JM4y7GwEY535O/RUHNF/qB5bDGVlvw4UOJhFP8+gHI5jkdo1xZB/WScVnGJFDBOK
vDjRvrFEjml4YzeV9cbfQUOPxbWcm+y5LFjZERNGmjkdeVojXspf81eXr5HFuoHLzb1IaZN9kuBJ
UpBILAWex2eSRaK4yfDz/xys09uhDgNkm23oJc0HiUyTCTNdkXTz4417Q7bJkaeloaRPNic+w8jg
IHNxz+IeGAn1+OwN1O7swXoeTqxYCycDaMnTO+7NZqIw3oz+VbR+o0UBf/HX3+5at+fS6j4aoE3D
dH5u0qhOfwBgasLTEPIonsYs+VhNNzgEvSYRKavsCYeV8ECvOGgP0tql6rCzofgOq6KJ8RQq/Efm
PSjTRrxRPof3F8qDl32ByeWQu8lWTwfsEiOWdU9tVW/Rz/9f5DL+UNYENPOILUmeR1ZxwudFB7w3
BqQGYk9VyKEB5/d+MqnVLcow0m7GR7MIfXjUtaZX/4N29gtdDgfdFjZkMyhw1Xb4UysORoAsIt9A
X9SKRNSdZxdfl22OUDODvr9EYjs7uD0yj8w6BehZYedzGHE8v21QMR1oNlGwUHg1mNM5KdrDAaP3
sJWtKXBytVj+JsdZARKwF4GmP9lVNNYqC16U+1CoR7ZxfbURF9SU/tbpXc32f6pPfc6mTLPSz9Qy
jhdlJQaoZqVUwNmFEGEIihtDlBpfG+vO1fc0erPP24h7b7Gn7/y5unB9IpbZ/nwRkh7iCMV06drC
vGF6oiqhs+WTIBPdGs01cZUyRB+SCPeHGP/ItFRzkWOhOHQ2LW2ZXxpdiK2Ni+ek2DGKHlLyhJCr
8+SYWjdA16nyYP2i8NBggu36IqHo0Sz2yX4ACn4n6DJEyDgQywjJdOoK1Dvi5yGVGHq8dDSWL/Ve
G9ng5ExBHXa5E0T50Sr5vAKyo1NXF0BzsCyuaowoXdlGBc2iicQscsa7PBKqlWpCnRz13d4o3uun
DesloxidhiUOIqBi//O1e+w4/NfzgFk+BOyTT5rkfriwmK9LU463+7TX4dgr3umbzaUP7L5Tl3NH
ilOwWZpc8p12+vuZnbd+m6h6LNRmveDqmDvAsQvhYdwa3m5bZpXcax4JC4NfChqld9EfaZT/FDbz
LY2W3q4YLCQYZ8Tix8+rgvPhRBugkkTR5A/30M5DjaQk8AkAtot7wwvmmeeAZbf+Q4uAUB6eAtEt
eNPLUXS8QnKm9ACgNgKsG1WtPnBWQIkP12lA9vvtlhq3vquHtlxaeTUCYqDTtnz0LWw3QEMgfGXU
uSkFZkr5Km7VUwBd68UhGXM1xeDEjEa+i4yGcw2ZwRJManHKh52rqYE6HpG6DyiTYfVZVkm019cZ
JgtURK+fkDJQfuHLcaSqxnHSV40fNXb/xSEksCVYpPE2vBE3nod+8dnz5XM5arNEJzZJ3GOq0E/K
1X0M8a27CkJBNuyOnse8MoVHhjHK/QVS8r+PuKWDCAVXNi8Gk2o0sRk04x/Txo9ruJnjPBIKFAbG
yvqYFgLNBj3Q6mbY3jA59zHOdRsx06iBVjYF1DP5RX5NcIJixF+5cdCsu0u9AZRzXy4VWD+HQd1k
2JIrZXnoX8M1BWacZdfNJ0Yuh4emOBwHMUFHoY0LU63kVxuKhiRUDbQAyyYbOqZZDIpN1Y6FCWo0
tIkF10JyTQle/6vRPv7VevWF0Ny3PFyTJXRxRPPSpC18dJo86k579mK0wT3noWF5ZYB9yb3rHsKc
szwVitMg0QCyyhW+OjKoeeIh05N/6tmgpRe/cavhJvn6neb9c1oO7sXxRbQH8eI6H02U0TNEngPY
Gi9nRD4AXt95YsjKFgGeq8eRGuK5njfCj1CrJNmtXNYV5xCrYXkyEIz+HuqMlwjNpBIDj5Vzmyc+
or+sBR4waqrhBQkuuJuQ4l96kxQf1E8C/XmVCxJmduQpMQLpJp1V9UUBRZbYl/za7EBMCe4AtTCs
1UujKf3D39OGTNBBY6C5YqP/tRgE7VermwRkMQNp71VhM8SD/BPSYH9KWZrvebNoEJhQwbVtT7vr
s0ZSu0uaTesJSU60mlHeg5sBuSC8o4JANUowCQ/NuE9WJF1mzf4KtMpT1LSzjPKXZgKag0i0wlVi
E7rJijneuI8pyR2P25pXY2zVMV4lIZzF65/IzzNpRsByuENlfLIHmxW7vvsbRU7XWJ0M76P5sfqS
yRZn+WbdScerL4XOqWws3wVygxO8yhuO7GdHhiKgV+KZfrwOlxbl8AyOgCY7ViY17xWuVxpMFw1f
+ZtzbNQnR3U+tteIKElTfrRqsvBeXipB/RU+6IPKb08yyX95LbpVegQBxa3dPdlUFAUwnOBqW//J
6T/fo9+nEhX+hYq1U09MaL9CnEL7qcQBJtFIc2gCNtx+pdseIPwN8Oy3LIa3KwIz2h9rry4wnJ7Y
96Tr81EvdKbU1d8WILzfuaxR2N61krzsQtMmwfcaJlFmq3V2/wplhgO60mC1vBfA2pb0i/aCHnDK
KGd12KFIj0cX4t326g96QsRkA8mc96LcY8BGe/t5lTH02kHmPZezZKJco34ySo/3e/qW1Iy/e88k
jAzrlGBNqb4bmRoLX4lV9TZrmPBzGgvZeMl4a54vVLjTBLNnZx6yO+jYoyDUGeTkAqVToS52Qukl
njiGoRbCRWd4WaMcD63bcdk/iFAE0ddOeFXcb3ZmO8eJEJc3aU1+OJOgf7vjGR5BJ1uU+c850vZi
q6dlEmxjhqnjFiUKC2scSxB9f8g+etBKRr7ukuLwRTS+M7i13pzPwSlMRyXCXVBPnMUB+OyzsDxD
uMpU3Cj/46PgAes2CXMCUiWIv3MtXBP0siI3zLWOYw1JKu8jRJu7YQ638r4HpmGh7w81Hjfr3Q9T
v8dGT/l3QepA7ANM5DAh7XaQAkTWM2XUYwehkgqAKDCe8jbiNZ9C2+b2QdQ5AI0NkCD58wnvVkuM
LCh4H3yfLwKsgSbvHSHErnua/WssL8JGAMcOolNQYizYen4gTBRiFSXxqnUudTRBCozheLrpO2Wz
BYo7sasb/Jsgf67K8uC4XMzzarzFrh2CEFoAidGBcbfuQEXPYFy2lLUFv8ysOEkcVOKmnNqKaDGH
7KuMTiK7ycVH08v8LyUqTzqQEWa4FYZ+7Db56kQLQA+0OYEgDqVoRjfk0awqdzLl9IchJOJbJTgV
qfiNlE+Fm7d31HLHfzQxusXiOPgRJ1E0tRq59Y3EX1PCEBqVK/rn+cuvhg5Z2t312ECtIwup6LsN
an/LJ3atugcDhEc+dkoxPpR+YFh4G15QnS1hqXc4hISwIoY7ByZG+iWppqSajlNbB10+KpuzuDzN
9j7eIWQj3mJWqy+OPei33E4y13JM0YAXMiB5MecL3m13ah/2MBGpj8hfZiUBBHBBZrgJOuo8/tsR
s8UUqKzmAAcBo7rG4g15aEmvo96Zj99PjwkApeWE8FnVXrky+slHsREBJYU8pQ/zmLczbB5Q91Jz
e9x62ky10N7xfSv4tcGKcLLwN7RCGrImIzt8LME1Gt5x1NXoHDIvyV908Rp5CEi6huVdbxg8DbXD
Dtpd5m+z//enK316Vee1bqDwPGCHBW+8pHaqeQi7/WyOdhwNTiPQsrLuyKu9snWr5zRtbByQMBzm
qTHWpdo+4Y4t0O1qQJ2w56DKKNay4RSMo7118vKVQ+B2AkMJetK62CBMCnlkzAambp4rA+aqlO7/
zSQAJXtPhqIEpBzMB+5zpDlCbv3TC4NnB1h8hO2lEnqo6iB7xZ0WYBHClJJSGBzItJGHw3+jJZ+p
zuFEHvcsmJaUuBx8tqkMk3zZM9T8FJjPqaz8QUm2pDYeJphuI4j6oz1o1uBKx1h8kynrlCKE+e+0
cKT4hJnEgYlbGk5IsQu+s650dCLIqnTfSHxefnW/bqiXZkTXUsHjPc3ynV2sKDlQJEcBDqgDHzj/
mtFAm4v+5jS0I9wZ25n6PEi4XZflsHqN7qi3Cp3rBI1zJ8PqBnzJVBlnToQYIkbS0e54NbEOXlhb
X2soDoZV072jSMoVhz8W0CtDAB70to2KDzSPiiRJ8An4Np3dnif5Jl6y/xgHczoQ/UM4SIsNmGij
8PIH2pLn6kB0fi0JBM3krD1VWYHBGSnU8QhGmSeI2lI+QlHUYp+Eotz+glMxn0kEoN9715mM3iVW
MPTuxzHTUfz4PDHsjFYoPFmvDPP1KkOKHB9pZn/+S5qdo1LZuXTuEGwsBywil5rKcgSbLyOBShNO
MmdRkQjKtYf68UixeQ2CNG/qezWt09kUaE9iLBaABB9sPaUpl+bsDPyG0cHD5/21fFlmBjaZqNGo
jP7dtXCUWLOM3e3Y/TGyQB6KYklMW/2CFN5oOHvBiSyJgJbGA9/xAMAp2C8BlJgBfjXSEAp86fRi
HH7V0N0ejnPTwMDP5eVK1cRJnByrxj0n896Mlx42LDssAzHUcy6JSRtAMZpKXUcarsLcawTKrPgC
TW7SFt8S5Gila5P6LRGzLXYJOIILUB8DTYPA0sKtceSQVmXBA5wyG4JEnKTaNjBYHmelvh+W3N+O
68HpfI8f1g501CWCN48T4gBUC2F+8++f+W+Q02VbPFKvPqoZ3h/tb0tYzmEQIU6eIvZV+N4hCkKB
zdyhe9C3qs8Mvz28RDWO4rJIBGLy7mZoci8gQI5vRXYpy3/Jj8KecjBk1AyCjEti9w6EKvU02k6N
pssWW2/dBJjSsAE/Ocerel67C6FFiWqhuooOsrOx7brcDTeaeTNvTLjaKx2ttzhxZYPs+UdtQC0D
lTDjnvs+0jecnv+zIFqiyeGDbEUrDTr2z5HVS3x3Bp+Lt78TkMX/C8SiPZ5Blgat39+CJ6UF5iZb
HoF12VI+aTln0IrK4+PbrOigfonxMPWY44qH4WBxDDWH/Wsuk/dMuAA7TFKjN9gGmsg5D3lqOgQR
RQ9z+7i96A+pZBO7Rw9k0RyA+9kSEPMphPPxGV2JGcyHP8Q9YLf79kiCMRKj3hHIq2dRRjSDc4vM
Y8DrbOntpAEWKFaCITO8zQh2QXDBMHVclXY5Tn1CmCirOkx0Klv/18aXfqmqSoHlveip2J9dBdaH
OSGVWtyKIP7ykGgQxcve1Sno/FzJi+USqzK6vc8tjtnSjMtKipby/vyWrdQuSP/4LA262xgIwuNw
OvPcTvLvVkUaZe92dGhNUGnRP9UIs2tNKeuZHUxsMGitzsT0zpZDRpP4zqS3X/4I/ytv6nePVZCd
ciwicj7zR5z858skhOLJPhWqdQrvhV9jXrgHUUMJfVkhex4V8LkWsaqTUiWZg/SBOEK+SQ6m7Yh1
JH02yY7KAr+ZmkSZ3tSuvlOaI4RAxQbusRU26AmluXJfYIkysp+so23Q3QZYflesAullU5GP8e5h
Ix/91HRzDMif/pSZz0aAB2dqQkudKD16C1Z2213kekXFFAwYF6pkkQ/MhOsKY2RE5DHks8jyHYGb
whEd2r6Mt6tFL6nFLv4yuYkn9t/+IaJnuPD3rKS1WmM54jd0355B2AkSF/ids55iYkJZpurBqH8v
r4hhoZrVnsOpe/tf5L6uYvBOY3nX10p4MOPPhIBEtZTODhJDfLG5NnT8l7pgJKv6sC+TGst2FShu
4t/3zj7bY4p3IzShFrw2Xq5Paiyski7KWH0KMhASByNICxuMd53qDlOv5Cv6wDLOUUf24dYcfWQK
Apfr7qTVmqslo5cv016bmNz1/uyPJGIW9VWBHhKRQm5GelIaC6K1uvOnlSuInDqLbFju6lcydw+2
uOsKx0Ng1c2vKuiR0njsnyngz8QHVijoe/+Z0XLCjBD/DbNE9vPp35C18rMqtkwxJoSolfSj0BRU
ygxAgVtrR0koTUfsfYST2nuXNPBjc8nO/9Ens33Ryyrm83pRRBPiooP2rTDoB1t3+QCJmw8USAYe
pThS438rFwfHy6VlrkGh02eyCxqcOxwkKs3bLAdqMFnDtpurgcSkUH7qnNqAGNaEBwoBpxRGWdcN
Vat56PnsRZvyRnByS2BhKClaGUPjoNEaDfNoV/MlIS3wTlu3/IAGxA0F4z8ZUNjGHICy1OsBZ+H7
1gfXvbTxOMlKUHeJnTzhsskdv7jHeL/+3JMl8LJEtdq+TkKIAou/LMWvYuXLsi6V4jZ+6ShUPsKh
4xcAfwFj9kw8GAL1fFolqQPxAIARdXip9m0E5/vB8vtz7WkpqFqdug0D20XDEHdiOESI/K2t+EGD
8L6U3bH/UTOcDCyEUE/CFfcOnfmayfuDqRMhJs6TrDCPct/Yx0zTWw8SxtSE0Ymf3c20uE4PoSm2
+vMSiEE4PDzUovvrxv+uVAg8ig9D3+Mj4llvP/gCKIq87y2scuZk19e9rCuoV/gPohuGx/cw8F3E
4D5e2bX8fisDDyR6JGpabBlGa54+tZiLnisCEEzM7XKeGmI3ZS4KQJSPHxJV8PjccZt4QqBHiYDD
C+TIYB2NE7vKiU4v6XkChdYfBsDSEIZfVHdDhBpwditPtkyeZ5et7aamnVM30AT9a+4w0V2zBTHG
IM0vFP5/owQM43uW2yt8lwqrzXu84sBk4qEahkXUGA4fl0cNsGMFOOB+ySi9tacGlDxqnYI+enfU
fvIzCc5ROxVvqTVXveT2tgHi6ztMbp+KqV9SXOcP8GgAlML6uGa+ov6NxBjkpvzjI3s6Pi+F1vbZ
g9gmMYcZzP9fee7li8YSOF/LqJQBCcatRnyOyHUb5BdWXBUd5UgaPe8fjLOaD3I2IDFVgk2Pm+iO
gp/m2kWj2/ethzVfvFl3Kb+oHHXgS6kLl74qRvaqiozdIh3AwZe/zvqfDmRrs1lp9NGfIQhskhoU
XFNZWAIEeKgy4u0pN2ikhWXItn1mC8v3q08d1kdNgN4QKu0hzKs/s6dDwHLTHk07/uXgIjJY/Zqa
50XsL1aiNDdpK41rDO4c64UaM18h3ypw367i+ChhVuGm7paWFa4tSot8gWMgAEWLwaqRj/1Nk333
iazEvxBgtwSMd6DlqnDa0tqJb0FyUA10E1SWcP9CAqCneyaQ2lfQrhKqZRrXZE3f5RbHrncg6u4T
0aXpItyNzZ0s75d5T4OcVi4xQmWyItM/wAK/p269o+u6Z9z5ykALj8EIvrgGQGg3Wsw38PZMAWNZ
su7eKb/P/enOZ7Q1jbZMS2ar5XL1PRz/A3Y5oyNK5xe3VBhHunjVMrC3P6NzBw3PXbMSJ+s8q78o
HgV/6r0TI2O59Qqc1ybj0lku61jUc04IWZzXlrqyFi9eSQI4pRt7jGaBV43STGPcHkOo14KtaRST
bFQrHuPgwZUPnBQERAGSTXSGI+Nbul5IXIyPf0jfFocSnm1RFpmsr6j4UEE8jyVJnCccVtjGP+CJ
ETou6aXxKo2qSQtDLAsnmchYTvd+NKWPv1HCK7XbyZ5djtLQJ48w+NaMgrKIZxV/f5GDJsCKGl0Z
KOmz2hvP8eBi9TCElBigXNt+RzWrB9CdkLQ2O/eGZUVO37h0S7Y1OPx0cfOGlBtBUBGtJf/5UUD5
y6B21xakwS9khHCZJRDuGVmcQIItU29UdoxpklH7sSxAfD6XEPzpCtXFx5Ezs/GehKwiwvjeldt6
i015aWv2V5Yjj0SlAiFWYVQcGNU9Ljh4DJb5lpCw21mFMA46/BZm9XpuUt0iRvdZOpIpfcy73Jnb
R6Y4bVsWrCyw3IP73v6RcQO1OWi9xGEF2jDtTYNZIj2wvoeTVHs8i/UM0SpaR5udkwVwQwzJ4GBD
ylMFQvIQ0q+xvxTyCl7hvFNtRcpsdDwq2qsS4P9VScZJromp/NAl0pYCUKzfSGwRWUnBmCazvGQz
r6x9/7+KkDQGNVHug6anwtVuPy2SBZPBmT7zfrWTAnWBOw+wSQiu3F6laBnXpZcHtNm3sHmS5e7g
YJJdsd2/DBGDsphv6FUc+8ZjimRBdUc2vdE5Ygq9s5PZvAKiBkcxx6qohStUN+F4LZ2KPZIRGH4l
1xIEQbIjgrFLwdI8gB8Ekw6fCiSRFmCQLXhBRhHEux+a+latqng9mtoi6/txfvSScoEKUjptXFOS
bKPh2v81CFe5KW1qG6GH8xNo2kc6IHOmMYzlge0K32H8upeODoZMnNzafvMx5FQB6sbuW1tymIex
PctEsFyvb7P/EDQEoE+96mhxKv0Vwtlx06gMw/q5AYberMpRBgoXwUZQKud0sJkIKEwfMhT2CZev
AMcGJ3atzj0kC+Ao98LyzQLJwQ29xTh8vQrUxpKftSx/sQGFHG3Q4XSlZefeVeuJ3faYFVYDqqdh
gvs5WgLL7Gte2ICGaj4hyP5xcI2aEDyvDmUPS2ZYQ+VCn2G0i0Iw7pJoD4mhRHdXbsNDXZ/5qs1+
hgh19obkeY8y0WcVymc7W0gZM8UxETz+Yi6SdH+wzCxZjgP5H8lraPSbGggNIHExE6pBWvxkqAl2
NbFoi3CFn3toJy95uch593t4KImg0w8DaUAYjhDw/gMtiGyNZYaYG3feLD1XWr/MtebKLfqo5WMR
ZCrLdECBSqPAakPUQhfmF29HUR1V50G99XvSm34O/WEzC/qKWXCVsVq7K/1g8En1kBzdgdX7taTI
c9xBhA46WmxaIbXfyJ/hounXMmnPoZP9KUuEEaXOunT5nZaVGoXdn/sTMKG5J0Fe7nnjhZGh52NC
CGHXQ30fyfpddcCHLTJSUwpRthyiHihE09PzlvcXsCtlXW6kslx1QKnzkx/4YwFj9l0DkJwofWFC
fpmT7mIHD62oDeT9XCsIheKkbeCXMdpZjvURLwVbV5m4hke3BjmTqcvwOvg9rGmiXpvfBUM/0aiO
Jgthb5L7zd7m0BdvY95onONWcZo6Y2K1XZML2jp2yoVhpMnE3zjIac89wofxJ4usxWMtxsjxn7cL
8m2vmf10+ol4XjHFYSu69rQx81xTKWfS9hSOQKBiW4MJQXiB8vE2hMJHEjr/685Cansw88UlB2z1
NoHanHMC2/3EN4mLBptJKP0QZgwhNvN898Amj2KGCg5HIQWnnxvgo+xIxMAHNhgxGdx/gieGE2Eo
f8MUDb1CSVlyfUHLE5DC9h4s+yAzDj/6RLE3ok63f/x5WLfjMSpUyWmp+1Xr1kezTzUwLvOYTKrJ
yb/xJZpY9HG5zg1oVdQOWSuqtc3Oy+S14mfjgqHMY1H+oXp3svb82d3lJAlIgugnGA0l+1aLncCj
PPpcZM4XRGFp0kJ7cgW5WKqwndS8hfYg7pbDslRv6gwyoNT2E2kYi4ktQq6Oz1pG4iqTSk+OdcNq
5IMr+4wvHIapq3/NbhKB9d8hMuQpW+5G3ICclbZoRtvlz/L/iLxcRUIv5dg7weOuqkoaTJMY6n48
LWk5QNxXCKUEi+83vhSQpHNCy6AbKuxTJo6jwI8MmgWhaHQ0hTeGmYiBLDOAGjqtoCbcWjDJlJcZ
j5g7UgQMalibugdEYP0uxVtV7spc/dce5AzQ+p8CA42AVsYdK/TSQtEzYsubLxbOX4TYDuMwMrAW
MuOGdeTRAhJ4egADzHc6c/jy7STRmpoON/aMaRkk0SGWhDA/xxWbx59xYZQlzrkEtkYbSUkx+jhx
CLeA7SrR/MiML5z9aSGDb0FKmk0L/Z5e3+Hd8CJH7cKqd15TENKhQBVwqAEvFb1RGTYQJzT1VHwL
FN5YaHx+k1bPiyd0SVjZlxI2Od8WJid+eJaQf1qezPEat38j/gDAvIFZJ3fiqehqTNkJnF5HFPAw
AmPI1qj4phkLccLXN7XOoWT1r1j2JS64YiiaeMsFwLe/cUl8YaHxUX0ataSiHm3VNpIg2uC70eek
q7eMd+b8GzMzF11Jlijs6pXuiypSOVAepyXsRovY2akao1D+iXaz9NOGGM0IBAL8RsdwwukHgmV0
QCgZsdrcgWQqAuNUgCqUmTN+aOu3c5QKnGDJ9D6/ufV3lnBYjyu7jbIUBZqSkRUNq3l8T0Oq9i0U
8yQfL8F/5Ffz52OCpswvW89n8WyMJPatwcm45snPtaYiFqMvGej/frwwtfUHi6bpKlL3+4GBzSvs
p9WfsEdZWBkmk4hCFC8Pn/6MrfOG4Sc9BZuYP80bUFzVDmNRj4UdZ9V6gfPa0k0pA44fxJ+lNIkv
hDcTE+byCY/8q4UCFQf5xWOJuk0ACjL9Wm9iRvuuLh0LzgTrP75Ufp7PbUVm08tuI/QZlVg8WXqZ
vxTXzIlPrnmgnu9h98SwGvYKqRcosowa+KIlN3vTbQ3X802b9FiaRRFKDCFu3j884ApT+G97Vbls
ucOXN7thMPz5OvRIcsNhROmiv2cYak2D/pwxWkyapUI1RPFr8giUJteJ7/qE1NF0Lb2WSVOKsnNK
SkRZJ6mjgCRBvE3VAuf/oqTOJ3/ng1vPgBDRgJ7bdvjSiXZZGpT8yw6/ajsUVOg2g2AA2r+dLSDI
HoW1vXuY9RvCGNLJfaFfzF3vLintOQB8fcR8/sIimc0lfJWOUk3lUwUlPmkg+wk+XuKfIsRamXrU
TmLCvI5/fcKdHP3HTBI6e3fgPVfV/hSWHGTajaPQR3w72jGlVQ3VzI57NqfAT44+fnj+LH6nOyCV
ximBWOXfDh40+FFTz2+/m/hecwj3G7+okinNRqbtgnfF4WY7vYYI7wE2/E3ktX6npHzKwuCcNodG
bY66DpOzfteaw2nStAkoo5exE8lAr9dkuJ/1GJIpaNUS5SR0tqsQ983pP3pBSSiK34rthKVpZKbV
E3vP1S6yvLMYVRLwhTw1Fv2FRCqlj5dStVi0JkQ2S7LAN5AKkI74c3bBQgD5JXVEHsiwrp851xvm
7IyOGw2GWi5WYKJDfcYnqSdqpgFgSOsWbhKHdqghwDLzPnf/YpwYZjAOJhUE35fGojmV5vEpvNcA
MGLdk5SGlTEF/ftRl0C45B90TDC/jqthUFDCGkDPMi4ui3gAYkxRNzQmVfWe3kJGJWyGr+vCSUts
gdGkdCnq+fRu3Bbmc/ir/sI9iqU3NvSPRmjQpqTD87gK7p0x/WfdmMYskU9tbUmf4Qm1hYtiPQwV
Ibjri2EBCslntfm2EXunqHzgReWXKu9Km64ZBWKAJJcRSWRz+EogbfnuBwkahBfJVlMPk2BjSc6G
D07Hjn1HXEb6DjVD7jEduZ+pj9bRy9/Haechc5yRrKgL7Jt9TCtNhMGYxwAMPCTn1N3IwpHmgAET
LG+0/tzBftHQhRCWzt0fjkzHV1sf3/MDbK9XDrzmSkLqpmTDFOfALBrnQUuu9pkDcyqw8nEWFLVO
/klo5S8WkWWyuJEg9l6Xduz5wUL9kOn63EeWVfhz0NnQAF8BmRWHJAC8unEFgfk2qlRvZfIAoWMI
rGdsxT5Bf8a2nj71lkIVvdZUWrvfxeqM42qv8JFpEvVvWeY/Fm/3Golym9Mn90oyhQJmG/yu6bsM
ggVi6Rzx8SS5sNr67wh7CkQwkq49xTqFiPt0OATozRBRHTO2jEIgx/Wwq8g5QtGI5ImNBhn/OFAk
je0AMPOVX3FAHLSI3MK8yxtT+UiqNLWvRGslT3ZjybMOTAUsIowRgjZ3TJws+843fZhWFqtj076r
kDJkZymKcUfKz/0rVLcTP/EIEubIKshauYGfeJGqygDnYhjgwgnPdtV3Dur5CGkqoNfxLqELpzWn
02ir+aFv8ZxcGT6AIUlNf10zZ8bl57+fuD9v7vdwr1rMTL/2JWNywezi7rcb5OD6YgOdaWvELFgD
gQZlghv2CI1Wle3jDla+UbQxrsG0kz5o4NHl6FrKQ0nBQ5TLoDDnkNWtnAyBqLGipgP6H+Uddm0M
v6IP8ZoatwRiB1QA2xNm5dwFNyFc59mDFe6DdxulgQJUis2b3czFctln/2vUd/NuIlPh9TJo7w0v
97mD9L5Q58iA5+cnE9Ah4YgVV14Voz/tr2PtD6n264ZDSJ1s+EQTsSRQzkkdkENytjgiOavnqZv3
Cd1UIEkq+UHTZlORk6Bbe+b1j31p428nXXaYQjCPXAECLwL6dhIhcFumCELKN8vm5Xg/qzGqcPXA
++bSDMGtM0nb7fGymveEVwnD8CDiO75LaccE4Xjp7KVwTIOzKgz//2wXink6rfeIbQxbgoF8AVEu
iCzqBlKlJmdxt0sJaeKwfXCMbLBTyWZXvmeF0pEy+j/s1IjR3PYJhAT3/VdttjTweJEWSsNYXRps
nuI2pWO/Xp2RVVP8UgPW6UWNtkt+J/70fL14uYB7EzuYxc/DQrrhw1CtxbLDi2/spBzI4q7fpNw1
CZxHxb833EdYSW/G2HuTknZDZze4PkoWojix0EMW9y8yYaf6dyvwTM3LrNlhFxkbh0chTOhzHtcA
O+/5kHQoRoHrBebpTFaAOzEsbyWAh8pjGLwBdIdGXcG2RBGAzKbD9g7oQhZYCr9x2z2tlNYzrfZd
efBnKxL6pWvB7gB8uGf/GJQFDVREtqbXt5TVbIP/fV11VZxqB3OvEdU5aaA3wW7miN/SNxovb4Ef
uGl2ao1Wl0sBfID5CfeQe0R4aSocy4jIbRTtpkPGviRXwENVpMw7n5WcVx/bBXcRcK5saVLvvzDy
qnJdKW0Dl0Lc6vU4GJn+N1iL9oL/VETr+6pH6aT4jN2xOAPRUdoc7Vks4YNQAUY+xRc13xVoSOh0
lLmGJoPi8Tjf25PKWMszl0U0sKl0pfz8k6WpH+qbX84wh9LGOjOW/Ecm/eY/Ue7cWqbxlxIj2FSN
3+a8BhhDSNEsRBwxGX1kr7fBWQkLmrQDE4HkoUGw0OFl6zGLbb+x1xrBgO8H/pGn/bIAZHeWpNgh
Y9+WUQA5qYYnbLIilyO++Fim3tZnYTlI9twfJzdiUV4jkOqlevDgYJmWgS6PJ1nwQEekbJpcu9gP
ytGxmkNDCMHYdU2+iKxBLMYH3TVu9hTmnjp6NYkrv0P0MDtN+dxoh+9Hp4YrucEgstVv3AUsYpFR
53Fw5KwO+vdO6w6SxEOGibpSrsw1JlT9BV8E86nnNTjVxRzdCWswaOg05lNNwTncplntEGH7wpRj
FNMEK8lfsnoxwo1bpbZMLLx+rwoklSC0lPPUqbHFlcVs4ae+oKxJPlPg3FMiLFJ9mMib5LOCLvf0
6drThoLk6wSLf+VpjP0q3xj2SEV5ujoKYVAG6xddWGlqpkKAHuJ8aahwYDxazpKA802VZTAvxTBv
nFU0ER0hHdK0qfmMX6Wt2PpdZEoF5+dwgLf0nNwJ1WhTb3bCArEtgCXXUEgRm9O9UTYjmTqgOMmG
WLPpcg75KQTsZd9VFsowF2tleOgrXCrUWcmhO4tMg9aHlpPSWj1r2KqKhn/2odaGxo3+T7QWdV6I
xbJk6BAK37Oe60MUHWU/R4DAANy9X0XI5RpsYqDrsJt1xpaKVGrQsPOmkePk7tNjXiVwGF7BQpgS
m82D2x0j57ZR38uZ0P8pWhNJ6kXWxeDY7QceQrjrxiMpdqk+/WA7DemU86TgCHfBvSAIZ/aM7/2C
nfOSY1UxST1Ix9oKQZoWU1uiu6LJ5YekQxsPcQ3ahcz4+mZE4HlXxcBKPY4U+jQDq9FfmRDLeafs
egdIHMa5YTlLuY5RPLmF88r57iNPMWTCTcJWyzpwuwT8Jbr6uc4oGY0Yb6M8szIyCufcqnF2DS5b
hfHnbnbZZonMaqJm3Q/nUia9ZyaA9W2+FMCJFCTOJ8HbMIC5dmPoFpyvwAWUNPTsoORGDlq4sVuB
rzy+IfboJQm+9p7QFOYNrAnJ71+wLIUd8OnZpJGdxEAmyz33mS2PqGRr9TKCgHqiadsE6Ajr3INi
WWv65gpyQfhWZ9yrTpRE/6US4tS0BAoCsdFPo1ndjwmWlkfyQjbZlLa7SXT3ntaetmMzX/w4AmEn
ajTdqpx2Fpdvgp5yljntkhS3C5e5jBGLoLz3UOrzTYx4wfnTPljlXHy0BWEp1WLL4oUu+3plLVIH
2Nu2vfrxi2Rv7hb5tVl9QqBz0zDoKBaI/3k3MfCpMVCEvaykp1JEgsCuA2zL+VE9ouqcrzdhPjwl
bCv5K0Sd2X1JFAqcSai9zZtjflS7sT8x1D6bD7QSlHEkIRubEozymx0L4FZxv076zI4ERgimGKTi
fYsDUglVUWNoyARkVGdfH7WAZkG7vV0SerIwnleastvXhWvSfKmXbeHjbEoKY7DVtilrDaOWnH0R
KG7hF4syIWLeaHUP+p0zFycLbw8E6O3NQouh/URCfmSc60n83vQusPlNvBcjmo07ljDxKUrYOSG4
9kum7hG74FsPvj/Ls6ytskx5nJ3AqJgnWDG1edh78NQzz1+orqTOCUn9dBvyx5IpkuuswARS1BGJ
U+K3eFVXp52i+2DZKqGjKxmNHchy8vRjPGYflODcLMtTDXP8EJYw4vnrEJTfvv7fmqxKYIfqEMI3
CrvyhjhVVMRoU5zIvYt/lM33axlpUoWWD1D8x8tYLbiYswDQk9qaH7pWgXmrpkzIpYqOhvHRvaw1
km9chFIZHV7pv1PArPi4vImHlQnsHa4NhS/fGzs5ZTr0r+xhHSZaehdBq56QE95+jPCy/Rwne4w3
h3RjU3mCLEpCH7GgD+dCLuT//6T2ESkrBekFxDKqr3vJcvaO9BiYiLXti8om5WcaeBS+2hiGGjyD
CF8VX7d6BSgx+sfeuDi8mVd4vAJtY2rYRJLi5ke1V4GqGzCjrkyQiTb+zJDT5p87zX7NNFBjr8rV
6uFCjQ6isqFY9hGSZnIPTaB1ALX2UqiEVwIlVZjoPTWP9c/DJJjZ+AX6BkCKEVoV4B5uB1txiCCb
P2t/MPrYPm0r96j6yKtUvar+WrcJrn0v5fJ5rNlfLuZOZRu5FevQyX7V2+BIvJjzITwW7h+hVD4B
LKJPsAWXy0ZyC+prFZN4my4tC1t6fVBT5SrvCmll/65dp/Rus5VHeOufbPCC2cBxXg83/ItGV3+a
eNr/2VEQZAJgYXC0fUhwCAWmrOXdXRN+ok62qqGXj3DAOwLTXN7ktKGOHUz6SdPsvoxe3fQVzBxg
5KdVa0xEsuyYgfn1rfix2OAChpN+87eKLWDxarjuUUx03ca9ILZngrHpVZB0zcC81HT7ntPMMRqp
linnPUSEJt04IslgRqj6p4bTvbw06uIMKXJVlWAXiAUxZgNg1y05hjeUS+dVLqLYvHI0EBkFp04I
muNcBNHygQ5ZEmHvJmTx0NMU8aLfr/f4EuqjeNmm6DCp0UPrEU208QOeDCpXl95rFvQD0XRGHtlx
4gFYUFyQZ+gnq+idFENJGYONmLA281Eo9vwt2y/TzU/7N/66suBeQqOPflzCXO/slYGBWG0an+ml
5cnlZM/c+t/YqKPZ+ua6TuEAVcwigfNavsQj9UGyaIxywh//mVs0LZg+Gd6BqmFxMPhUe/gzguE/
5FetIAlo+4gOUujKYHGPW5Ic9FyRK0cgdR22T2VLZk2CTm9Qwr+Gqy5eCLjyI7Kr4t2EctEGbpTM
6Dzkx18w0ikebMyzgxNRZWxwFzomc5C+P9fsL57DnOQ5azfn/wwvqr5MdIScwWIFvYX29vxfAeOh
JGmB0JgJxqeScLmyf3CVEywy1F3UEEWL6/ItjvbyViijvT3fPH4ExlC21Gf3z/QqNoB3xOqmuWYq
psgcR0WHoXHtBooXXfFA6TceeClMJVG9xkmuOatbj9TfobGThBu3EMGXi7LI4fNZ5pcCdtLAgNun
7N1WU4+7DHxiPThvc0cEsRmd0LUpsIPL0VAEb15OdrRGrHhPqrk3I6JVQpi1G9gOiScH7FS5hQOV
7GPsjl6hOGViRNOYbDwBJlp1A85orpOxH+vsNrszCyXpTcsXOSVg/m9Cr1XTEyPXDQQeF3BbxEsK
vGHXWTwNFP4tFwW7JP7Oz3SED8r6OWSojwlwbZ3TqYZNMIfpAa7Go0HMD89GxMofBQAQTAGUoV6h
xsYQpUTdMU8jHkKDz/FOrlcp1MSVzipVdsSJJsx8P7/F4HnMHh6OvhtNye5Z72iFOfhQj1RHB8a6
CrHPCYuyaVfZm7/wpFp1eU2uWtFcKdDJ9Jrg/6xzxQkSsesPK4DLM/gxYvTmonyXrVRFdF3LqlmS
RAuLZ1U0hvmD55Okefw8gVuB9J7m1YfTlzeSAQJPgqk7pUaqjBLmc6s+vRshR5XJqRqmgaHbiV3q
W8LiqJgh8Og0wgFMPInOleyy0pri0hKdisVEHggR80poQUD7k078l8BVgqeUD4KyTYlSSqGQhyOD
WWqJdmm9OztaHlrJFpQe6S8jXJk9i8IA8d0YDU8xPNwlvatN2xUj1yI/jEEe9lWLSyYGzyhRoD0D
SaByn3oIbvepdvdBre2H7BuudYhqlSlet+OieS30Cz9pCburpFdl5eqRg2ixCQj0IZTg1hqQGc1/
d0pKY2NjR4HmQc8BGRFFZirJXMhtkjfzikdybKujzfmLfqMCTKj784cCM2dsvZMuwlhogFJDs67j
N4eT+9FRjsHXF4Tb33PilxoSdW59Z52z1hsL1A62Tvm/9kaHPPqdj664j9wWgZaCFHskoVPlnZ2P
YoJzwN+9Bsj2v2izZHBwPb8gxiNF7aOJkYqyehhye9ntStpaKVeCCiQa17vt7M3c8ffpkxaMqxw7
CLvxVSMFhr49VnkTgXaAMxol3rn67FOyh6qQdOnkCXim1nFRTi7rP7938tUdPKsqLIHrAUKDHVv9
mhQsdo3kvQV+26M/U2KYgyDzrNWD10HYOSzyGZ4cNIVIn6WGxkxEHUwjQ19ob693NxVKy5lC6QUd
ieL7Kt3WeEcdu0Chv6Clnk7Eh73DsPNli4afgo8P9Sb+I/9LdqcfCERD9LKjC8FP90dLK4B2VZE+
RItkDKx9RagIk4Th3E1rV1QkeHZT0GoBqUQ6zxb3t3dg+jj/SthW2hHH5s7+masdpnHBtNfCz4eB
3pyKUKmpz6TklL30ncE1RpBqgWk2u/hdIENxUGgUwINMTXXSv2kTa6ZyEPAGhFbKRHEzMPL3BQm0
eZX6dLbW7m2eCsxEZzL/cvYxmcj4geLuGOWHnoZt6QNyflylTykn3luZlnL/+E1EKtXXF4woXr22
7CudMeU0H4c59sQckaKctT4nH8v9885NNAD2iOnYbJnZxRvmzvU8hXsv24eCveJVNgrjCnXN4LxA
MYNDK6EfiZB4KmNNC8EwI1oPtz7JV16On2psd9f5lvd8D++KgCp+PH2jO6NPr4gsZYR6LDUkQBhw
W+z7h9Ifp0n/b5/ePJpU55uGXaj/y9c35K8I6wqLanrv8IijH/8Ve36KQGKdeD599wnoQy6Wqrao
Q1Bcdi2JiuLP/zB35Z7YGqiddpwtr83+mUb9nHhkPYxMwHIDquLWx5kktEJrGVI2VNOAkCOgT8EU
5+tRC8+mmzjvbwJi4vZuC/eDCau+zOPSSe2u39HdeLjOsyuU59RyjEyv6MReBJ78BZqyIVoCppZ5
KyD8maxk2QMZ5+bgzDNiBT62IAUEO1YhU9mWdPGczE44wooHN23e696it4uBQv6PfteWljrtSRj9
egE2/B+Rh4WbuQd7Ec8rYs19nco/SGJ1QdFoHhOsT1AtTITI6Ch2YfY5JCndGk2FgucE2Kdx8AbW
EKXevXO9MrEgg1iFBgHbQUNavUE88dym+bCMf6cV88ZyL0crgGKoi7LW5s4RfJT3DbEwUxh792mm
O7+r5HqBv+dij7RzMXfctOHXoZC09eEw2T/BWnN5HqBbLuMUMZmgiwF07yHn+ur4+q8x5jOqO46A
s3M8YfK99Okyg4GD9hRlFaTm0YTDiyhRVfAPUYwncYQ/jMqEBiCQ1vXm4dHlgalTKYAkEYyp8Mgl
yBpM8J+xeN4qyf/AH/tMt8i623XMDc5FbVOrtL0YHzjD6GnxxLsQtctLww89cYAs90sHKYJiiXsH
CUK5ZeQj3mTXuNh55iVCFGPz8jpDaDeepj6dAfc6ErpxtJcoRQBemGUWSYrkfw+IcPCfb7TiXQhu
FuR2uV0a82gFr/tp9zudJSSabqacUU7gUx8njT6DYULQcebE/NoNB1oLq7uCeB04OK52x8DxCWTP
J3pq1aeUZGLcffB+ICJY1uxVgE/p4ciTNU6U4S0OuUW9MxxLWQg+YK6tuuNpY+ixuUoqtABYzfYq
Uwe8qrtnQEf+8VZmzj+Dk8PhxMroFU9dF+kTj+sTOarpQ/NRXckSv6rT39xD8nVpGZPie4I9PV8y
8uTwDu3k3AKfb9rPDJGeyRrdtWOWoIvIO4Y6N/SBDlU6sijtkedJEhfa3+T6mzd9oc8q7vP7yINu
jArBqLuQvTVt5+fyzgj7MqwEVtLS/4PdMLb6QOD86JN79Y6pOWR0BNeVUSv/trzl34LnI9HPInEN
dW4OFvGu0845Yc7TdEZ7kJHqBhh/sCpCDoWtNe66TyVDVwbRLOhw4rlaoTy0Yoase2d2HxxTuM+5
9hyJIeFwmokKpgrBBFusviGefcgjHHuBuY+3MWHoondG2HtvmXeRUoOd+b1SEvoVK+o/RDtxtExO
Smqk0Bq1agk5HDk555F1dL3H25rFvPGl46dQWJQwybSo7cs6q/7PoVRzBIMHLmF0o7h3RaKjvBV7
Kj3mUwPHsf0rW6jt17z5+AM8dH7Ka3FRYOXYxaOpDNn4Si7EbfN8cU4BIPZxdQ42u/8XbfOKpOPK
153gFPATmxshemKH+S3u47/fm8RBz+zOw5+/AQjngDoyTu00XuhlP+YD3RC6IVP2v/2LgQj3IOHc
LHsQgNLindpEaPRljtGP4NsunIvnQ3GCpqiCPNUxt3jxNo/M3yfSRi7581yPzYF9wyUPJRL+AJ0r
ZACbyDwlQDB0CVsbFLC48J+wmANDTgvXfVTfzkNKPDruJHOHDjAiVjplGu+DlaPKSoZQ+qMu8wz/
NNOW+CvFlG5LPd2IEI+ZkV3AJONdGyKp0a1FZrMCWTb/dHAlBZ/ssel1UI/itTMz3zdTFIFiNoBB
qp32WzY8eAIiqnnI1KRhBf7RQEkdcoxlCB+APu3zo727KQBKDraxFAA7iIMKcin38AeFXlVwE/hI
wT9EPrg70ux0VSMC3UAXtMzWNIdCeZ2IAre88b7CDPuX2t9169HahrNP+26jIaeyXlXGQsd9P2oI
jhWXng5MJugBxPEAY+sD+UEnJdzlglAvzCbuJJyijwDo6RBEyOQtaRF189414tD17IGgPqHVqWZg
wzePrH1ZVpIrT//+eyjnvgvm1Xh9CavkAHWqGQ9KEgtWPnOqBbp7kj7sCNq5pOUVWnn+eAlTEJ9H
XMr+mY2bKcMhy3m9BcJ3fBUgW6mHLhOba27iL5IqKfq9m23OkmazmKfYofNFO/E/Kkhz6t9hiWlK
0F4rWPQ8iZX/KDqgfNz6GH7uN0N1KLRo3Pu/tC0GfohBkKC2T19T4BzRLCkkgQu0cTxV74MJvuws
Han3LCfK2CkPsfr0RiN/gxCJiyfs+9Hdbdh4DLWY/U/gCJ+loxNHTLKBXgSCYmare3gfvpsdEURd
px0VHzkSNfPukht/w6778Qn+aRvB1o1yYy0vxkG7EWdX6FOliWXq6eLwgv/21d1GC4L0pPVynrj1
H3YJzPq8ct0GLbfhs86PSy4XjBFPjI7jHiRtuFvm3C8+BErw52t3mYvuG46ap1zNEJHbbXnJwfg5
AFbNopU0korieVn7aguB/TLB4klXW2CROEVnzNbAzoDheR/Peeee8/4UB00nYnVhhadOyn4iZ0v9
2mEZTaBkPPjQ2EBj1rU+NGmkTjIEY+ZjAkB0Mk0CDow4xKvy5aR9RNJ8+HZpXITqEwt4KTgt7XPF
u0Vyf0qvA5MXTQ/gQ4Rp8kdKJo5GKZB9vTISCEctlNix55toeZVa73YW6b+YaCG51R08ylEc9x+v
S6SE1s0Bd8pLJmIkjdzFSesHDIQP5+ab/mCqqkvDuBJCxJHZX/RTEjIc0Ba2qJ1NJRUjbjSF6zZH
uk/BuBnwxjrFYgrS/S7US+mdMPH1h91BPsOEh1ElnxBq+le/MQbMo5WK0M2yCZ6Nxv8vxLD9odtY
cdf0BZR8cBPAKtdSbzzo+qDLQDKgKDSSGtOc20kzcpvPIoePo2z+M5BJCITG4L92irGzrvtcpATg
z5QmZ+/PfwHDb1nFZOWZ+rF7XrcB0ZriYB/KqWWE64wVJOSHanmGOU8TiY9Xa6jesHmQTyHu0k+/
BeH7VdL37s1p4TfFcTEGj/8FdLSrTwJNNocUFJAAZ058BH1ZVKwJzddJkFRjOTbHomzC14dd6JFc
4MMTMNrZrN4nkInTlrKR3/isjicBM8tzO4Yj1kVR9gqtK9RaJ5b0fU4jUngq+v8K4xb3ugRkBYXV
74CyHYvptEOh9zVRPB0xtNKftGRUS4MCKUN+1d6G0rXrKN+oxIBCxcL+sw7s3CC5yZdhMLxD1e4+
3awzemLiwVsS23uAlBY/RAzrLRolq4Hzc1E6sg46DeJOJRS0i6bwDK1Nt5poTm0ahj2esLxiKOEo
kA+ckatBnCbgehgvgI5buzwdhjvxr9kewGEkYTGI/PmznwdUgObxAFxkxmYL84V1kokKs62L7POU
wDtfXrw9XfiJXeIH/Me9d2XHk1rtcHZltDRl2uP6jwX/D6fVWtBs41xuqc/y//c0pejYfq6Dt+01
3Q62su/JB26gIkTl77LhdBAgqCL5bUgqRyYtAZ6flOter1hs7G2vnQs/nUcz7eMqAVs8rS3vnfRy
9RwDWosf4Tch0p+V2bgRpSOoRvkCLiyB44GVFZu0H0yscs2ANBqH07IVRZ+A/gcGHFx75a2eDNqw
M84lLus98SEWreW6GmQTf7pSATdg3rFVlLiPv0vgOInkuZB1yJzDaiLLAGFvUzx55BktZZeyCaZT
3NqOkObaLJGgzku775ZnFIfb/uQzf8UwaM6C3xMH1MzVt9nD6JmdO2ojj7zCUiDbtSsGFNjsPkn9
VqXGHAmhhti4zhdKb3LLMYTej8I7L7/xd/byvHkSybylfBfaGk/yvF9EJiQFleFK9ZgOWvkxEUXq
9Y+msv6DUzQrxYk4eaBNE5O/FdBjrj9h4nz/sgRnS6WDBEGi7bICf+Yc4cXkTEMeFhTOl+0kM9AU
3+Zmdf5zoEPcYuRAW3jy91cswVpGunHOVq2av+61hCHHoGN2wUvufBTb+pHGZFZKVeYHz8YmRCFx
K2duxOb4rEzaaFM3WyCGb4Fdsz1whUdFpj21V/oLSf866ZQSf9Kww3HH4dFy/OTG4Gqtq+/7ENg7
8Rb3orC2/O55zfSeAbJ8qBWFv0hVI+d8xSBM4cKIb6/BPITN0TRyAI5ysIUxXcgsvCHlwRXX2kM0
CwN6WmXr2qDkbSQJ9RlHyO7INDOdeKYxeamrt6zCwAP4CJ2VBwHwKxN1HjuH8VGH3c6ylPqv91wD
Ze4JO01rr2psGtvsvzpM50xK8xNiX/22fBDL7i5KET3o1qiu3TnE+FYqDn0AS0Paax8wEhjdIBSm
G0mPWktELouoxQIyU2RxXH7E1Ki+CYlXag+U0e14zh4vqDMEzHoALbbw1mOpwGVqtrqq9OPXvU3X
qRU8PvtDLszmYQsKb/PMmxPgCzmLLuUAK/TAa5UYSp5fZ/aWUeQqQwkpYDmFkVKR8etm/FB3/afX
noqTnhl/e07+lSVuT6yXFBvj17PAPuZp57FOhaAB4mE6KSMnUHF5YDQV+KTCze253dcOj4dY+CJX
c8+euWTCKLL0JMkpGAPAlsDN2ac1ejVAHhmX3iU90+Nxas0jAyTlyZLJXB+svIM4UWUf6CWcBb5F
0ybK4DDUlnmbe3wr0kEVT0euM/3pnTCTnjOM+WjPmSkNX9TP1lo7mhojEAHVPupA1gvb8QV60d57
pcjG80OXK4RLM6V9Tv8pZ/PfcFt0wWyY2aC6vbNnmgzY8y4ukqzn2cMeE5h7/hsV4cAGb3OuvP7q
7ut33NS8EQ/kopT4Brh523VMkm/IN0K/qCCEMMocyaMX9bJDmZBH89el/XevsHr3VujED9ofdTVI
N7BZt9X0bw4LGuYz03zIRuRhDzve2hOU93TMae1tMuEo5SWfWCalSc0aFNKVodARZF96q5eXgTY2
BtNFMjor4x0u3r2oj7CvGSKaPnMqNGBsla03u4fNqU+GAcwqkQsGllKQKI7cW2ZcZDBq1QlAAh5Z
o5/dv1jPU3xSJHLVv1WY0HKoaYpfQOnFv4hovAGCrf9eAVv1yz5rDVPECakEe712r+Rk1rhVHQZ1
iUymnXSJ/nuW3saPr5vIAJA0pUCZB/AvM9lUqt4Kimc/bdvq07JpWrSx5mKUhOquyG8ZJpnl3Srb
3CVf0hR6OjGfpGcQR4U7vZECKaaPGcmUV5hQCkpGS1S/bX2pQN3uBB7GdEFS+21Bnw8SYBFKBGZA
dx0nijkuXM8C6hgeAQfys5YsOVIAftHYEAqB8+buzEe5X4DMhlSjD/WqgMPWdM5jhooe2Dj9jwmK
v88vyAAMNNXq3YiE7bk3YT6NTgpto6Oq/EC1pVMjCbkjyve4NO5hTsN3mH3qswldTSXFv3kib6I6
aSP+hG85F/7/Q04RNEbs1MycogdxKnjcdJcS4vIfauQp1bG0MflzeiBA5aymMCHiEfHS1pljGBi/
KFsTbNHgbAXE5WV6HSlwVLKUlqrW/HlBbOji9bkr/soLFnVw9Fq9sVplC87Tj0YdblphfspHWPPf
4BbiGrDUjKkOTocp0cyvhArXWLGkXgnV/s6cX0jhclqJRVgHC/xlGoCCd4NH99ZQdTUhF/NtilVs
tWiFKeY6z/CnJsqI5y722YKJQuj7VKwaG/VO4T81RmDTKZu1LZXfE1I759JjqLUM6wkKnbYVoBkp
Vxdv/KM7+zQoL1HiLxFgpMiCJarlFDyejV/+PUW7EGHVWeW8sTXlKcOUJAU6vgX9/pXvwQEGJ2+l
p2FaSXwvhseK7VtEaDiFSF5egcHFOVsZ26ra+Go6lDLksc4vE7tM7v5sZvbaxVP3oqnBimGTjvu5
/r1rc+0tAWPSmaZfMH6UTxaeUWaVrgCxUgFeITRLo598m0qdku1TyZgi+MHhsAa3BUHkc5p93AIj
PC6L5pVf4jWlpnzmAcRnWCRcI/39EFCCH3Lq0k24QJn8ftwdn3y6ffGcd2rwtai9/Obkm/LxAngw
mfp6nMgIoGBJqzt1Opf6c1bqt+rf5UVD3K8NkEuJ/HCwSJ86bvabsddab6StzcPk6ld8sIyeGYOM
SpAZRXabLV0QijkgRQcEW5MyP4rG5MF/fba/Uq9FxWHpZguhAItHydC3WI+RC/JUnteiQkfjk2/x
0//FM7hSWdQe3hI11Pv7sVAWX7zf5iM1vrwvncgY9iBjJILIKEMslLcNafDMSfRlGwhT3+6fdVOQ
Q1SrfNAxJWdFySUUUTJBN5O1KQZRGOad1pu5ZN8uV71O61cGmdS8kCebD6MIPw9QeH2xS53xrfrE
P8evg2PDqznvTo0OlON3s8+IskthG9pHjYyfra4XaDzfvauPlKOwwrKPkPTuwRss5jLqjtawHnS0
6fsyT4RjJMNxegcRjB33kvtBsc0oQypqlKdso62WNreG3OPpTBA8dvdTciJVXwrmnKykrOlIrqij
TJYxTtHvDLeXMSuDt20J/Q8+LTVZUQPO6xAqGTDrDIA5lyf/Wn+wgn4zg4N564Xm/M+dryfmrbCp
xjkhIr6Dr9ELx9XbML1SbqiOT93gVPqpp1LH0Ex4FR9LYvRGv6e7HQPRh9K9TgjkAwqpuKcrsAiT
Y60QVhCQmMlkCLMcHjDLNsdd2btZvPV4/xy+54poJkxvnJ7TymzUR10fl/vbU/EZ0BkCyx900kOQ
kZX2WYrOZ9weDpsHy0relk/4tBWw4DR6t6iEHV+GfabA9mbuqS0tYqbUouXq0fK3vmCu/P3JUrrg
1zkSosQ1DRQMeTRBoWnUXW7D3rSP4K3KN8u8SptUYWok6VCUxlLRU+obg1I1Mh3BVKFZg12aElKA
BGExsFbw2Vd/IJEaNX1sv04eVuC7Cic3m6Oxb4Ej+Nf/raf1G0yQNhWYGTtEKnhmi4fQt1aDRcES
0PyrPNRTaIjmRSuJLX85BkyC6w+wR7/pi4Zk4wz5DsxidJgrWEr5GEKEX9WFzJvpB/Rmch7UWvLN
xuzG3JOTvJbIWreDlv/B3l5m6D1sSnfoJViXtxD6PvApSUgbtdlUToNoPfmSF3dKObiMnGOs00x2
Cd6//A5czSIpaRvki96m1Ldjhho2qupPlz0qjMhqt4NsJaS4gpJBLIJ56U0+T1Xt7atD3DXz2C7c
RV90eLRXW6B/7KMLCr6iYbZj2TkVDcqp1snSqyDzxJ3xcjG5OuN4aRAISc/SbBZUal3DKOXFW6jt
ixiBbJwzfJQ/AxHsC9N2drv8fr2b135grKv/onpzzVILc3Uc5Uz0j8oOCvRF9RqQt8e5FaaAtbrF
3Hnn3Y3MldVkLbkJFTjdvHITzp62/CX66AJZ372Vc25TV0X3kagv24qrMcxeurcyWlBLG1D+yxhi
GtaHvYlf9Y7BafZrFojv1byhUU5NyFePETrfyq1fjlPFfwIgWeIDJchqUPQ9owBBPQEe+2K7PAvJ
HVz7gZL0kijgTrfo6cin84klJ1qQoZmX1TtdskXBiVb+9Mps7YH2J4uFSE83I+zTkZ7EYR3ePBhP
eBCwM715JFzBc17JG/xP/IJpqmmbhWQcAhDhN66I7W05gNTPc2mmB5Z6k7zf66Hzm18Kx/t5VcdH
5xnvGrBPH35pPAtV1ZkEF/zH7zE19qnauiWXyOtHWd3tNICVC/J1gDI+bn3T3g54q7FyzCovqfaq
1sxa8Fa5O91NT/qooK0XmpvFY9hH6ighdaUtjU5+zZWZW0krmZIz6ZQhOjk7IDsFz65IaV8B8q8I
+sxDYtFfcroVCP08Qj1DYniycOC36uScPozk22UpK4FR9763XbXc9dNiEs3Y9raQ2UV3S0fHMP6j
DU/X9jpcBbc+WJLbHDbQrlvxMJ3/7sf+Ir9rYWJEb57rEwDsPom8XBqMAXo1nGDgeDfvU7trCN25
jKdqcYE07ObTlbHQj/iGVKR2q7jeC2YUakPCjnO4eQL78ED+vrqvKgf8keq973MHN8lgDK4qMEcN
5TxXPCMoPmcRZodj5PLRJQtZgVxraQT9sVegCzXr3HymIAH8vdObFsGerdc/o/YiEnKQKfhKeTuT
tJbvdk9i0iGANTF4l46qjJGj3LEqU9EZXB+86hjVyhZIHD/7qbuiQEhuONDzodNUufkXKYvSo4Le
IAS+NYAn+OCRaad/x3SOQljOA7TsMjPDAp0H91HzWWVMEHCRJKxWtKmHLsM4Npx6h3TTcwIOyjck
WwYNxl/SDZu88TvjVJHPlafGq+nFwAnTqTTFG1e1cedFA9Jy0QKdorLbMze1a1D5ZazJXeQIIiCr
J9GCv/rnSlVfTBqBrFmkv3RSKstjo/CSOOEsQEBNUQUPPxq+giFsSh6K3V1Q1oFqW5AiVrzvcEnP
AbPMRPJ4Usba2AmJ9EARo148fzlKT1Czm+ZwPJ2ody4G1wqin9dyknJVioadY5c+0PgEpIpwZPjP
EA4VtcfcYzxnmoU/WiaVW+rg9ajSlcPdBXXfOjnIKvPQwCWFUnii7OfjFQqTcIO4QOS6EhSN86jB
kKr3rl1/dVHL/K4OCj9sY2jpd+HCkKbK+YmXtOv5/UEw2BXTMJdf1bwAMnR1j3OBF+FMbYXdi8JP
ZmSIrYWLrxObXK7p+DQBbq3hX37A9RS96bTHr+L6/XNCkeHz2+513wv5jVadEseodZw578F58m/F
AYkIpBDDMEH8ktSEPSJKXuVaFG5B+HwpUdkZfC0el4htBGbBzJ0PPeR+ztMlLiOtG1Zm9KzhUY2/
sd5uKXiq3FciSYpaNEkJYc7ycNfwMNQX4kPHnLbRlWEqjiJcZ1ffsQAqWMdHvG85N6DyjQaJ0m3C
tvgrVC+I6Y60I9dIdoHUQMT8xP7c8XMb+Ex//LEzsKPVc7UK/Dy8S5tK9I+SRS3suxaGs3WPGHRs
4mYT0/CcE3WDt6s/9JhCx+W0V75pK35V/eapDX1ou7Ogaa+iok6qDfxfSz9jyi/xHgQa/vCxan+S
fNv7lNVuTewUXTBkqPAzT4tkHBQZ7wicPioGC81SAUg2f/jSoyLULo3+g6LENp86HHjk7i+r0Zel
4KX7mmc8uKFn6R2MBE9xIZQshOBz5wv66eNPwpUGalw77Fm1ZQviAJ0NPJcSdEBczGGeET18tpVB
4lhwDl06yzmnRbEUKo/u69JENwUzZJSa4E4mjwHELW3RjEZJD2TY7V7kohqLBejQzziCEolL806a
IXeJTDDuhnvYzStTGqFKXhQoGFYebBTo8cm8ncmG/Z0MjIU/mYg5mYDn02LPKi0d7A3/7ZuBOKpm
NzpsspdHyZ6c+v/8iIPVxfFms9cI5Q56eGF00TAKaLbQZEfLxAHX6LDwPGVr/8YmcdvNCK78363C
NPZGyAIF841x3unxxnG7P6vb6A1/zIvOANwYLbY3ipb8kmYlMp2Fk5ZuGpCXQe5xaC0T6PH6nLW/
T/im6uiP3GM4L9QPdiBDhBXMoFiXjejkw2nmdEr+OrQIm1BmEp/AaJJ1qDaZ9zqS6WuKCC90uU5g
pUnW8G7rFGGjws3A6si25FbrTpk9/llpaksj1x1SYeqJQu72gGDgftiswReAKLdTi/JdgH+CCKGD
deb+SuMwJLJK1bhS1/87oZrVEgifTODRcV5GhSqLR6dHDvveWALJdf/OyUm8uykIP9rII/o0LmF6
9mOL4mN/vCVKOVfq2mLqYGu4Czay3mRbLQTW0jEXUsP/DNDkf+pmRboRXIFnYqjgWLj/9B2D8ENS
GLn1dhrwgLaRkNyJX3OzHNXo7Api2hyRewfH3U833B1OMcAlAPEFGpjfT0Xzb/xhDZZbgo8LKl/H
8hfyXvD1ssoGZs5U+jZ9+ScM9vrbhwAlJV/llu5fPY8SSXSY3oQokum635TeZfJsTWY9JXq/N2rw
SsSoNiEcQSsjPp8/nALlP+sVjgaGo4CRtcVL9iaTLqod3rM2KNO49E/EVL4ZormGjiq8cMy4+HIg
iFmtCLoF9yvCIECFyW7PbSAPZqdDoIuonF8nwHzMa6CXfNI9fZVwmJwG9giXQmkrFwGyxkQBMhXG
FRdr0kMLNaKf0L+kWhf1AFNmczOqpxa2CaR/jzys5XeZN+k9SbQRj1IMLvefFq/iVDBMmJ1GNjBL
OyIOxS5LwDj+pfezh7dgS8oaW09Ose/7g3AvpBdW5eDb4CmbtAMC/NZaxFQzil7tcPKNigDFs6e+
GOVScd+wpbiYeLzkOQCQVjmoTp7wow/5gkxWh0FhdQ+ejS5sYLrAGv0lnmwQNAeRkZhpUVsGss8u
TCzVc3HZTimdsFNT9RfOyYXtZSTWPV3DOUj9NTzHESYETsWooKZzuj+WH4yj3G4dhHmMtKN3R8mn
neeN6SfzTVEKWtBYxmLpJ99DtCNvcIR8q6VDMii/95ot60URh5XPlzW0aMFXPi8gnMygXmFkUigP
Ykr4JdhMdF6imN4IkngFsgpmeSCUBhQoTny80Wz3V3FFzhHRn/Kls5J1/mY45lPw1r+OWkzuYRSV
1alFQ6tkh/bIA/YQm/0IBlW5eVdQW8Y1w51qSwEUWBROeiBu5+YjWqPk/n/bsm0VqqwhRa48RX2u
1eOy4UNNqeBDYtwcfkZXZVgOD1nY4IENurpcOfB8DRqXJqlZFR98FEIxT+ZhmUmkL0B/jHt7JySG
X7Ni4U1n038RFvOd/wNQwUprGVaIz8EsX9peiHQ4JiCPCmuBRYkLc5WCgYok9jBM0JCCgL8prB0N
9DnR4y7n7KRqwtoVbY4uwBL0D/7YqxSDeRpk1H5E+QZXKkmXbq5FikR/xPqooi+9xn6vin7WrsM8
W/QNOvmPPPz554U5JZUZFPArXesy3HkNSbiEKDT59YBD41GaVZ8ycWQ3//sc7DSnKXc2aMKmPhi4
Ow5p/RFfQPaPC6/BnLkIl0tm7Hy+P8h/adTjZEyBQdmSeq1KWPQhGlndvHu63eE7v9gskZ8q2hxu
jUfDrU/YebX3Xf6ME1we7pEzb8BJHNNWIS8uSHm9x8ADx6H8LB/jQiyYhsUvQVZ1TnUIJ+cc+zgP
MuYOFcPu5WMFJ+VmDEhAo4cVL+ciSJXf1jD/O+SNpWdZlnKy2kuMwxwpFxldCH7JgGUAsPfI34Ma
BDSh9RHpgRRLYs1m1n3b2DySh16oa1n4uPLHHICdBqtMTvOUtX0QgqRb3nle6Tt35UHz6pdQ/xHh
1uxl1JVA9nijwi7aQvQP/OrOfh4MoBNbTYE3fGgBR/0q5EfvPzpIepTH7hg+H5G6de/CC1m2rB9G
1+lC4eQyf85ghOfrAs3UGfRBUTDga9ORAIhH7XxHnQL2MqMwCcmVfqdB2JlD3qJpVBZP/g9NNju8
ETLG2DUtTDqAz5yIQYr43DnPefeDZ7Fenwa4N6LN6qgsERZAgAAItWMSnOzROjs7SPcVlgMoF5Fg
CHGpL07LsvnNhF+2Vz4lqK3gBQCPvgpuWg+yIz1NsURcU4hKqurJmX3IBf4P7eZgpVbdMDa6RNnz
mae6ju9ZpfCrqyz+Rc/VQorTUypFqMndfUnKinXwRFnNFoC+26Pr2G+xGNPKBaiJMNflx5eNYh8m
orhBsvshinkRvVMMpyVdxZOeSyRHSlsB1XNNOcB6fcck8EkuzpD6cyanj9JJF76VOffeRpYoaRwu
UTimd22emuKdphMQQokPoFJKsvbceji9qHDagnnMsNRXaZReqRLpriREa6Uh6NCUw3FYFQL9pC9n
CXtpBgHsQzQ1tiil23gGV9tyAx9GyEcqOU49u1vW2v+wjUnZXNXL4x4g8rSphWLwBnFfnZ8b1RvO
JnvOZo8s9skwZ3nImlBiq7WpBbrl1mNYd6HOKOTQFIOeJbYDCZ9VjMw5VYSj6OsRyA73hhctIFZT
If/0BTw7gHBfxd50y3Km3K/eBE3hrmR2yzUgQQblne35lsfQA8sNgnJgSw5yd48PzPmceWF8cGfH
LKW0K/kbNJP/iGJSysNLLisZlrowiE0sf2cwj1g6UEC3szR2RmfRJ2Rn3LQXQ2v7CX3o9fMZnYTQ
0NVQYLRELZHDvRtZsRNK85iwOm1x6ShNhvxcpE9sIt6urUEAmoss63z+FWMKzee3vDK7SPLv9PM5
C8kRXg/Ya0zHgCE5o3PCe3wtVtX8dp+gkKo2t7WkjL2x/4qfihesj5JO6zQ0VD2QOAyj6IFtNo43
pv47YtMMvloTvnn1+SlRqtwvt/iFsHFVUvuco/f2gXg7P6wjfFLxsk3aUN2QHRgLQZ8grU/Teqjs
dgp1cc45Bn2Xvwk8+gLydAy4t5gr9Io4+Swr7vpWB6ENPX+rWtnWVJSd4Dbv++LZvGFGRCPkutBl
qzcpD1IcyFPKur7sfmHyLdZsV4OLwPbmZdwT7U7Brfl/gwIN4/i4MR00o6RFmc+POc0vYEJuz4Mi
5YLkAyGw4kWJJN9XmNWEABVsHogp487lwTQCWPJpfLzzotG63kAWiziom9xqckKIezj3MJQf1cnU
/nNHk2Rg+wQjUfIPXTS8NShw2TRetRguw3zBdY+q+mQmHprFU5yjMg2Z11lYYAbNpdusULFG3Lij
o+vUYkP7mi+viWrlFGpgh8u72eQgupRReopGXiQZQWoynRi7UQx0t8CByzJrfAdP/+Xr7GLS6awl
buIGxyfyQFP2cml5r45RKtN0KELMVbLXOeSv19okGo4t7EBOiq55sxK3N+MziVMP288PhiQtL2pJ
NOeY7dR0E69ukRa9zuvqLkOZ5y2k+/dNZ9QT4hkMapdHyek0x3SLBUvJ9djzQKneJJhLexlkBppM
cia0vf6ZbtgE9JmhIjlrASTv7FOJuJ0YCVMrhDw73hyrYlGBSRy2Pk3JBQcZ7bqGiqMbp1hQN0y+
BlBtI8pp7eXYLXOv/6pQuPQHLIeZCNuIXLER+TI0DtiVt45OlpqIius2m9mTqVQgCfyxtuUzMZP9
glqe3X5K+UCqNJf50P9Vr0TUVE9jRu2GptZWPCjamJMecSo1WclvSA2+CZ9qj3tn3KqiastFJ2z/
f/FF5TiQpX/xE0o05YAkjSGzbt2h2qzCmozR1CrXyLuQMyHeETL+b0ZYat5ttIVMXsYVgVSlAV0J
3+CeaKsPm3OSA9HTfkB/PyJ7lHxWcSikr+wiRdcfm1caMf1poPaVYCXDOCPt7s6AywV/I/Up5d4Q
F0gTMEAGU6T/SATH5JHB0Ew+z0MfY0dQFQi2ZEtYJVg6f6Uvax8OcO2Jt97FeMN5ez6slvbK/1/R
71efBXzw3qTCfSvHOlLt2NJFzPzkYvg37eLQ0YL/lO5lWxn0N0hK+4e1X4Ggzby7kay/4Qtup0C/
uTZIYgPpZC4Y5I7qVI7yWDOraY3XpGVq5dzVhJgwcL27SJeqZi+gX/v3PBsDiPk6YwHZT9wqgFsh
t5zYwhJx6JdBTSMUW86kX67uWISkDEzil5h8OPIvtN9lo0b2Wr7dDkRiBwOrcCy9X4fsBI+i+Tsm
WWoasw40k2t6TScoiWuN4yLY0+YzhaaVCLc/NXROd0ka8km7KAIkHuEBDMKIYU8vtfdOhgmAXQSO
1hsY6Oa1EHWeYo7wWxf/I64fU2Lki9VWJcRYtnUU8o5JPEg8nvJw6VCf0AQGCWXq9Z37G6mnbLUY
dpBAgAB901t6ne4wJpdsh6f1Z/dPfQPYw4Fbrq6/glsTFew8oChnPBnAr5i7GnDe3oER7Vpv4lmK
YQi4vlyM8EYBCyWOAfOfmqI2d4luZxuz8RfhMm/3CRaoQu7xT5XBRVpnxfWNPlyXM0l6YAvtSx9b
RRTciM3N5UbzeY1m1o2sG0rNfXDEOFm8N63DnhOT/qYz8SRdwtjI3mRC9jWA1FCirWH4oLlZAlOd
1HgjLkDld7ETtlX5QyL2YRH0i+e409/Zw9us/xlIibMHWQ3IIaHUamKVa+utWIG0isOM+DGbb5iz
vciG4++M3i+tK0pNQbZJXodBpnc16ohdn7adz3sS1s2+3/GfjOaFlZLAvp07RKm/ULp+EMDy1iNN
kRgRn5QQOAiQ+Tabj6mT0+Z/AbqIE0Wn1KYhlA6949zJ5eL3nAZOdpdz4Xb1V4DVgFsLpysuGIdp
c7+KgGLBf1BhAS02pJ1zye3itjdfkORg6qcTh5V6SwgJ1Ozpj6fsquFlWfS+vxiu0bGOduhUTVcc
v05w3cRdMfqm6WVNLDmx/NtLWB+UmLOZO4ORpqcKDuLgu6PlcQ7RT37w5XpA+itUSC2+0HyNlYwP
9a8WgI6D6LNqtyLulm+x/9bjMdMEM4Ec5ck5oQ4/+F2xYbX8k/KVdk6xmxWLHkK4EHQb1PqDvceh
JlVAevTEmJvDh4cK/75Nuo41il5qffDfQnRpefmjRRbyyndXtoui8pZWi3B9XMnjd5Gg4vv35IPt
DJkmIP2F+lrZwS/mOA8EphJGOabIZmNw3WcHNe9RE1jmDg5TRtBGMKiEPB6ckeulPj+fwwaguPH4
DOitoiwFg/QcO8irZ+CeDcLKaCOfm/SeO6otvephJJsEXhmIbawNH5DTfdvB9RX1Tl7oPAtYVDBp
j867fYsafii9MGA+6BoqmAIPguBo7SDv7RE7s2DKkURmlD6rt/HCZwMAlHK+EKXpyr6qD9QOBdom
0oq0dSk/sCyPwixp5XZBzF+9FJNrj+HOvnHWLzO0IDK6O8UbUoPc4ExyfDs+Vec8o4pU0LVeQxeM
05ldozyMnC+Rt2INcvMVHro3ytiBqvtJEffoXMNY8nFGs5uL3qT2ncaQJcECCps4s0k3ENxy7KDM
ceObn9SPkF1SUvT+h3GTNzwU1zVKspTfWPq+WnGD91npUS5daCOzH/V1QkYvDLK/2Teui9QXXERm
t9g39RwzLWfENw5YFB4FWg/f4UnEeH7dhLVDucdXiK3caE0zpZDCv1FL8o69MMbn8iIqdyEcJVYP
9eMEpt06GhSwFMA66nrwmrPxZyKZq1Sf65k7CSiWRYxuD6/3ocgRS4aSdM2Uraw262q9d8KBHsMm
b/U+yaZkXsDppNvcVOiuqCk8b3r2TccHK1Thtnxi0icuBjVyEVXz1/gTfwO14i4EFacZS/QTHp3t
i5WmVF04sCWM0wzXqWgXxGcSun6ZCFNTHx7SoxApACv3rjJlwZndGKfT2WMEA0pvCuMTl5wiWypX
GVpi9b2SZASrCoousRQrPm0U91b46O7w0hxpmcJZRuFqeoVjY+B5yCyZcpwAERRa0ffrM397+d57
U+FB2p9AI7A1Mo9NoAADiM/VKV58NIg7ROtjSe1Famxdz5O7HtFCyDmync6KgB7RmWx67ny+vqLe
ra0Rcl0ksPoKddRCIrMzyzXUfiG2Oj1pmh2b15flRHHuKmmW+uh2L5oG61x0I0UutAuEqngG+/Ln
FPQZDi2/WtDiy3BTbvGDfcvqdxbRhlrkSRh9YzPrG29I/zh+D955yDyvTGfsZDL7cUd9K847QaBS
74fX4rduS32eQtng2RFR0TdvkCR6FDrCzB0y3ML/tT6Osz/cNNfhKY8zZ3Npg6V4sIgGThO56uWz
dJ1ZTGO3wRt0BQl8oJmsLZCGrkXfcpm2Aa3brbkmr/WU3rzaa2+3e/oGLG5oQAEqYTQTaaoNdN13
T3qgwbQ10+Yy4im+sUNlsaCoq6/mo/PlT5yJJ05hla4TgzlNTqyY64mhLGSAmMduH5IYCNm45Xg8
GgEGu/hl6IYWU62t24HuoGqMo79bXGkpylfDfJJuWht1p7zmzcWZcLA8aJXmer+WZJlhkrknt6F2
UXuQOqgm9AbRzeblDW5WimzxVLmmghYBaOpwKhtx9xUv2Lfxux5B3CCIjNKvPslYi5xPMl04F8CL
5/itKy3yyZsDRwCGojbgWvorTzsPv3vAdxC1ds3FWbp6oRZ5mTzESAYeEtCCheJPlIjSAOU96NX+
NBRP+lYMLqkcZMGKALWIt+cBQn8XIWOTlxYzfAmDFHzLZ7mXUJ0DYmT/QkurjkYJYS2A/wZjiUYA
ejxFnDxuCJg6J6R1Psrc9gG9q3pZqLUrgsjN2/SmLSSawYwifqHlmXAsT8lWOZLFRlcGIOn6I0ed
U+/KOB/bRL1ZUqXmrTN4787AahU5eXYU/9p22WJ7DiNKW0OVnzLg2FNDjyQiShy8dc2F6IPppkHC
WD1JA97mYJcK2DzV0L9/SlhJWX2gzDJLAxpVRUonw7/15220CmcZLmYI57gGvb57SkN8Uqz50klZ
Qpp0jkwD7M7Sij1fB/PQsuTuB1WiHXU3vNouDcflUiDSlQN+U7FTcplZffvY5DG7w1QnP4OkfMgi
xScpIl8MZQn6BUgYgXtjUcfSnlVl/WeLtr6x+0o9B8MTOU1RcJWfkzjEiGZafdklUBp52bOYkx6K
ApLEstYUNKaND76tH/dvXSo83d6Dnv2dfBu3AdgwKUwDLLfJxSg/v/asMo5SOvZ7iOxTss+mwPiM
StZ8DXP+1CXzX81RP8qez+r4y88D4GmcskL50gDJ+jjeehrBTr99XwHWA41Z1u6f4kCt0qxYb8Ha
6H8NUjC5bAO0bXgwSJPyXxBUAbfS+5MWKQV66tcz4pgQEIs2EC1bqdLfwMy/Y5K4dt6cOpLTH5rl
DxHprvCNwftB4VF+9S0oKt17QgQOrS48RrAys4v0SbdlEd8PIjZY7hPH0gtvhcIIqIX1WNe+CrAS
1R5a56rKihfGamDIizG9+qHji1TYVQ8UDohJ7ggCJkI4koCNHTX8db8fOBo6eFvE29XhWAsoL9Pu
7z3wl0hgkE/jEfljGRQ7JrtI1vfA4N4/zPAvJtxui1yiUDRhoHpl6okD9akKubOc1b99XPkiWtw6
8hXmRhD+tgR5assTB6nQYMwCy9CddetXaI2PbsaWZq+JNZ/bnLRlHQNK0dz27S7cU7+07vpVXCq+
txtfNUSXptHqUuXiqQa+ekuj1L+5T4Ads7fBaaFJ/48FR3gqrzMsJi4l3rI4V3HJzvFDPqI/6Qma
AHZ4O4tuukQwZy70EW+cBoUNeE0nqE3joOPZukJik2MhEBscIYgCa8xofYFWs6EViF6pjDAnB/YS
ppfenFI3BdFEV8l5m545WgYM3vrbzp5Oy1n5lo3vL15RW9Yr+jXGeqPGM+Xjo2F9WG8xOamLuH+C
rHfr9Aw0byyl+iAUYJfKYtJlLfXfCJcAwV0y9UKCWT1wJzA2IiFvgK1pk2lNJRLMZWoOsUGT2v3M
HoFgDWZow1zXqkgT2w8XU46bdlN051yL+Bxm1/pmfQk2byDzVmnvWVBtsV9Bf0YyvrPiH7ur6Tn/
TaJdshX1lNNIOEfVB4wTtUlVzBe0bTds/gbCgriuCYVxCi480//XHGlfwfeqT+uEfH6hZigKrO+Y
UR0Rv2ZvNUgVKuUFn+nWZelOeFb91PmLhviv1ihZnsBhpaLRGmt3D0AYaNQ4TOigfqSxEM8woAgJ
Q3+PoJmFiPEOAI+0Oi+3RaQ2tVYLHNkmx1NHWhsfXbSKlpZOP9NU8Wq4UUTQ14NZReUEXrGSuOnA
361kne2eILz9/onBsBYaegMm9xeI939pJz7Q3hLo5p3JkOaeopl71GFDsc7Xf+O2gih4Bk1Qftbd
l9Nh4wfARUEh+6gxistTqPZ1g9EgzbiAF7p0cV5v64ukTmLkvyo+4BGcVBuVB+lhSLqPjXnWktGe
NOGUz3MIvzDDVk+OHEiq1XgJg/1XNCKMI1YFdVS23qSOD61wlmkQVX/pgwHuvdwppWvlpcG6YLKU
5NtwHAE4kqUZMTaEIzZquYQpSU5WnY5pdAQlLLQeNQc0te4zAxpx4KQ3yboNtXF4NFQL4exftSfq
PrWIhoJzwNH+8kAvQtGa7cNN4XOzhvIv9M4J2IWvUOwHcYInokFeZ5+zMZiUzN3gttxTUpSAqTsH
fhUwbRJrNJhh3KbYq5fKCO1Xqx8Zegp2VX2eGDfF/XqSWVOwaRpwlJZxt7h1wvaFTu8FBEoSRn3z
bKGOboxQwN2+6G5qhpIBNAyzOHwwdQ/i8QkHI9Jgl5Sf5WibbiHiq/sCPGRqiaw+gFHKmLOW9L/D
TRTARD1lFsrkMQFYagaKlEDOfuAFsS84tCsuSIb1BujTBn61HCZ0bST5xOtnOOj0NJOe0LNlt/qO
U/bfr7NzkGODWXq1PVqX7zWnHcNngQafyaHCgejuulI+xervqzImd7Md6c5hFhCo/VUgN3qVwgmY
WCLXaliZBhx3w8uIDuTaxhtEC6GVkxWIw6UAkxBQXODTx5mvsIUaY7ED+SBZ4obNW6dtHSp754xT
00OAj3rmussnh9eLjaGZmRSpE47Kw7M5OpCq6dGLZmh3hRDHxBEiHjCR7gzo2bw7gsL3OzT5BWhK
r7YZbAPSTu6BvJ0aEingEgWoM4XfacEoRd2kNzG1yNRSUnpViIsIeUnAVdF/oBkK8u3az5HKA4SM
oiZWdHnydqt3X6Oz3BJx7Kt+b2gKr/FVEP0I/2woz2bVoyyv74LPke0s6qp56v8ZLG/MMtbfuzsq
byMTosGilAUrd27bt3HTvWFUL8JW813yPmQPHzXrMIpBau0UqbQcn1NqPhqxlHCQuCPKZm4Ju6IV
TDmM/VINB7rwbJHd6311tk12VYF+/6bgUyAnUurLVW3jWE9UIBkFRW3E9u6o5qKadlb1OT5DGzbf
A+/Eox4q9qsZrSEsmXrAIGZBwdls3rSEbFJ3jZFQPVj5Ojs9wmxMICHvD34bwIw/DPr8et/88zsv
PkdhqBQWPsWTczKIW+J77It8bazAvadMOlmvrzJlu+G6PK3s03XvphCZZmegV3m6CB0kFHc2S4sL
iRIt6pkIs1Xe6vJ6LTtn2bDmxgl0QhfxhbdKJIoc6vElc7+R0LAKhRXNI83jDX//uXybHeTaEUdp
fnS2uE/agqzg0H3EsEX8QIHaaQbhvtngZ9PiEs0TrgC7XeffPYL9SitiBLUBsTPL6L/UtBRsT2qu
Vnngj+MJI+lp6qxdsz1QkdE+siDHpQkbjZlsoCzJyiLpOL1BmSOjsYEVh1vfI2y0CovaJxx1dZ/G
7c/q/QOr2TcP53ftRToTYJvXeKrvzWm5u99E9WFvB80Z7OX4NAGTvOKfyLcgiCE9RXTRd9yEi90i
+PWYaxQwVitxi89xqmyFOSw0UZAJ+B8SXcI+iXeyuKC7SaGVaQlVylievd9grng60yklbJHwW1A1
vf+M3MuMAfByy4+OdwKJwDuAokxQl7cTyfrwdOG9OYCsouGFREH5d7STIXzE/hx6rwNIyjmjAdBb
kxiuxboLZYtWHegoorld6EZgrAXI3bRykY6km3BoGzWzqzUUz6NTzL5hKuKsHFHBZdkHtMAOSYqS
cTGqp7XlbuF4l/tUZENkRYc8/GbxYUwiib80R05JpvD0EADcJ54FaHayH/UM40k+ZVf32hZGXzVR
KJa+tTbJzx3m8B3YDOeM1UrEVVUBkYrfvNgpzTZ6A8ecSbT65osafFR+Mn/YLT+BEsnUnYIugSec
XLhVQdAfSuPq1PJN7zX+J2gBasreXApZ2yy86srA+G58Y4wwoLqQr8KYKkJ9DXplJ8JgqCp9+UFW
Jud4VPZ0ZlIekOQYFTFsMtBVXq1EMuIVnTrXX4FwlRcoQQ2D08VPiv/kPQRhpfNfimELnIPHwI7i
vFaCwORXNP3f3wDAjiCACvc9QdngEkEwjwwS9E1CRG8F+FzMEzWLkvVSlqhklRg9qFtXPDZfI5lf
iS+UTVort4nMcd9mXEd9UrwGPjWpfcVUownzyoeoo3Fqhqp6yeabII34hFqUS6x0A4HS+NKdheNy
vittYQmjcO2avYhxZwFDwu2jTzS5pb+mvSb3MU+E0QLvdDVcDQNXK6uszrOrN4Y6a8tlzKdjsGgD
2gpiC09aBX6fGBFNOfiBe9ycbKZgIcmzGEr9JncVmP+bbGNOMbMuc2/8//tbKQMDwdOGLnQQZybB
/CmKQS376uF5Jh/yUSU15e1z37KgLeaHYErBqwvSrqYhV62QNdrRZR0pJl9yi4H/itOlITv/1xr4
XX5YII9H6cMLe2R3q/4XtYTmf3n7pLTs//Bcp2a1YsKmoRPugrw8u5svfg6qE44i7vojBMzZT5BO
gqRozowF1+wfcYlWJQIxuq1fLP3IyzD4NEpDlJgPG0Xl67Hd93AYgXLg2IXh3YH+PztvmvPErqmU
EKFbtB7yi7BsEARdrm1cZySVQkYJ43WV7zJSKTAW7Zzlkl3+uno18PuxrrmY/P/jMOmbTvJrMZJo
PcyCtzLRJSuNSIbb+2/4/q5c1czyNIkEnxk8EjynwNR8aqOpjaP0QYPuljaBvQcI46beMhD4RVO2
JfuuUA/ge1bM68kKdFj7zfJO7vzM1cGG5Cs10KJE9B7H7PWLXTXxf4W0o6A66Cz0SVUg02jleW2i
xiDjKyrA4sLi+xKM3teRwow3z9NQyJ4sgtG5AMERDigyIdGIL6UUG0T9ZHV4+497DaUeBNEnXItz
JcvaCIICwfa9yupS/XIO5Yce6wgDsdbmyatm4KuI1OjTfFwuBY1VakjUexzqgJPg6c2yEt9udeK0
JLHKl8/DbJw4mMmiCS/hQV5n1T2tqjl2WXIWhZhLChj8Xu7njzvpQHEAN1DK2exn56sx2/L3rQ8e
SddsWYLrHkopARKmK53yMOn5gEi8So3/QtfwUGAQKvSxQ9lvci8olsni9sPdWC0QfEeHksrYP7av
ntJa1D1qV6GIJG9CL2GcWFaBAfAA+COVMs6wFXvTW+u9cXhyDPu4DOPX7NV0LK38Rpfzs+acMXqq
bSMBSeRLPt9DhfSJ3KItKI/nn0aQWG1vebgIH9tZ5OvtwOVgXptSQGbUWEfkZ0PDXjGfOghi/1tC
tRBqBRk4bS8jRYR8Jq25bsuaP+ri0HmwtRFVAtJYiCLMYs01uBQMf6BRD+K5nTmr0oKBwai8EgMH
ZfWnVS7X4l9Iz0m30VdRodN3LOiOy2dgyBT0/iFDknoX8Ipim46qXc6h2bPjSUFYJZeDD7kRP9lL
tztoV8fyRnqDQwHnxeeaWKj4jtVztEwKpdOAqwsqXmGPSn8RaWAwrY9CRJSf0KDPVOqQYGGrLozy
G1BY0c69+LPdRIUrDroQGT1MhqPhojDM9ZuSDPeXimSLbQCHt/FEhWZWZdMbRcjW6knYmYF7rRUA
bfynlnowMwfTzYuPXPTAIK6LQ34/z0qyg9zFtdUu7DWrxG3iK2tSh7QhDBXwTQMQHmj/1LEAGFFQ
69UubrEem/4iRCTafNRZJmxYwA/3jB/j6OvsWHN0Uhx/ltEDlGDNpU+BFFU792n4tDOmdfj/vrYz
lHwLNYG4y4Yb0gx2NnjHTX1nQpdHOPLqSqdiqipLiuLeqj4F8DaBU0QRwHfWtxhOpITr3apobw74
68qmWbvQp2T/0baBSTIC26/95UHWS1JKe7IO9joaK8Q3/VP0tONFARGMYatSkoUit1gCwQeGtI5D
i6ZqyXH3AY/nbt1IygBEssKnEsAuN69w6K6FD7ehAKwaiyr4ZLbpJo0YWGFfelQPf7BRE3nnF6Ia
3bvRxk/HKiacrwCal8m23s+NBCLiNB8ckaEMTUjMgovp/Ym51Pm+sHwmH8VEvf9MUHmSEHOFeqYL
4cNrJgcBEiMD/wSIOQ1I82Ywp54ckXynYllbJFAunbiHSMRR6GSHelKFAsuwiQKuE34csFo1f/mg
d/GY8qLuNGSvYbHmI7k2Jqrbjrrseu0JGyXYCaxFYZKHTU2kbulCATWpZyzcUrP8dZTPcl+pzN3i
ShjIRkQfW+eU84YRnKLMhxwGKOnDcvocGS6MbmXOGV+jgInj2hQDXBCbZc9Ne/m04MX3jWB9AOlx
BB8aIgXnY4gkwiUaFS2nCRskgR+P1dKo/Wy9VTnG1NitZHiQZqO9AVX0X5WNu//SGqrPvZrAYRo7
jKoDKV6piDAK1uPSRHNXBcaxr6SfiPizxNvym6hg/XG9c729wKtRkRh76oFwcDOzi7UyPdc6Lfyg
TNGXEWKpZScKAYwmWutjtwwnAgew5FO0kUMmjUDU1LKz+oLvtAWG5uauQfj3UN5xg0EcCyykPP8e
yqnW077C9xY6q7HTiMNKo0MjWe7EA6xx8wpkj3aqKkFNkV/Irj0fG5Vb/YVvWzbbdhVuGNjKf1TW
PTsIkrE/6IBEyOhtgS6cUPA4HVgYGXnWCOTtAI+xZvVrfewUyhSR5hMUVisUOjXtiP7G0h8Rninf
UmLaBTfv/SMeqqvHd4ySVZ770XKkuedEBQXL3Z82frXl64gG+fhTGEjaqY2OtoxxWvI2pGWPe/iT
Cv/JdZtD9gHGOH84cKk4QqKRmnXmOQKAT8dLNIO/WwtjnCcKKylAoYN0zFEnjM78o/+OYcONUp7x
FOWmqifF/WqNa6FU/ILLvHbdqn8q9UukwcKPt1cOQu8I045XJp7K5w9bv46JCC2OJJxCwV5uBxzj
KGjfwqBCJYSswH+TIpcCqx4Gub4bN88cFfZCsZnFFh4BYldVrL9y2SEmeXXvf4zqOiUV2uqRa5LL
ar+MTTI4gGkWkAAQNeoL7AAfFRhrCriSDAgDmkoN7AD6KbHt3PvdC3u4Ni1QFQqCWPL4XLxr6sP/
kK+iUoB/UgWlFtymbXIU08UK+qys6iU+QBqpQbI0bAR74rYjOBuHSvhNM6MHjkP4iLe5GOMGEFEq
yMkVrb8mEI1/aMfPxeeIIsQiSFj5yNZdn0r9vGHh2uSIml8vFQUO0069KWc4grIyAL30Z3gtwG1K
SjTcskIw0LaS4snRtEVC/CE8Brxpttk6U1IcWw2X061ppbPRXpohyT9dniVnhvfYDRg7hl/rqn4E
s5fVyhB2o2f+FyuCqIDaoS9wxejNWavDVMMylsXR9F9SlMYWbc+HaGJjh7GBA0z6hC39yEDkRFNj
ddRI/9oNSCrFZG+qPmleNtzPvv8254Gn8c50OxDpBjX9DowTjl11VSNC0Nfx9JI7H0PCp704fehs
grqyDBm2Ze3ItlvL7HnHmGameSP7vjELdSMgT11AlHW0F0xt6JnbVVqKbPORfvMj1AvpMpQ2Kk2m
5V0/R5ci4Eoht+FDUS5pNhD5E2iVHefLJ+8IvKIW1NVpCqml+9WWBxb8BMnL48tYX7mecLRSauOk
0p4u0bTVCffFWeAJoJzkSWJ4SqJGjhJEwBMmWJ3pb+Kevygx6khex2piiVPe7yNz3K4TsN9++w8U
Vy4WUPtDc4O70JGEzud9MJNK6PCePW7SRI9kXb46jgCcuvP3Anzi9NRhGbw48ND/46evsr00mTWn
/cd9A7ACaDVQ4wNMRDxUA/pZI2u3FE3Gp47hCSOT6AEtsPJCDJ9WKgGDuTGTnF6Hr19qDOPE+a0r
JAqPT8cttxRGa0f0jeil8UGuEfsWGsZTaHBXgNtm+gZRsOoYZCVMwOpWSmuXRUNF/mCCdc683uRN
42wGnke8KX7w7etwVR2WYgJ10OPPdaDk2clK7XYdov5ehB/64CEJg/Go6KTkAFssqJszf4Q8BtHT
izhFLAJGSEkj09eGWHm0d4+N25ZUiyrOg5vXgSupp3B0oY+EhtqkbPbhL1I+plE+izP8Xgb6Ar4N
npiuu1AW0YgMg8vjdggYSxYs4undj3EgdPb9OucwjpnB1a+DMZyFlpyHEr2XK5x0z5S+8r/TBjEb
PNGxowXD6eSHBs+sd7uMbtaTsZGQP9TMdyhqr+eIWKrqhb7V6tgIg6TaOXdjGVZbShYYEnwBkONs
jjneHyA5oAGWf/tngoH4dwv+smxP5HgXgnv1qYcf/k87QkwWI6iC08RmqmBuquUqRSq9p+89oRKg
LhB/U8MtANE/0KEunj2AuXyuiOkbdmBtnRAHl48q2xlrpFyHxaKvctcF4C2Q2K3wxqXXsvr+XuKg
Am6D0xFtSd1JS55nw0tZvkp4WqbzIlHrve+kn0MRl+UmV0v30nzRYvIUzscGA9vsuhdzjDdGc5Sg
3iMpshcUwO7186YoPHCy853GEb2KrUpe9CQMpLeFPvitFiJXKHZC0Billv8+u+ynjo6xaoGdh28/
YLWBzNiZdcknhaFKGqu2puJ0aLUUtlLbABFf9Fd3yeOvn8G6nrU4vGMtCzMocsCvnUQOXIcAu3XO
BcIJcH6K5NGq9Q8fKjazE4eA4qYhEwfrm3h2JwB3X3KgE3Z4Jrdectv2mmBJQ9KluANhyUnHTsHx
PSjgugFpXkjsn7WSFleU2dR+aR9FgkTVHMUJSp4m7vC0UeSEsZl7ZKdz4/zO3wGYt7KcthSOfQB6
PVcSyyNVS5sZT4U5yLsnFkrK8LdGBjZzQCjk2vc/01AE1aQTRAbr9Z2YDoHUwFXBBNr+OSj55cAj
iK6qQE02Rllj96S1SCgmmdQfj6sc9q4tCKHffsDFv5kbHny2JswpSvo1cj/hiS4BgdmYhPCVooPi
C8k2QEXdP5nsEnm8+y4uF9OMxfu4CIfpqbQFzPIyn5sLKRmuBaUaII5CjtqY2PwB2Y9ghEen2lsc
q/ZP2DXe71uyI/4y2JKSrAxL3HY38f7isLtiX+bnuhplO6pFojbbH3gVQNFoyMVW/siuIIEW80DY
zZs3THIFhf4sR2RUwdaVGFD0n9cXTN4Z3xngITO8RrCmky+LIwA2S6/wkQJ3E28Q8FyB2zNep9kB
A42rJNw0Zwgq8RhAF7CTq343lGxLHArL2mC75Dt7T5pF8yXiPr6XEki512cVzfoNIm6h+z46RZS3
xw5hyysk3sJVVWHcjtgSTh6Zw9kJZ8pJDYrnFwL81LINVrY37I8QodYVc2BqokDITBkuc82fu+rY
rdD2+w/O3AfYG3lCp2XuVo26+vmKZ4LwtH6ToALqd5u5MoRbMDMbVci48XN7BsS9k2p4XBY3tECY
MZtkQSCDhWwswetpVZftFKcUSLfYlIqcQyGXk+3ysRRg36ohXk7X8/w1oNY8ZC+qcZit/M253JE0
bV3aLyc/gphw9enN+4J6es9tLap1khMIbL/laC7uXdPCoyL+cBdYidTFkVTgXeDAdrvyXzRyln0o
MBPsGFM0vf4ZW0JedzlabBw+tLEyS/nGw82GAos3Vg+SFlhd4fGFSRIAa0GXYFiSvCWGBeHoQ/WH
zSiurZer90RIIimbv78klq1he1jTg4y5+XsPr2CW9eyOMZVB++d8x8xIQ1TJUVe3niuPifFr0KQc
PqJ1BifGb3vHMaPVA2esPCQGW8fm6Y08GXncw5NE60331zSpD5gpgiHIU2cYERE4pqDRttBBL0w/
/1EPmYC5VV6KITNV4E0xQ92ZPrx9rtjpr+eeDbLsFj8UcO66kdK4YylVLSiiqZbNFLIge1cTIKEM
cSPZTVhuplrCn9HjW+tnOUcf7tdvstiwtmyqMm9gZePzhbDo+RmPRpRdt9JgLtSPaK7JAn5Q220g
xsar2WgPxj9oi0MQKaqNAFy8xCmOmgDS/VyzN/JINjwj70JZcEsaNDiRbgoh0yMweGdJkuhg09ju
24BqhkfKcNfqseWthoJxJFl5tXp5U9xt+kElbXSmWu67L6dK+YLwhf25OeD3205D6RfNnJO2Fn4N
8zYG1eML+Egtjt/VSVfj5k6I3Cd9q02M44k34lDXg/cGhaIqWNAHIcShumYSufIIq7YLDVLtuhbf
BKWXr0YBj7nu1HhuM7fTSzJXQcAGfx1xUSww1GBdo2ibIqtodWDL77Nciz2/0lvr/ZQjNKrpseZY
UmKfhIWxMTAUJzqKBu8jDpQXMd4T74lOyGQNZDPhdKFyl9Zga8tQd0M25hNyz1YCxwDC6nG3hjUc
lVkDRq2/svijaaliN248TryJuzbBtiFEEzwSepDHG2uCQoFYfg83kXPGBbykLw92/n5uKybOPeE2
HCHvmz+xpR7qgd/7iTdocvN3lBsDJiA+DWUdnfbRKmcYg47VwVltx2ksmg4r0dgKgz/HLWPfsqGW
NUkYYPffJn/EsG8jZ7zRJxoj9udvlpiUv//fis9a8QS4N8F7pMUgYoNXzIaOIUQa0AFX6fG/hxN7
nXHLjkpmtP9Wp+liirCKzoXRXE1vD6isM+hxOToXkE+3f7YY/ngO2LkZ28URkzr0r6t/jUDXorFx
449UXG1uVR0mKc25M/7RycAqLw9Nm3uf6IXlYDGX59d7nPR9DWBTzwjX5ZsE8B3+WLIf7kKsIgm9
Xq7VzZWeMO8n8GT+YbcCooGnSDJMz/Xe9AIJxn5G5UpsBDPeXzHCnrFtKSgB+V6Zq1LKuGsvpZ8B
C1GSjXf7qcIHESVnpGRB4KinULYuh5ENaLmnrFOScv1tu9GBNk6IEceHAi6pYxE1Yxj+wEWMV+2m
DmALxvuQqXbR+BcVq+Y1q3Qj+5KsgO6tGvza87v84n3yyACrLdN+Lcs72HpVlu3EIUWsL0O7t3T2
TUfd2ojybsbt00Wn6+aqVXD7f3StuG6Y0R/BAFb7Mu47D2encOAj8OPfft6DB7/VJuN/iWNlYWx1
Qwt9jo74zHSp0YcQywIvofBK9N3j/Zke/pEXmiUQIZ4OjxVRvwo/x72em/B2PPiNVfZ2GmrBgx5e
r75KBRHhJ4S4DFRb3nCX1BBV3Kc6U97ns7rr9XtLzSZy/YZso+6ctimOYWe4eRTlfqNfD5pVgTM2
vcgKNasP7di5UeszJli/yU4HHCE1dwHCLeaYwvsIvOwcn8iTNFKKmv/dNc8+vRaUNNrv6+loM7cU
j++OlLdyfIVRTTYXnHmXwpDq7mt9aBb3w5CmWnny8R+z9PVZvqv1UkXEOlIud7vOK2YbHXRlOeBs
y1vLH0xi1zHGhhR+4W4guAjtxh0Z3OgGiZpqytNpOwagLajVdaPZLNi7LwBFPegWC32p+XkjfNSD
6E6fJISprtPCWMtxMdN9PQO28/dibjIYyI6Z5Ddt3g8j5bjRE2rWWehBxPHRMCk18rQrMQ8KalZo
LMrWwmcSAbk1GmIaHgfOxTdzKRVZzM0FxZMiqYyxrvq+eNYNb9r5qdjr9H7Y1142g8YbdVPoQT+w
MvUTYGD/43EZK9jSnYPDZEQ+RaUTLXA3qm1NQz5IkTH8O0PXgk1fI3UvcN2+O2/Gd1jlFqwiolVN
tccoEKwbQQxD/KBIuYDE2rm0eQ9YBhRSzguiFZmSGI67KKlcFM0A0RP7ZQw4vdcwJtpiTH7u+5z6
KF5QDJqVxbFSzBkiJdYQ0Uq5xMj1DcpA9ZyutJ0QZxvFrJRnMbvTTg7KiEi/LMMvriPbH9lDIPof
9L3CFY9IDl6uugDxWvcDbXiu1r6sKKJfFH5j7OF6E8w8TooxoolqdjlL+VPwUSKT1S9m3OvZATrM
cnxq817k0J3enxQs04Nxd8wFv0y6PmuB8KJWf2T6x8dFs2hvluqcN/4GYYdmm/pBw3uZsgF662r2
LrkAjn5eMez1V/edLtYZm8rI18bix2fXax6m5YQ/FvFazmDeJwgZxstAA1A1lzcfXkcMKCs1snQ+
1Y7zzExSYErMl9rsB0jI0c4ThZUHKod9zbZC6Gsa3wHI6K4jLtTSPH16WptCBaAkznzdnfjVQSDn
+3IEm0VmzZl7bxg42U7mdGdSbSga5QdIsjj7nIA66Og6kBu9MQ9/H/YE1pKYtlkkimlS5YsntPlH
F+XF/q7oPA+FDuF1yv/DHFQDD1uogIBIqGEf1CgNVjgOfk2gOU7Le+CCnNj2oFiSn8ar4Wj15XIJ
0u/BZ62s6w3tMI+q/X3eXXVTjMMsVNRMkCt4WdNRnRHBumi/yfrnysnBPOHzB97MxGW2Ji2yOjam
emo9n1rtPuAjkjqwoVBsGOjLJE078PuEjMNlKFaJobyfBRUEHIuZ6LMAUQFrmRmurCCVSEVxTnj+
EYzWQlwWoGkx17/YA+DNR2ZuxFJ4ytpkF0w2fK2PlutwgtOJOpUJtfWyTcFV7r+9MLE+zLMl/1tQ
j4O5KbHSEZ677ajbKkFZ96PiYcbJjuZmUQIkZxHoJkYxgczfYnog/15mvOj47MNaCYvealsMbc0U
3xd9m7+MbtLvW66sjqYV2nVHhb2DMN6hzTreh/1ebFSVZMM/6zeAgCnRsxqcAqXKgT0hjV5tjIe8
Nyy5kmIUvXEYZpJhAi5HYN1tc//1vM/b3DOY2styzTgv2r7/qFHVOVlM86VCXIYBonBjZS/lhbbz
8x/uNikhIy91erRktpmDlWZwGsrSUWYUXmNBBrDMCVpWHnuo7wz2qD0UJR30SQ8P/sXtRoBHyjPM
qRZWPC9ZMCl6McBOw8+w++1Rj3BySF1TukG1U++RW1JZTG5gaj93+4T+4QO5K/G3VdKSTeWq1m8d
F5Kn7wJ5l8wYRuuf2CH49Uy4b5x1wIKf5qLZmIi0cP/p16dWcJgYcUuWoGM1qABfPLEnVofVgvGd
SAkexytxvcPFccoOWDg3fxVP0us6druBCqmmfZlNjgZdoy58M3OjJhov7FiiaxWJWHPjfWkOz5Wg
+WoWPBlY21Aqo6fKaDVkmebPH3mzzzOAjEOPWQoXVvMsd6WYDfMJROQQw5nYLP7RszgS4KeH6BTq
i50qenv7SI60umHo9WPuL4Ko5JbSOfhs47agJ1ahYDhgC2KpQHk4peMA5/FL12Wiziu/xpUGnlSK
1YcrJnFXmIY9vL9i9mS9Fvhy9IprC9b+s/1Zg34LPVBgoHZasM1HNGYO3w8Yz3KSqv3/VwESr3BY
udCSPCUnTXPRD9xnvveKrag06vXR9LToeT553IhTEUtJ2ubnXs2coCPVNoFkrG0wjGB0miYZww3k
40RnLst/EFhrIx6Dm0yeYL+usyFvWU0bBH+6hpHyPzjqsvEur7rhssQd3wnP2rTwlFp4+liDJ1Cp
hcZotu7cTfHinziDf+ofyunKX5SLndLt4A3YTKXd4PwYW6lZVoVuJDEYI0DERf7MleHneNEynD/j
JWEqLJ1oxLa58QtLoukDTLPKDPUkwh81kpqlfhM8H0wkPCgxiTjbNAbH+KHPqgZpQ+g/QgueC7eC
2FyAMHmhMpz/kvSY8pQIWPJw7LWp6qn6hCxPQ+KczouMKTYSF7zTScoqge8/6CVYR42vOA05KIzM
f7/T3XnHg/dYK4xbl3LuPHecFuFgl5lCYaSyqfd/oq+STkuJ7M4WxAuP2rwz9uk2mK7J00g4KsXn
239Nr6578oxWsyY2YpNMU1zEBehuhINVuKvhMYrRomYQ5CCLANPv7GMU5jwzEN5W5VABKsKXN9XC
gAzX2v1HhQZuGVc6jZJSuC0hy4P4b+qIPuFP25daWI5alqbRhir2e4fJv9cTVagXgMps3XU/iavg
FlKK0GETQRDJvy4d5t1bN11CxJa/UWZUIQwnhFQ9MEA7Lp/Hr8ZXjP+yageb3C979K/PhSBZNPoG
J0I0y6JhEcF1cHvwe4EU7y60H3bTKS9CWy40VTsqcR6y2ZngGk9Dlj4QNVrWLs9F/Dr+IhaYKsr/
9gEJfganWQuHFst9Xdt9KChiHL/eudZ9Ga3DOLERYLeJLqiUkjE0lsB4PUUxJoED7eRX+vfzwkyF
o+QiYz/STQIaK59bdOg9a1T7bTlB/GBmcOZQdRnHfcocHAc6/JTC3yQRHqmtCjbN+skt3Wq/Haax
Ioq5OrBLGCEf23BWjvDsXQxNQJ15qNTfxt1WsaE+24M1/QIPlsQHFhpELlgSV41L2fQjh7pTkP1s
T9JYiqWYeHR8LxKaG5cSai1sxR89W18NnPN/zu5yRkBF51hXnl/H6HfNwoTDiBv51vu/hqz0wGWI
NMierrkqiKfUbHiffbuxcTvEDhbZRSo6KWEQgrCKu4nR9wBS/byLaljk2zBwrxf718OLR/a9JI6v
0xPiYQChjvEfyHo4VcWsxPpwitigxN9MCTyvLUkHLm4C5g0NQHE4WtQuo6W0EffWjY+JgwfGtW/t
77Fp8PdQpLE/6eEj7Y48dZaQjo2ATufD+MiI7WunzBj57yYDPe5Zn00x3nVjS2oyuBOvMLNfJQ7X
pRyvUDotZQC7Lylpyp2sHfVXiEiC3mnWPSdtJnwlp6+z8d+RSYPcX3yHgNrno2qsTVWgCU3fESJx
cXe0VxmmNnNvfpPH8unc80notKOtZVZ1Hv5sWRb9aYVX4n+dFaxmorRc4CZTAzkytv8z5yHSbX1Q
Y+f06Da+qZFg4lWmz9gh6ymvMKBs5pkllre6PqIqXV5VXyxIjwAVJoZGpam2RGFvhM+TemyvWmfZ
fyjNM6OPjkEsMFAIesChk+g/+4ZsvWBOXT01FyRXProWYYIVbySgNUCU8q7GWiR9bVpdFsMkWjsx
ax6CIoS+Pl8N1Tm3XNa9T6025Z1lJdd4N1f4G5fCdrrrZaN+Mw0LMRo87hbCRzd/LIzPVqNwsPWs
3QkcOXYgNsLq6VqlCoTFzMCXu5HTc/I5J1fb1E6zJjuET2crCqg2QplhbA0SK8CNoYkDduCNQrLm
tgIQqnpz8lrcNl3VBFo0VUB9EBrq40Oy5inDa2FQVI1RBF/qwSg7Wnf4wVQgC3GOGENZB85iOKzn
kdu/llgymvmS+Txo1uOfLd+22hfn1B3boVhmQYMc3dKKQjF3dVYQBwb4Hv5Sz1mPhBCjxkVOV8iM
rREwxD0Ci3/zdk1bqK9egLHdJgoNekvd4JzhqqYmdVAefYkeotb2+pr6d7SCKmiO54Jinl2ROkUV
4hJF/YdI3GDKfZTuyZQn3YFP1dgn/pBu764ygYDTmuYqU39JngE3MKNGF4okZupxQhnM+8GCnugM
0y5b/MeJREyDcCUndysDmwVAsUJF4npjABYgCe4NwfYe2JeRXiN/wZ6N6oZsKx4KCLgZ2tmSHUWO
VfSsx4J8wJJZoF7ozcRyQXp31srdFDcSW4rbXrxjpuPskOl5Gq0b658yWn0CpxSsk592TsvZPR3U
UbhLRTbdFUO99TIMYhUh6QZd4He7vGgRcfEFttq7iwxr1VR3lK2R6Jomoijjeo6nIVxYBCpEcMKw
QfUTl25ThU1uYVESHrOEBZzTXZFjNMQM6kp9P4UKGwYmkhNfef8GhWkz3bxJm9LLoT8Tl+DUOefv
3i32AMVaRQ0vBqNso/s3nYV1IOrszUpU/ekvD6lakIqSczJMogVTIFiYRHiO+P6vZZ61bSqaIVDW
bjY9ouA9123C6Lk5OKvgRTnZvO0AUB78XMHwZ6c+ESgtA1nWu/o8qhMZKgRsU9CcoDpO0txeEd/H
W7UMisHoO2ycfkna9b10kplZyf7nhpBTjLdYjAouldutwpK94aiMSyv9KhR8BIrBo18jCmIe4uVg
LVlR3QAAYRPS/+DjnFMypoixoX+mlqpUY6pUccf4DQ7toHliV2kZt9j1UaGZ9KBOAqVvvs3Y+Gu5
GgPmN0YgJTZQmEdP7CB5O1g8K7wx7sqKQBvjp6wovo57hb7lN4XcBjLpEINing80r0WhitE7QUV0
c7TAf8C+zav+P/hztz7CjZ1+/R9TB1WmYqyNAH72IbgAvkx++QHToVyuLpKUvHbmsMcck91Z2N+j
xcFRFE+y7wDWjQnWXOU+ieztetCBmRhKVc4MekdUKjumqQW11yzxXSlyhuBeytHOgXuNGPSkKttg
6yt9fR6d/jTpJiUl7h9oTfwHKwCcYI9rynbdUjwMqDNmcnnOu2QTnmeV9MOO7wi+l8RkmvgI9X5N
T1OlxwnXTAMNIKvuHEa7cr1P4z8Kkg1ErGhmCnCY2QfJLUmD4UV6uVFCOjWfURzOQykiTxuqFdaQ
wcANYvmtHHr7Lt8w0FLwMPeDBVbibN/dbSkp5U73mRdXnRqKJJfFhDNWUhmWfcCwr1v8+qp3EM0J
XuYh2/Nx2VhfBWEDhPA7ZulRzVGbKvRIGodvS5yscz7taw5YrftOfEQ97UOnAGzSuHNLu462tG0M
7yuePSAnXvFG/PBG73NgZkN0AV3cLvMNuF0U9aKs4zAnpWLLpnQECQkqwt+ZrHP6ZzS/NwKHLRTd
67U9bd/4NtJ0lJfayTXulxinXdDool+NYi/PqNp9pPSNAolj/gT4CfNaRKy2pmBP5TVXqOgkfKx+
vSW4dZ+TFrRB6xZxQrJMF8+mMcW12Do/tXES6FzUIVGQYTHahnoUjT8pMnU90AqK4hbdYnWIKxLj
/SEjrvF97JDO7KfjHQDQjS45xlQ8IGp0fCPliVbo7t9+mvCX23jeU+3B8Fl+tUAruhpWh8ApLCzd
lRv0K9Gq1dgLnVk5RUq0Bk2lc2ZB4SZa031d4uE8Kh/z3LcAvS1TrjnwkPYZgOU8Pi9qy2KT9xm1
jNjoQsP377SZVGKpZFySfpiNOFsmPUMyZUW3tvpDI23ElYvjhWzPKZqMmM7Gh1IUhHMRPL7gyKBW
yD1k0DOrdYa7sguuecM8TGtHzJcCNdeDPmjt7CBq5CEuXIK4iJTpVHKU1LXclFGXjaNYQg8mVJb4
Ej0GyjrpPEpKogb2EfegWZoLBuQGuoLI/782Fe2mVC2Iz+NwOB6rMKj5xR5a3Gej6WTeUbkkHkvk
nNdKN41zF7lY2oYA9fVhzny53smWVcvlY4ufUE6UM89O0Dv1RCpExQoZ5Icp64bb86FDSOAN08ST
lgTnZ7M1WPbvniQoQv0U9RTM8HqXB5IoT7/if/Ao2DtXVHMDRXaYxtVq8nwhlFsTzF7m9h+a4zef
3bWEAk8xe3Aem3NfLiomjYCps+HEAKfsCJWcZ5V4bnJA+FMUgin6Jc33KCRYvKHfIF7tgsSVkNai
97SmmDHBxbwmDccJvS0It46Nb0in21MoWa7ejKF0SmRPuFJC23btK1CEH+sI7YwvnJ0Tuv0ixT/K
41v2ZWvROlaeTj97u4Yv/eVPbnKu3eX8RHpmDmv2lNxVsIgohsSe43HN9pwrBSuNg1fwVLxKDrJQ
48IbkkADz/9qpe9riD1l66jFQwxhs+iotTRkYeN+xJomKaNQz8GbpnC/RPTuQP3HKOqkbk39Z50y
6xJHkXyIDHLA0QxgBpRbsxvFvarcC8pLluWuHfIfwOmQQesfDZb3xxG3OVLcfNev6WVVWG//IK7D
vuqovgJQJebXsOr/YCrwhVsc22lig4R89jhyq1wdo3OwjAgbNBmlOIyQBcY2JuuX3OsUGOhDlodv
4L71+ASgFqkWd3N/ksPxSO7F+lF1RIkkngX8W1YWPQDVGV4Bn4r5Bw5JjdeOZFof3Z9ABkwa1GcQ
fwLN+ENtVcVBtUaMn4qh6vWYdYt4M6hfPrKnsnXbpxuiSpBV4/NBipcyjf9Q8GvKe5UcwKVZANkp
ju2Cj6Bjml3Wt6T+EYxNooZTm+RD605nS6Gs4qRZa5KNDlXU41NrVA7VjgB88N06lHXHRMTuIs8s
0bVg8F9EmTjTwXJgG0bfm1ikb8luHbNCh3hWOHeKCJyygwbq2es5JRk7SM1vuFAdxMTyxIuSI0BP
k+6U62TLRssDlI/RIZN4bLx6BDQ/NOjQ9Z5RKkTbgs0FW2gm74PLoWDAsKL3Y42fHLwXjue1AN87
qx8PxlLt0EJC8lzbsjy89bdaCD5vN9hmNJJ5dZkIRNDnuD46F/R5WotKvO82AUq8gy6Cqw86scj5
aeNgs6fpnPPiSdAGJkrZzyDZ0DfIwfbqIBIRgGs5I/7vOx1eLjjMBiMPfjge6jo1hsG+mKqEaBKf
UfG3s0FIkiFDOwtyRIlk68ndgseZ2/FlW8oN3lJTRHO3W+Jbkrxa1WFFFCuEhbYPa8aCX3ywwAEB
7REXI6lMSzmr6KjZe9gDsd2xLB0dQWdwhOE6gm+Bxvs8MmnSG5yMXmfLdaGPpbeqm8DIymQINmvi
oKqWyik2hIvmzkP7lrkCLC+WHr/clHQlLcb3C5RoHxj+avcLESKEDpY8wvSb39SncnyMn4nu46HK
vlZQydmpYKPVvCUDZOQLz0sce4NN8CeQ0D616y0q4Yv85sUutyZRaJCYKPEey8FCjl0jiyoiuCac
evc0i2oQf1Mzyw3xG0YnGACLpe0fJYSErQQsqn5nZvTRgePn58oMvrsOvDYuVTAq+uuBMopAoTcb
73j3W/HJXPANrHxZlEW6F13OJfyE39uwsK5ezl4QLpWTh0xO3ELHLRv2K2TDdX+xugpPN7uIxL+/
5+tB5wsCV2PESlQiKdkFXlsui7GrlVv+Q0XwHjlrdze4CDV4qWEiYvAOzP3yLUx0qKNjHXHdKQtB
KpvivYwdgT/piVi70lMXfEjbZKJsu0JMALDyJZc7A/aOHfajrpB4HgZvJq38qeFXpBNIhJdraT4L
nxdheeak3YN2ubVFvSlwK6KR5bqVE7cuBswW4KvdXFJr8nwQaA7v5HeV1t4EARgiAeTw0oSWRF/2
BO+VIwGHr1lqcB2x0WX3+b7+Wkr8d9l+KW8lgNUbrldXSctpsebhm1NVLdF33aEfzHuYDOeRbMp5
rCgE7XU9hBOgVyPb6C5tG6tOp6GoPVGMVvKmvg80V16Jp1D/EvAl/7CcgwAYulLPpF+XidZeHtcc
luGSu8Zea7aoug6F9zaiyDj6xXWH70bI6XrWGad4Hmbflc/nkWetHHt75zpNZM3ynf2LZRGWaNHo
3wnBVl0t94WoiHNfCxMxHDOgEJ9zTvU3IVhAfXwvJT4erlQhQGybw1MAKS96CWfR9aumsH9ZWM0h
bIkpVtNfvIvOJ9i2K8Mynw0grC1dCdUiM97M6TVApw4SlL3slao9lIqmjeE+H0Ss5tJHodTZyTKC
WAsHXnEI77C0EFyyqe7oKkylcsXm+TYIOvFC3iMASNOa/+qmqzUMB0EPOjwNYq45puqucV8ClUti
eMJx3xGonyuPZBLLSKrfOBG0gfn/Q34lemGUyn5YBWkdOOXxK62quzCnyO+5Ex1Rl4r+lJTlXS3G
CicFtGzdDUwLLKkawkaT44TNbnwOn9G5pkqD9vtX9twxGZR+D+B03wyz75nuzEYL0BpnRAFTq3nQ
LR+ahCSukj7CNOEOgyQsGsk2AEDkyxgaKuScEYSzGh789YQEDIeM40Aqfv47dLVYXfYXWXZaaJt/
5HvodZbOrEWUNX8em9eziFSPLrBfJBxTKQA1t4g1k61nROswhaHmCkPEtb0AAUbehvMlz8ch9Dox
g+zbXjyIyWjIhe5ujYv12oBChZYgp3fHzXfqT7yTpKqMXTbXXGsCE9Y+PG1qLIcmMQCH9GdhAgyv
kK9P4BJvkpFKtOi7GlgDMqB4V3civP/kVTZvmVGFiQydKAGiJ3Hpo5B7Suoav2xH3Hjg5pRXygN0
t0DTyYqDyCk4Rr65AWEZ6DBzFJ9n+xlqGh3CGWV+dbZ1PbFPMfcP7oPjMMzoS6D29MYoBbQFk+a0
k3rqnRag/SzzHKxyfCKb+uZWGZCHl3Ey3NuMtMtKZRqDRH0TWhbx7AD4cMwoaEz+SEXck5IGH701
3RzzZAqaVJQnsJbawN9ZlU2E4OzUvnp72DSsgQFfbWJyD3F1SLCoGPla9XF7vXfBp061UMbewx4Q
aSjdW6gKaLiTJvx8eQoff0UAoG1R1ccQrwg+G2pGkRCgYW51+wbXKM8eSXwneEoeVgdR05Nx7+nq
kLH8tHSdup90epbYEez37Cf/cxjluJihJygxi36OV83OURCWHoi4+Ic4tHseE+aTXlAxRMqUxU0t
ULbl6y95/XL0nRkB01BFNLjp3C/eA7Wg4zdat5pfaLLxTxdixfxC066epvqHVSIwYEJzeSAx74Jt
wBBn/xjNWG5uxZFDUJYIdiZqPStXO0BvDUit68jIAZ4DRV2hQXYv9BKUT80nrKeWFWn4zi0uAcrp
gUrsFsjzyqrgxfzXOD8GSMmHkL4f2WLG918/yLW7+1RZRHeJ1/3Pi/yCkcatc2HMqXMNu98PkzrE
XP53CzJ8SALVo4euD0c21luS+kYbQzkMVSo4eDpqzyCPzXQOnYARJ5qXCBzWrtsQJB/rMUw51NRi
Q3mIjHjk/+BIQ3JuVXnqB6ZRIHchFg962IwCCYn0lJWSRl874Y600J3xOUrXt0uZeaeLtvchpKnx
OzUwgsQ/YEOlQQ8i4v8ESn7dVmIPpE/BkEnDkFMCUimqgpxSE7UNFLRLCLiXFUiEQ91FZTwRbC5h
sg1WwIAxPNza5pVzFhjyLzZheZYp15wM0KB0LpCR6qvUvPa68T+iG9TSUe9STwNbfX/GzuQeyWAD
PKh9dE7nvKQLFSFIJdPbPWi3xKDMeTXmXUTV0TCTHPqTyKYFMiSuBttKOtlNxPn0xbMD6ZddsvkY
Jjvgb3Sne89PNEHfFsIGIk7tJJaqWK21Pc4Av9BuloDiB1TPKx0rz30I5j2Q1VWS4o9+WWXYY34Q
+Npj5H8Lu506NULOlsrbDpRhQjOPXY7M9DiNsF5QJzS2TggDDz0tTQjUMTtuhyHErd1PPVZbwTkD
6+WipcfCbNstqUwhUnfEJ9xTo5la7yyu4vv2z6ZhI59tKB93nYZBmtbJLzRIzbfYhtYyHL/2QKxv
XkbxtxBQjWXlN0N2VQSaSg0Pef9Qq4hH7hy+eMjTgTXimq/Azmkq6Cj97TILNcoaFt/FeuOzX/Js
4fY/lKyRShsWn1D6IkjLuCaLEnv/lwupnDkpi0NDDcFYvxVo694sTnxzzp+1KFx60m1c3/eQehDS
iS1XSoK+li/tSGRVstojkvAqh4RMiuqdJDmid7tHZoV06xHe5K5PLAaibRjefoFE4y/n+ddD7eJ7
yDVxpy0ucLl33ZbK1RZc2kfSXPwSBNY/B9tNX+kSf5QLzXCH+5n2Zi+bhQC/To1s2Cqy0xeb1wZR
Gmb/Ksrb8lZ4aG230wpM6zdX46sn6ck7PaTGjaKxLPlyKXE3kpyTXgSswD1uPfaWRBy5SyOXWKh4
5D5f4tiaR2StdgD0kqPqlE3a1fuGEPG1tpYpgXwANDWjrIZYXzW3KmIrqBu+aI/0dYtTqQVdhmwC
carlmXziDswGvkSmV6PlqIvixYRuBlvtEBHOHxXuqnJAvXrQi1z/VfEn0Par32/1gJu9wpE/gyK6
E86k/9CSq5YR9oOJDAStRmWlB5RWb3wbRBU9dG3PF9tH2w5VqtAOqXfV2ZvrX/fcBAofyz8abfRZ
T4ejyaiRpuq8hkgz/8fZvxLWKu/TWmO+3v0ZU3y5sc/YH5Y0hHfx7O1Ti2PCfpGvkGtfgM6Zy6lt
VUshNKrhILGsZoPn6Wk7oUilO4J2OM5cO0jmD8iVUlJHEQGW8fWnZIZHuECNQyxjWAK+Z5RFJ7fd
eLGekeUIL+T++KM5Xiwu+Bov1c1ecIIhpD068dN+kGToEQrDF/35ZisqVpUZHPeb3WAhJ0gdgQPq
sGcRs96Z0J4YgGikDhTmZD36pti6vHZQKB9ERsZik/88dpKj9Bpupon3X6yPxecHsC4WUCXdvLra
IzAdP+mEAr71hOd3+pvHrrlZAAc0C/xUjZYV66jhoB/I7XRedRqrzyoj0qynIYFUXbH8lRIWKMfx
ybnAYJiYKEZ3E2zUutkfk/l9xg5FuDU2i+YpKNyOvtJ0dx0E+NUOh1NTJyznR0GU3SY8zu0bSufV
1xyHUs/lks/d2ZYv063ex5OKy1p3cIGRlhTS77PemIpO34MfeJJ+esGxTgIIFf4V5JjrByAxD11p
t6aypkALUq5sk1OEprxCd4lKuHKObFuV3IQwXjnCNsJvqEpNfaFSmEihgXVvNJomhP3ajVG9BkJz
uoNy/1v496D6b27d3SkjTwpRgfWfDL369BIxzzoZMVOFnhAm6X2BnJ42Kzn1ykDdCH3hbsAyn2WA
gAXM594bwXA1XAokKrLhCp7+Y/3ftg6srmyC7v7dppAmuEvKWV7rSdOk4Gs8It8aFD5J3UEnnS+4
UUutYbo/pf1BKYfyTwtHoHSD0x7alShRCWZWq9Wumyz+fo4LcEnK+9GUV5hHtuTVMAJbHyKYfUCq
Zn4jcyNt+/kpCNlGtxVXuWzMDOrwRGjjMsmYM07R7BWyNE7XGrW+nMzexgwnGNgOzIS/Yswg7Aql
nPulo3xWBRFN62dg6oCK7T5p1ZURtRrjl8a6NF4i4GS4WXxpiSNuqFDrw649XIbsaijnQZZTducc
8303kMDiv2maLUMxQaERVxjNw9bhb8jH0DmkqrxH+Zq8EeZNDmzphWFV0OT8HoIgfZjuqG88yBQr
toEqTK/wMPXkA1gYyH/Rcsmf/aHFw5c/PZjlMSQHhHIdi4UzXvJqPobNugHJVBp/dxC1d5J/KreS
XanWMEg8H1GKHE5qm2l4N3VsoEsmtICHBFyRlQkDAFxN4BYhR+TOjngm1P/tTz/7zEtVZIeGcLuC
6AKx5VjxIfKnUWQYrFQtJkwDLX6DTFVLCjMmi1RlQ0S0rj+b+EaWBr7E5krgEBvdm4WBU/kma2JK
FQ4a/sRxqFEc/k/+BEUNVRkZaFP54aX7Kepiie45QXMEUPG0FpRimzZQeVFKgvzVNC4gf7GBPtkr
jaw+9yBt+PzBwiWnOPx/Y+gjjie6wrk0KUWU9rx3z1A5Br71YIJ3bb9tskyoY6vwMXuIpgXDpkjY
RPZn6xMDIQ4joWM3tuK6hJN5PokGBfZCQb+zvOruQp+V+G6LkJY7ksqc3dUJuLUb2zZsjTGLgJIp
D7zCCBRSp1FL/LIrC5f39wnXr5M333v/fW+MnPj7IoVmejyDuBCiWxnTThLDdHHnrW+6vZ0svD3T
DF34E7tNb4UOpO7inGARmYrvsxmvI1hysYZhP2yS9Uey1Y+0rOVKEKkHHsTIdFv9BqzJLfwCdZMm
fRQGlEIwdlaEiN5eUinNdG1L+bA+sxfNcYOtwEs2FyE3mYzjvDav+bjIWT2AOAYCfayIscL5tIZL
fwFWLQ4sHAC8KS9S5jBkFlOzT5uVNWY2y8spfpKrwI/3AiE4PCTvMxLeoXRuV70/oblBngIbaF1i
ZdmeuecWF54oRUaa22pb+ftKm7vQNmYr1vA5Fk98zg0rr01qawSdGMmFk1We2m3z5DKa20+oycsj
mWbSE8TPYuQuRyxy0ZaffiueFKfDHxVcersblGLTyR8saUUbhsovYkRnWcHzIoTTL19MxmtF4HVL
mXi90+x1SjCVRolgu4/o5apUb1nkCYk4OXpVjaZlv9fjUyYKkWlyYxrVaYc5Re+bpIFWY7bz31FS
Q5Q6DEigWEhCdj+z6k6/5eJgfNcAMqa9IP7zN/7U7RlMGOcfTABWDUUshh8JYoPOFXPpMw6Mw/mb
7vfISIM9XV1ZWyU00VIu5hPv9tt1R26V5PSNX1nMK9oqy7drRJbaupzFPT3z1vQwIUnPmdMheYMe
d3wj4Smptyw4iEPWxYn98/JISwv7Ybk5fnJ8hXezRI6iuqJCe3kNj1yOREWbqpIFUu2JrEH53R7c
xVpMm4kiEDBSgTQGWuZYbxtOB3yCn9XIZND1vbVqKJvZJrk0Hbl1flw+8+/7nH9DvVfKXLWGoP+j
DEJj7nFj0O0h9Ct+6mYDTJSEpDGUVfehEEFRl68UIrBRmcdoawTCrW81IXkkEQFwvJe7RBSYLaKV
loCpFo8miHL6PeN6tEfw0ZuH2qUFfOEN1Qcozcqn0wrSEqj66TIhBXWFdSW52XCmuxPkCub0DnkS
8jy6Sptfy7WIOFe+iK0DSkzHtmztRO5r0U858hBHolVGOAbYvVWNBBO+XjcbMRBPGJm6T35yArma
j0fxVGZsdYzsoOGRCHFEklkim7hd5XnbVZyoNe9kHoBragYQHo7CiAEj6ba+hCC3vZjqMPe77Nfy
QGsDW++U6p14wXVM4WL0NMEdStsHrpe7AE+OPGZzrfTA6ZG6b0wyh7miQYJtmZPHtDErJHfsSD+W
iz9ijxjhlZpU8T3jPwog48x9gawh8H6RMKbYuE0GTwUuh3EO9Rwn8Wng487XhyeyEcjE+eVu6liN
mjDz4RNAQSBmo33FTx6avd6+p4hmC2xysGyw2Ox62DofgvMmNw/2EoOeuW41qQ131Skx6xuKBR07
DoZWaff1tQRv/CZQLwPmxTG4pCvES+liLih2cR1/I+fFsYXiDcfqD+ZFtrTAHrEsJ2BmdRD3TBNm
1ygPbjREEtNAkd517uoXjSlN0JK3vbYbV/y1E+jeqQGaV+G5U6DO28OPR87hlzKdipz+nMxr7lZw
rO4Zu/RfmFhPA01RhQQf/afjWjPRW4sWIcvb7Upz7K+jyeEr71GSgmDzcHN68lVUuPgM+KC5PUiX
N6djxZX1fSwi/vW+9W9kYd0Afmcjov4GcgEvhOeGEEBFRSZo3jvPaUckWUy9lY/g3XpbsDF4UB65
CACmZ7NoDz/dkvU/KSb47CaPGhvY22+fck7vBEVYZWKYZuZSzEc8+JqaG7vZwBgiZ7do56fijM6/
dKTcV9xGOPadcq791KTGn70lYm6inNAdig6NRkrTxtR7ccU6RBh93ouI8sfcc83vgR9bQ/X2gDyO
+aAO1o3SFlm0QHj8a7EdEwLYIJRGzMRwW9oQDYaRIW6Fb89PGWs8t1/lu5TZOPLoMOUfyKDwUMYW
N4XxsHkIdiXL95ceD9kojZQcYA3mc+Z0tHDnMLE3TkUXWyPXuIVzytzUOulrcenmk8QXxrEl8VZW
polO2EcNXtcymkcoeQjzYHXivtwawHZrvI2tTgHS2s4aQwqD1hGD9TVp/AmhXwCfS74zbhxI+lzp
0iMuGxcl4spsPD+voFCXAxPOBhgfnTzmYbBtNX1NispXY7sOozjFA1TnsiFRd0Wrd3eJRZjMoQKQ
82JaauYQrqJrxg/PA8cEk+CogCBwTiy7pEhlGDvO0FlsuyUs8rldLpto9ucUNeXH314z6rSuEh9f
29PsNAWr2HfvykomWXGtBCamGmAoBpmdHaJMZk8mUD/hXSJtDmmkMUcVS6XTh6t2RJeixR7YnUCM
/QYX7USq4w4dDbzZp2lFRnoL7Y6zWRPvtnSqR+ndSBjpwHiRcXmHYx3M669u78EDVNMa1QuMYLbw
lIbNPUF4pbUDRAxlwGda/w6YPwVLAswew17r7RDeSyjiXN/NLSfknHHyk/ujM4tO55ueOmaOK2nt
cOf+17YOPAnzJDUs62cKK0zefbohXQ49t/4cQYDDqSX4oAwY5uBDL2P/w6Vx0nZJRLDFL7HUw0YV
+DM0sCb1GNMc4+g92F882oLebdt66VzTBEvBiycdowdMWUG/RSgTHEonI1p157r9rmeYidiWG9jd
d57JCAakkxGmWjS6NTATEvzYcXMaZScD2/98QnT7OxL2MXsYfyBE+e0e+3zaoDMAlt0Kt4COrk5p
XEjScnyC+NsMnB68rGjJMbJ1zZucTrpEvHMH4qBv4z2Cm5acU7lneQz53ZoSY2eiP2rROogkSKmc
7Y83AcpvTr/v5K534C2dUC/RC+N3fUW8X54NssPuJff4qlfop5yANFve6VLN+FVHRxpv2tFfns1Q
Jv2BSfhZotz/wqi4AuANjtOf4N3cYddsI1cZ+HQkLZ3jjSJQhMAY3WwZ/TVYqCcMYrc8gj0qSsHM
yCkISS7569wZJlxhPbRYv/ppWtVWR7BST/Jb+yS36YXt3u5a5RL7sVIeWjVACl13teOV1LHYh0St
T+tBmtuPmYpZHr5FiOCvylZJt7qaIrumgqXwmCtOAbnGuqXJK2/j5M5YyjbgkVfKhYInHDQZ7Ae2
gsAVrXk2xBtYeRfsBuqHpmrwpaoA42HcUfWxit5Y21s8b6DjCU+jzNhUmIESoR3bx+jMM+E79P54
pEipzk95CpOOV4hYqzxqnF0PjJoMSLePYky4Wdb+QGwht1F2UjA5cXn7UhIDhYhrLkwAEJ3q6+xm
q7RN93AHWhEuh1jXxiZAHKL2xJn6qwxyZOP7Xnryhm+wb9RQVCPxFZoUqPySbc33sQstRJ9dgCaG
FF9EUvk5igBmbKtX5/tz2rYZjEvO/25f/xXL++N/QET5lET0mlxwkq4kWxK4z/Eo7OlyxfJ6le78
/T7Qybr5+tlOOfuMfI2jgui78cD+y/4JSM8Lfgj09j9M693dJkjwujuDdGerCvLykKiSlm7qTuun
pgDGRUp0edZ6I4L/dpKSwcQS34vQEY8V4rh5S1mMKW5IoPL157PNcL8ZVCl6aHBIwDXdJAE7Rb0v
HP5jaVAnpKyFJKJl7Pt7iOCknOmmSpsvk4WnSI3EWln3Za/S4xNqrqZLtkCaTMxRr/mhoO2BLKOv
qQdacr1Itpkc+8gTm/zud7ueUfiBbuc+CBFPCNV/BjAOc0aY0v07j9GiD6qq26PpBixAyhkGAKFr
xd8soFB0BymfRX04AcD5wKb/R6gVZO25NzwY5xXkWg1KXteiL7BK74Ihn6bvuqcRqhp9lD+H8+KO
uWJEMPmroR6NbJhQu9DXAdB2gWCP0mKeHpGdIkbgZTv2hALLPwUA9ty/P75Ogx+qcx50J1pMVsvN
SM+TTJGGBN7qL+H4G+Y+Reb4LDSpOoj94pmZuVfaSFBC0Sne8Ed0YfDh6LKvgGsijsM1C5wnIkQ/
wLwSsF0NP6S8GfcfK94rYxHJyq8I9N21WKL7Fs/5mAC5NAfgmmhMkGd217n79mQcoYwJQcV42QL9
wNxzW5KKcTruYGoiRaVPdo2j1A4e6s+IXdylhR9BlzV72UrlCQbTeD6gxF/kxAjK5uQm9lqr5rzt
b6bKcOHtp6Gy4Ug0J4xFcChuSyF7koo1UNYmqbmz8bb4KuE8EmSOBcEFNiBwtIFkGhLHrIgDHoHt
VHqNaVltPIyP1rYER577P5YM7Ia2GSP+lkTGi9q0LT1np6hRbp8ECf/xqdG94JzopzJvUzIoYARZ
SYBn2xN7FKszVVRAeVHEs98MayR2G7VZARJObHaiYc1Zfb8UsWlXCP39wAgLKMlAa7xUcRAxtOHx
qgbOsqvhWEYRD2YsPfokTVNVOPNjMzDSKEfCD8/Nx56qLuZRv5i434vLwGPyU8QCyDPh1cVRlVFq
NChPHvtKmbgJTt+GkOJ2P5Lu+V3AjUicOVyauXhZur+/qx3O8/jn298BXNg7JgU9rcu8u+7+ig4v
kT+r4pTPYC4+DgXKeBh18jY9/IDCfakuQPJP2PTKGVBvnjVP0U8nYaG14Bgo7zZ7+HLaLoV2rq93
bkFxU1lFDgARd2a8hMzBY/4STBJa6MvfEcjyc8E5CojuHJhlHza+1OjhQ1Unxaa0fzavW23L/HSm
FvDKBiL9DskZ/EZuAGjZuXoOMCskxiNpxG6BDSmAIFfTHtnhbAt7C+gdS7Yqe96b2KrmdRzrcr1I
jSrLE2eM3N9TiiYDlHXfcNyunej5CH5ifReyvLG9qCk6wbslZ2n0rp6mA5JDToQvwli+AHC/GQth
/RR8f4tG2zBqHdd/fZPROaCRxgpa4P+WpUAYHLWsPkbtJjS8mzTZiruD0d0i8P6Vt8b78VONMryM
PpuzXrFMc1oME7cZWOo3QOe1woUcEo6q86JXWqpvzqCHFSRh2vaZwhsIW9LnQhO3KB8qItQrgdwi
eRJgKJ9fOjLlPBS/jl3ad5tElLCMkFAzJJERDTUuxnIIHdrwlNl6s+rvf6TRYDu235xTrfzGiZrf
fsLh+xJsvX4Jo6fySCbhsCrgnpGTvue4EHTl8Q/YkXpHXxJkJ8B/sIuxnbdQKC3SURffWGFx66Oi
1pIwAkqQCdxEP8K3Q5bp5l4I7WHWinH3rO2VtvdCyGcoZKkyMEg87+1GfE8B+fNQJMzmpJHyIsUA
j6c6Ti8VpIaYvYa4F8nadXsnF0eVhi7cA7MgtEu0XY7sCgUXztsD5Ae9kZYzyfFF8fy4FwK0XuD6
v50HwzVxWK2/zQrFgbjzfVWdiw/T1oUOkpuRXhmc426Bh6onUVsZViGARjuEe7duijZP/s3+iku4
WSpcQZMyfjYvXfTdtXK79bEmy6Xsp0MKCqUX27fM/TgfLOzE9SgyXlfL2mgBO01GwofICiX0flMX
dCqqf7I+12tkjZXCLZ7Czm+lo53hQYIj3g4BYQP6GDwEX6xek2N9C1grPmuKXRyh8xsg36Hbx2xd
fuO1bBIZ96wfFNyS7ZgbxwH8ZTefnzQnmwHlbdWfHq9ygtUeLKICYPV6Oc2lQKVoMgiTZkhJ2eiM
1PuXQk8Gw29OKHhUz074ejtszv6C+xdcrfNsETHDQbcZlF3683x8M2SnG/vrDhxUIN4aLc+SnpYa
ez9B3XSiqSFAg1dWfgEt8Hq/suOcOkQnBOaJ4G8M2ufr8/ztBF6jknOmMMAsQ98aln+Bv4sedZ4l
B4ibxQepexpEVY4GcpAi+7HCTJJGyYjVk/SHkAT/zk44Od5//TRudwF/LNFW3T7cOcfVXDwsEX+G
WxpmV8Fbt+YoSlwpOPJ6nktBsOCKfKSh8sWaMmDlak7JXQx0qGcyIq9DLSSLfWa5G0uek6OhHqeh
7GYbDeIHDg5rm+4tVLe/dVhRkemH7ByU6JZQmdVi3T2Qw5GNrM4lJ+SzRbjqqz6AOn6Y41D02I4l
ItAsIq6gLL+/qN1rT4FbXXfU1Kvukg8K1pQXTKRSTXbGkyHruStZHc6NM9tljOjSlVXfw2K94Mkw
Psi0DvXroRypIi0CrqbB5hpro4sFMMnE4RakbdLSnJpEnVMelThpWjkkra652CjP9NaSQg8fKJU4
dp3RsonBWY2ueY2j604lDLRedr9XRiVcRDt3WomEB4vnnnU9aZCJU1EkXGwATm0otB3D14dGC4zo
Zc38KRJimzUPBH5JR3MrhopW8rd4PKFscr7b0MNj5Tego/TXCUlP+2FfTs3Qmq3RlWqJhYMdFdLr
Jd7115wOz5kPZYi9MlS2z4nnvCFc7UArHnqxvwPKjX3OPgsvywYYJX1aP/ugedcl/9gvYliFnj0x
Dp3v74i/wL7cj5TTzQG/lcRZIBVGw5EMTP066/a0Jp7rhw6L/rphECHGoeYlZ5+VicH4BS1KryZj
IsYrotOqjbVn3HL+7YvQMz7lcacbjIGo+n50vkJp56OAZYmmy715XV7PpTN1twTIcI9bSf7qom3J
UT19S+53ctuvdRCkC5ii706xucL2D22im20I30tLB7FA1gq1Pw2luIqyb3L7t3Jv/gssOu7YvDcQ
EQ+ksehd2k4wkeSclWlRVmcUI5X4t6b36phXI0jus8C8NNOFMLx0hTb4RARvMpfCdf4Nu70aY+21
zQdFkoknrpRrDNCDMcHcZiWbQBvlrZj5Zq/yVxbB5HyiwX5Qp/xI0vJQPlSJ6YbJedFCN+1D9nqk
0nwj/I7y2E5CfKw7INSAxpsu21JbJFOJqT59tvtuutTEuiC2O5krDZCHBX7Q1U+U3cWvJiiCuuxo
B82c/NqgAuqo8aFvYwelSWgyiQtxJeKcwYtOh1MVzUxAs4ER3Dg1POMMYgY3deuiq8o5fKyLxo2I
fiHs3ENhe9WjZE2pDFv7bDqQ9EaR8LH/CTH+/ODsbP6jwluhjjMLNLSFMYtmxvpCXOuVRgPNV9y3
0inQ+qi2hkIBfSwYsbtoYW3zZKdC7j82zZwht3bjCZNud45qeb1DT7nTxB8U1PIsOjOlFIEcGHQ9
kQrULpsK4V24gEIgA7L4HvCa8R77SMK1fQAWc0oyyY7Rncf7ZJI9K3ua7JG42Ubm93QhPXiGno5n
ArsZ+AWo8qdNeUh4o0sD2RbmVofEeddc4uSq3L+WqPxj63vJNTZlmAJ4kRcIua5B55PpKBbRpBC8
aclbLmQ7RJFyWtUUdYkg+Whdz3irOYZXyyuBapmLbezLKEC7QNbovVbaE9xCQ4iTpk+vJWHMkr7N
2puDlt4gX7Cp7TVzmViC1tbVUe5hqvbNO8v5tcv4bW5LnUfNGUn99v4PH1/uu3urXEWgIYkDlXp9
6dQo5pBG95B27Ay8u4dAZr0z05WjhAtm4DO7F55daralpb6xK0QLPtSZhAUldKbiEg4fFnGfLLuk
R6Jq6FRz1otomMB2ZfNLnO3h5E9xyeMwqtpnBmBsG7YInS80FuaamrwVL7gZQ1CwA5h0GdjH4a3w
XlgPyoY9qB063pZKoJpfONCqY8bQFoH1o6pQkOu2q+52NujqGwd7eQ+ZCBDMZEMJU2Ny9dojsczp
G53LFCUT2RKz1jB6R/yofPcCcvGGWtiztiBwtR2902yrytvkbuj8G6lUx7dwylOv9qUqltKrnPNP
pSjx/GjAkgSegzLq46JLdCm5x93fX8LTqWjH1BjcOoTV2J8kNNRb7gpXgKQRWIz7bByQ5pOniOpP
BTzheenK7XnLHSYY09bUW8FF9rZpl32T0E3PyQQbdk/wRoWH7By6vgMoQKI4nQ+Xy7yDaUcO62nN
i6GRMMx9XjLhbW7NzoiJcVLkfdoRO9lUr+hjKpI6kwRE8PkZ6oGrVg0e0z19qaORDitOGlthV+g6
J6cL6hR/s7Gp3Lg5fc4RVBCiKRbLTIJZFnbeDxv/bL1Qd7pCw1SbEZ8Y4HBBYb0wcYOkOAvf0VLh
S5+KvGb0q9E2ME08EenLON3w9U3tccZkeSzkL9sHRqDT7TchQAe3z50o1z1665OtuLXv4wBCks3L
gmKzhiR+33HoR5811Ashmvqtpp9+TaBp77tGtP+8NxEmWxQBMUWQhJhud/cVnntT6mXMe1og+kZr
PLx45st/mmC0l5nKHjHGn9MZ8StwfEKq4nOa+HJlyXKq13qfVyNhwEd7spcZ41igA7tHqFUbtSmy
5rrEfoS+XKBr4AZP/mpTfGd2Hc3YuMx2d6GhHtcg4pe1gvpq+JRnBVgZzgT1eyzA0GWrxEBFXFCY
sylM/I8KQV2h3XNrZg2Dy220Glfh346tyJbCAXeOL0dIqL/x16jxpOlZs6Pu6idJcF/nNFZOWsrU
llVIi/y9l4URsyBBArN4ye3opWclMLU7qxE2eX9KLsJqMTLMta94r2DLZY4OE8dTGXYxi/WpLx6O
XbHMu+IUuUdJh4Y63zztrqpgUNOUOTb/TA3L3jUGYtOj1VVhSwT/Qak/g9gbKVe8bMxEw9Sx8xKH
DuTo6CPU5i0r/xw+nJPJEmwX2cKqpBod4FkGZhewx0oH/GuWmY/rF5QDm/7UeM3jaP3ihTT0tOXX
VpoJ9Lf1Nezryo5Fu+/lbeMEYJuA/sBThqZP9LcJkJLTgccK6xIqsY01Rd+cjYcsb8TFIA4aW+ZC
fZvywylw4IHGPRlXsoQXuWVjhUQzSkdx/UxPg1MMRAm1lxQpomZ0wN5PR1Om+n8JNauHixYI3+78
fmV7g4TVpLhdC2q6cdzQmuyQPW8ZUoXSwwI8qPkB9v6o6cZNdEa8CoeWDYEq7qmtfyBCPP53lWEY
knIGrfFWlwJlCLWaC5UsEh9/anJbk1Tbvh0GECPi6p7J2nwCbtT96Rs6cX4GojsffuGoww68W0z8
Bpqd+/EBf5dfvn4X1H+IdyWC04xFEQAgGFLPXjsGMqm1GwNYlWWRzv5gBsGODfNcqA2o8c10jXAX
9rx5vDJYam6IsIi6SotBg9xKzYtjDrHjRrRLJ4mapvMtJDdaUj/+th3+QIr6jqlLvmRAwjx72bdJ
i13cuvWcDbiznIRVGWSc8QGjZTWR4kGToRHc78TTbbZgUgyKnKskT8DksB8L3Mlno4SZRe3GkmgG
C0zNSvtmIPy1InHMkwR9T83hO5jAt8os9uzeIlDGMnN7Vtm8njdi9eo+Z3lbMRwUfuTqneC0Kg22
hC/jwuyCnVOB9hkceKz/CO+zXPB78uDhs5PXlAAQcIt+hEnXYjO5Vj1opoKUBeZhGA3bpWA6s+7x
PQOqoS0PAsAH37HHXYNx/HkqigAzIBegEDisV3k1k3CM/oakxr0ds5LuptrafFMxJ7K/hmYdTCDh
FNgYXu+rm4/U/zPEQk8vxwZPyfu5Fyle0mJFZJTJQzbfXmAa+SCgAq4zQv/itIAe3AA+mM8ilVTb
O4K/mOuZLhmkLi5HH9lrr0dltgJWsfqhSsGWEJcuu9zL6tmxHHF9OKPObMfJ3zOwV8TJBCLvIQmS
p3ywExYPWVA4VfkB7pUXI77IU+kjvRdMjRg3mQiIIROWUzTya/hdOTvxbr6KzGC5voglh/StltAr
tOaBLDBfU8kXXqb1lNeizOQF/1seq7lmsw5IuMMtnq7mfOIx4kgV2zGi3Oy59lnVeFNm6wBjiH8T
AWKNQahkShT0f/F+jdrvSlC+mJxOfjxHcuNQDjYfuGPFw7Dqv9untwRPIiZuoJLn09XnV5gLniaL
6rYVWdxDuYQCri7W20/Hpzk5rJg3TLHG9xu7oTqwuAWVmHL96FN8Kni+crHKz1q7iATxqY7c2TDo
+m07ybmVR07hvNBwySlmB5mTTAQJ820ZQP2+zKwsUX/58b6etjjoW6yqSdgfUh7SybDUhyHWULdw
LQBjxEpRNgZjRXHB7cyLCbZTb9u3YH8hU1MsCGROAGtM0pGXLqw2YSzuZ7hDbZGfsB8DIEktF+RC
PyGSVToiyZl3rVzDbBveAkm6qlIYsKmUfX/0ap3t5dko/R2MPacLhzeVNCyqgb6aUS+6lqnVb/5m
bpCeuwJ/f/uh7i111US5AAu/sIuENE/0VB+bBkkZzuUrpzboChNZ/eSC0yC08TGURjNOSOP5pNmp
ZzkqWZDKa44lk0OtshNXM4JrAE2+I6HiwcKWLlfTex1Bujfw7KD0epkqPzYYuD45gbOCqsoC2mit
s3MNb8X6UsrDJy+Qq4D4u+eu7EU5Ngtt0JRzsZxl7loMX1JAxCnesNoebxXsZsAmTE6t6LgOcLLo
lT3s8jMVY2c1W4Z0iYV39ihDyqSWE+bmLxA1tQqDp9ysZVMAMnWyNSIuWqS4WNg8suDcLDwH1dt1
VBxycvMq1H/NfG9I5fdaxXeQcta/C1m6SHkmh87jKN2FNYYOAHjZLJF+VFsvQYpZee6RZZ9CjnMo
3k1GK9pyG/XBkXX7ksM1QOEgs5S/QJRvq+4jnw56tW9iUI/RRqbbIDM5P4x2lQeCo5wfDIX6I87m
DG9IbU0nnuyxa9GDJSUb4gxXwWCiZMIMLOT5ZNvXjEZBFudMYrCaU6Ldj7SfPp+2w0LP1/CFEErS
O6YIw+siBwo6WdYuLBDx8cAwsBOh8+w3eW4TZzbukYzvCKE0SGjRslAxeM3hEU0ZSvty9efn2mw6
YvPUrtOc9hI8pPFaXqGeOwl0Dl2bvHeyIsfHnK1U+G0McPSgB0wTnwyqMpPvNjB+NMje2yVC+x+b
4yEmaqLoS2eUeKcuK62ymVNn2jRYHr8emz7vWNug6RqoaL/+vxTNaWSrz2/Ai9KD417Lm7k2yoen
lgvv/hk57tRNUhxWoDVWXfApkHtv/tcE7z1/WmjqrZdxPrpRR6B8iRwrPI+7pY69L1xxArH35s4l
tHNZxwEVVdDzfUnhkQLc2biveOc2dR1/9pTut8ctysv1ElBCBiJ7RjfdEwR/sJYiB+05i9f80h2v
22c/Hen0wZ6jTNjQqb76a2foDic2BbXSODsB0FX5Ab/26qQBcs37DagTm3VMxIql/77W/xCtLHjz
PEONwSNuTVy/4jjPWMg7oUdqwCRF4SFJzda8aye7oMIB4MUIVA6vup1O1Q6E2a1VS0Mzj+vYhUGZ
TFBHWv8tlJ9eCa79oFky7pxfrcb9pUg5vU0Hb1Ln1eF3NhQQmjvwz7VvucxTnOb0mSNKkUZophVr
PfUKysrYP2DonnOoaQnQRHhIWLU8Z9eVLnnrgjvzusXZV6bCGqLCwtBJu0qYZ5id8tX7DpzPd2By
uVRxKy/5GF/8KcmMTYI9Fkm4HhZ9ArjuCZUxuB6+lpvG81M7s/NGB/tvagm0Z6+Tneop21WQh4fE
efd4ENFic9+yQwNZslKR3cj5jkAoP/MJFFHNA/Vn/m6CkEMZ27MXWm0AQbOipv/X0u9FwI3H/PQi
X4X+NzVjliVGPI+6oaYXSQNR/pqV7NsoP+SGe9POeInHr6O8ZH0KxWHSfwjeTxIVEs7VM1G+jHbq
QCbAZHawy0/3BtxT/TlzboUHyK7sFrxv2lj/ZnaGQ6z1srjeSylU1aC7h+xuhSEHAKmQYBhe2UY7
/TTzGt59h7Cl5jniDAE7GvCU6YsMw3Kj78bwX9bVl7IFLR7uCozPVaeIZnGglpxZLLd/2fmFXb8a
l9TkBpnF9EAxJWkwYlBtXDPH3Tpk6VGJYPA5NSqns7hYmWMNtG8KsCoUiMicswPg6howkck1qZWQ
kMtZVtJh9grAqbVPCYciDMzi5vKEmlxprdIDgcqptmgvzggqQotq3HE7NVfNwfXSGQsvw2H2/LfU
mcL5OMMsWRfmTms5cXBhVNSljPXHnxGbkXhCf64aLN2jas9tY2E3mf2SlfPHq2AQe9r5i/rpRGVA
ba37UBJsUBKXNmoUmcziU/EdmyrH3d+hXhj+yKe56+TQ6z241op0tXZgePqI/JqvN6Xfy/4PUNMP
K6/kcfmI2zH274gdUp+w5IczhoJcCvf9s3GIkhCDPHA8DHQFEfMY42YsbSfKwmkF3Jcs9HSucXr9
qSn5Ur5Vp5rWUUduke02faxEV7v1JrZy6qZQkAKAVKX/HoI9110cJaYp5fxUfiltmSC6hplh8xdT
esvVOEGvse0jwR0/2KpZkltC4gUr1Mo4Noa5l6bH+QAodcCXZelUK1YLj0WgAW21S5W2pJcyrBqj
NNGg/4AUcrldxklnCsp2zkRZwmyvVEsY77OevGrxpH1u6U4VOHaKbpm/U1KfOcHUmSgz//FC9IyQ
aR7LFsZQdfginjSgzMDFjKybfHC2BYpVy+PJNZbNAVPm4hvMNT+pRBSSTTIGtuSVVX6PYIpJUdIs
6yUi4RkNqdUGs8hAsyAZTRxTipOew4yJ37F0B8JyszrUxzpw60iwMmTMxhvZ92sUgUbQSOyJB3oP
1mxLTmIm7iwfBj4eALxzKYkFon6YzDXHjH28qfleM1mnSKkFndSagpz/QOcRu809cQETzKM65McL
rmqjTImVRPkiUjFFfDClctU7DUJKetzCqF0adOq4+9H+i3pdSNKQ49vgKU+ff6QYYrINGQEQXb7e
yXOl+rXyTlAq2n/NmGFraxv221jguVBbUHL8qTD/SCLRdZ8kkonKlzDnOyAh5OQbOL7115krvdBo
PbfxwwJwz8YH2kMf2Nlnkuczf2K6c32/fXILN6VP8hOAv0udGFn5D0BLCQSAMBz2OozvdoOKV2tE
qSBQCV6CM3Wbe6B6Cqb0n3Uf3upsk8JDjra4hBEnhqA+5kWk7iS1ltHZk3SjSfskzfSfcMi5rR4s
3QF8F/06Rk4zddSjJRxsn7FE3iQME3RDUz5sLkO+DiMlHTh0K4Zo6KA7iDQ2Ie9T3hy4j0hcrUfq
UgwCim4foJuNTpJCJLsO9QZW+uUCWczKrih0P2prFPPm+pAgzYfsR2zssHBDphkQwMT9Y1Phb7TA
46pThoVCh9huy+1NCstyHoOp1SVyfyTgsblsqaqrTPzPnuCNE9SQCJq+53PY80f/ai8ONxvPMPI9
w9S/qzzOnD0OE1bPpc/DXwEhNLncUNxTIbf6Qsmt8A9uamr6Pe4tWSSxOkEiz4kmVeHuO142kjUC
wVHtxNhs3t8eNYGqrjwXqs2wWEPXo3QbF1/0whafIcz5LcN1+82KL3mW45VYiR4DhI6WCHGcn5df
WTPin4++P1TvuGFGwlSlUG+WrSTH5TWpY5A4IFLn/3gS1GRFDFHLz7rrsj84EXkQ9J4NUIwcjrJv
+NKUcECtUYJz4XWmRqQjpeET1BPl+UzpxF4parn5dlG4FFoomz0gk8nVWmAWia6J+4pWbSjsmAqF
0PCmu7ZjVaBUrUTRrB09Mdn227PygRVJt31vhucIbxhUShgz7K6eJnuH6FDmwPDNt2EKiPdUCNWf
uoqOaMS0ySB8iVkig7eJ+eCvUIVUgCmfZWX7+zgdx7ejFFAg7CIBGXZLyysWHfiiTxrcHhWMV/ik
FDCabr1nmJZVxKI3THnXGHhY3JEWwLsfaLD2OmQnM+jHF/RCZIzjFSY26aQUidtbt3cWAy2z/DaK
eS2DcpWFTrwPx+vlazItDNRiMDZmpt8V1odDwUj9HNyfJ5HluDMO0l2rs8X0T4xtzZkDsrOjbi1v
npp+JyfpOVOSnC+BsRfMPLlhJ5qVPsZ1KWjJ6Kl2nf5NXmTUa4QI0qtHp/KlBeEJojWSoHTHEegw
dkkPs783I03uNyPzkqtCSGNmGLyU8O9KBdVFpLaJN6J20nv00JHXpFyvGk5vjQxQ8lPemXzBnRQU
Q4XVJ7nNVQM0GkW9f2pqjoVyviJNh/CSiW4JfbIlRoda1MqE72LOFcLn92XPBIliDIvVxo5Xxc/O
hl1TLin6NUKaKh/Ew2uUIKSdflFKqYXQ+KicwtMnLfNKI1+XuQWQBFU53Qw6MgPTQFKOta6p+SwQ
fT4xmkX1by0dQR+ksutHDPcPQzOsT3GtXyyUWW1PlnLKyLypxNKu1ZHvB4p1X26X2CmXOZeElN6h
sKMcU9bFGAPROiouVJ/WfLkUVftfn+xCRFYw5FlMpZYFZcprZ/vJ5F1R6sIFEk8WU9kMnBg5m35B
59FDWknQp2RQXl8SG0fLMKSQfijHo4WRsdnHBhQd568/VMmtSBJ1teiPqHt5p6flem88qhhEC8sF
z8uEyfMinEQjtOPh7BYyjmQea+amdKwww53Gi+qfRT/VCZqi/+Ou7wj0MwIvdDH+CvYbmzdpQvVZ
YfhB2Urk26OR+jcClJpXMpJVPfsLJI9iyrL5B7eYNHpBmuP1XCt87CqQdm9YAd0BneqvwLWNvKw4
C/564FvDcdoUX2+zJLvQJDd+fZLc9i+EOS6L/tty0mXLDA5FTIrf5baLsYiqZ93AC3uU6EWLw1vK
saH/mGHIOalkcALcboVOzR26Bz2RMG8ZxlsUKNdCzzRjnJQOGqSTZpBROrZgIUK4/LgXOkIr9oLA
oyVsbGDVQQcqAUu8PUSDxzbL3G93l57TFknDv4U09CSmYqwY026z988CdYUmVKh7oAmNbGZJSwLd
/8+HwXY3ZqEEOfRptlw1khVosd8kjesRd0fWKwqP1Glr1o2aT57V5CVc7WA0CSP+ztjeEFlYw4+g
gcLJ9C6BHzvVenYXTO2ES8+7HssEfK9RR+PmGzWNgyWYQTX1h4lxUItL1pqgyfDI6xoiv8mC9SjZ
hos2pDLpQ7pf7YiWi2a0TftOw4XfI+Deeaqb8balvNSNpOrPdAmygFhjhTIGyEmiYE5QHztiqyUZ
crv1r/oa4xap/uecHYGgGG5hL2diBQopExlIXUmUMIbABubhuiAmnEUH+EjryCYGyuWyJC0rQjmE
4qfu/KEZqTGvZ1EfSwzS73Fwvz3GFJ2ztkKJSFH6USrrnIsKejFkmS29SVgjOyjze5UtfKC1Bmmw
SXZlWh/sqPcSm05axaF7yJjWIZOWi5+XtTgNIou5Mbz2BC2u+iFNlwq5uPaJG/9C0KGOXjsvBIPj
HisXpE2vBb8WoyBGewWvrJWS6wjg7A0GY0lwuxiDRSh/yAAJIAT+foXi5GbwCBHznMy3uWDtPMLn
dhejvKVfh7yjGVZYSVnNoGR7OcmISrc0Z7rXaQnxkiDjv2nziJ/f4qMGRC9CHYu17fgogQsEfGg2
AA2eSY5a4sanCnHtyLyUYVHFH2OiwkIef5wwNVFLge+3OmVqd1kxKXBameRv2o4lcQ5kc1eopT4+
g97QBGgzMysYO7SCaohTUfCptdC+cE4Au+BsQ/wk7gCC7bPL2uvK3zUfmfO/kl5xuUwfM84TiSor
BGuwe5pGxhG8KMsRsgjJ4J5tS2ba1G7C2LH/CF4pWgdLePhu6mG+6rEFsb4F/aLDYsbeNd8eRTfL
vFtNig6R8BWyYoTMc8iHxWN2qQmZYdOaAQNNd/sTgX3iKb6TJpj5ozXaelBMlTIuy9v1nsUwXLVj
hf38yBcu9CyFeq0s9VR3I+LmHijrFjOjDhtaadFFVa064d7BEy1qMdJEgpt4rqiQCuqoKovmWzBl
8fRnTt4xIWaJdVkT7QTecmWwKn7XMMq38NjTTyP2b6CBwZqRDrZ3Z5BXNhYBE50HnebIkopGqBtq
fIbECUumWwYYVpTPbQufONN2bpKboGXplbWav4IZ8uGkln9yrfGgXNuZCXnQZi6WgKdwWWLHKSDh
s9uUdcL5gihZkpK54egoMEtJjQUx8/qcRE16gISbjFVOjr670MQU14UBxvOuB1K6dWxhzdZ5WpoF
vArt7kNl3gE9361fYI5zQSqh9RsMl63nIGoMxYlmOCt5RTMz0hzNEOHonFw2mNYo5Qf2oolknvUR
na1+u5TBR3fjw4hQcbmiVa72KPRXIcUDNCG/amgyv4pArNoEQWTYvg99RNlDRI/KJfTQu9rWjhrE
oLL2MAvgAAEsf8WSYtaoV2Ntj9glR/DBDnNAnRGS1TjbobSdaLoYYCe9hL6x9xXlfdjA+SC3cqgs
JYp94Flci6w0Cvx6MWOey3tbNx+tiwF4HAECgT2C5OMm0aVtgW14cVJhbRth3ktzHp1y/zmmmun4
sHqPvz0OUeB77T90XJte2o1Z9zwPs+56V+S28ITNnhPovuHoEEEbf7XhrLJH+yMzn23KQPklhseH
Deu51yiwWiE/pVU9jDCYvw4vX0esRL+qLtCEJDK4OKa3wmNv7wMEICwPAcUNz7/yXI7MiKfeIfWu
2bIXPx3kUYejOeITZ9ANfNIwYqmUoGg3O7Wp74oJmN0NJq9X6gsgD6r/2W9Zd+BnuLE3Pui2p+Iz
ZH3YYFF6/7lGNaugHzyBo52JUobThzj77eX8jnGbSpOXQ3kPGODjIj++g/BJkbnNGi/72E6NcGYx
z9AkeprhGf70qRPWczNENSgoEpuxIjm8pPrzQ1UXGyXfHhlxIkGjMDiD+mBlhvOvBMkV7NKv6ek6
c5TxAO+JPTqjNhPTvmUr48gF5oCyFvctg5txRj6WAu1iMFxltu9lFEEfNrFKmvKRnUjwDe679LL4
UgqOHuqcpe0ZRvUpgSDIfWJvIIwJnYFBOBasl1cucB4iwpA7pcPsE34GETI1XI/BwjikI7wNfYAn
+S1br/SgXt7zqRNIJb0SOHDcP6FfYglJoObANetWvSHvce2Ctq8AohUY24r+c7aEMygmHj/TTkTm
C1iSGfnTHO8qc+kkS0oDzL3yGyqQ/Cog+/yb6dQnc4/JXK9WaGRUIBgGHrJDxm/BxxsV9Yc5fa23
yiAGFQ6uDLZ/ehkfBgL+iio0ZptXAESNpSzLxyJyDIP1gtvnwK4+Li5klSGeuFOXYqJDw7fKuHDv
/wQcqO4qn3JPeyLEJxqEM0Co5dVHh51Y4ai8vUbVjfdKuNLZYY6EwukDClOghWRKkyt+uxQ6Su3u
WcFmNUD2uggIIOATzQ6qtMa4uX6UubWtqFuHQP74PLz7HGnbKKaPcnTPGe9DEczU7xgTw10tJ61A
VzMjWqScIFnklqIKhJZldQh/dmMiC1uV6qZSF5EjUSX4bMZjNJ1IwFSSHsJK9LYjgKkVT8dndlJU
Gu3cg5pk0ZFuqP2aR0uMDuSNybNrHwIBFMfEcFX4IXL6QOmcIyLaEvunQGpngLXM3zBVownDyrM1
s+6KbSoOlFRxXVgU/C8BK9oScFeU4fXzA/X7Sn4sOTTnCzB9dKu8vjG4aXYZ4PpybpTn3JugxB91
+Lp3Vr19VSVysWlq0KF+uZvRO1gOT86CxzXDMrUoDlC+fprIZG1AhXRqO9Y3aXepoXIo6plYT4x/
/6omopGb8mHeS87/wKR5T1vzE4OiONtNdCLS9x5bFElfBY04vijHT40s59HhlGGvLNZ9uGAFQfQz
B8H/fQoe10BXRoZ7y43+biV2owtGee0SwgANefKgAxJUQjKUsygpBNX+GL5XtwWjUiK6AwIA95n5
VXg0UfRl2E4Umyt8064LWRUZCisSPrSW7pbvRmBYekSQYsNk6XfY8aWzP8aeoMGuae6/F5lzLe6h
LgzCFTXRhA/08SK0fUihPo/P9AgwgBDxwQNd8bo6cisUg5+qFC41jaqDJGo8837dkc5xXS3G2yUK
TRt/14doCg9de3hTMiYuhcO5NNlW21iEYXetIHmAG3Utl5NhQVkjs1YO2Pt+RPJbI+EU3oYkJIao
xEAhQzqRQsXHDovoOP4/DP4EVs/SbfmoBCUKePPk1JAM1OC8zsygs9mmbdWdkgVCmNJEoZ7qVXe5
TA+0PwASD0FgxLEnBWVRouQAefMiktPbfM3cjFfSTsx9mybGucyIvPqHpEZkUe9EfUEGcnMA498L
UT54g0Tc3fjYuww5cOx9SUISO3tNyi9R/F2BH68VipO41tmmUBEMYGN74nnYctRAghT1RxXc0Efi
iFoqK/6upXoajlz+ZsijAI6zYR9Z1dwW9qhIRoTR4Y7RF3umJ+c0VxgOgyvbrZiMx6z91PlE82ma
QVBB5ITr4l57lu1IaTriLIr17QRWfPWQ/jcnyiIzz96yMGE8+weBM9l8kvao/VU8F56wPuf7RZpi
hjOK7hslBYhvlWTI9v4HiP62EtUSvFLOFxwJqBi/dZcGKDt1hyZOyXvEDX6sx77HfQycRgq9axIB
4ops/GzhMPAbx+xbMFx93Ae7BPTtjj7OEyBz/ejuWc9XOkl2Ek4E8NmR4gZlXhf67AbRP3EEJ5Wj
ktifC2g+7BfPbfUD6cxEbMokn7wgUYOuwSdYlOgyMyPk6vSTkPQOjQ98ea5gu7EQEIm7QwcmDTMb
5ZwtTnZxXzvqe0PTo5LFqmNbETxLrKSFaHmqQVoa8cygwImwWYwD93cBQflSblWeilOpaewqJFwL
OAwCdKUSJIlNCSAn1vZhXwSK1wWMqr5yahno2GeyVROscHxa4OC5eWKh6t1DPjwM+akxC1sVT0dk
Jzn2+AOC83gPwtprek4EnukMnkTjAn6CqsJrOH3mQMSRk47qNMV/gFGZUW4W7CjNpS5HpE75xEFs
0OmP9RE9GhK6N8PiTlpapix2GC1Sd2z9Qnsjh5lTDos2TfPw2ccKU7wL+yNJS/XLQuezXDPv4+Kt
pJhikoe2wAUo6WlV3HplqicQbhpGbcIGbjqqmLUmYxyIJz8e3VEbp7ZtPVIP7by/0pHBrCXW9ng3
g1FihYQx3LPN9+0Tm77ifZ65I7eWNEzR9efj4NBbf6WSroR77maawfwrWvmOSZWgxfYOI5nefa8x
hMoxkHBXxrmBXfT7/o70ZwXYbD+zl93EHoj7O6KhRxPq//gehALohoJTUb589NOLFH6a1V7XkbfL
jp1uOgKR4/2+e8msdt8e1B+o+hIkpBej7xqGcXgco8AnrD4oOSu57XEzaO2Kofx0um4s2kqByGrP
uIemVcugDxnr4aEyARx/3ik9CroMieexlRcJs7a9OWkbF0Ipaszuk5XLLqXX0bQ6TvYHcqFQTJYj
9HwPp+8msqdv9pr+VUxlm7dOV38yU+Db9PyzZSsGfgTLo/dSkK4mVD6KxNdA+CLlrHdovxUodLRO
tL776rIBXo9IlbrY7TciOrKhE5po/ivImPZELJ/pQdmBDA9ZM95O9bvryJl6O0RwwSYi713qYIH/
FSa4T+Klq96EWcirSZBXyT1iEHqV21kDlnnzIi0FidUUjrplNDBV5iLCjLMtHOHABNJWg1BV6JD6
hUlIO6FQxS/rsujDA9IpM0L1SaXDfeJRwakwXuO9LaBBoM487Ct2Ibt9SeW+gYnTaZmQZYX7U+We
b9ndp/2jQTiGNTuadHTu1lKJ1H3Xe9pDbNxc+q3M2PYwlZ90QnC2Dv1p8q5ba0L71P5S72xW5cBK
sf5rcv8Yy0AkopSM6D+ucVFun2dWXmYVjs8yRaTLq36o0SAmM5yLLIrAVgPjDbPhVx1LMsMadtiU
yuMXKgjraaGPQhkeFVGXONHO4c+nh+xG95ifsQ54Vsqd6vnP4QgdFMYVK1yhp9AVaKWnlV58/y2s
Ss6+zuMTlKuyu6UjmbbTgLcN3xrOL85DbxO5DXgYOUSqsL6ty/5bPZhWJ2K6QhGV9hepR+gya1Ax
AtCx5SUgJhaa1e8bdEvAfD0HOsIzHUvpr05bQVcchyoZR3IC7/MIJNNtNIpMkhBvV0JCsp7pTuSy
aB5D6HIzJLRY9hWJCJjoohxOpoPf/E0TNdDyudDuZ8fnPEPDf+xSWc64mWv53vHwIaaMaZG7LHIH
VcCt51LQ7kzL/4GJ7Q1nvpQgc5JJ1aAIO1CXYYppVlvg/RY6GG2/apNzN92PDNcnIAcIMOfiFXFH
2XdEbAiv/0G3wRdZn2UWVwGPYdMEA4Ij4MLCkmBr37CPOiJU8pdEoylteZjbYkyyPLQYycf6So5M
Y32a+TzXEv+atN19Xl7sHUZs3sXzTOgPSHGyY1i6ln3eiX1JHIYqGVQXya0Vonpz6UbAXLQGTV7W
hpGK95GvwiBovk4SyhheHm6TDQJDRb67Vm15GwgINYzezptanAbWAlIL+fi28VLh5BtBXdQZ3Dur
00rk7guBv8VsfuJHLYitlQ2BAuQ5qkyo/woZh8wDHLo3bN1db3RteoY4MNiuRPPFTVs3wCABDojW
L+pw4p0+ABNcFicPgnooDyrC5Jq79dZUrTNktHPWWwgEI7yLJiWTxEyxaCDn5rnhcUhG8VmSs/5z
bA/eQRGsTBntkm2kumrwVHozJWG4iA6F5/8YQUp6bBqJGht+NPVLNfC3I25PhsbZj2ahny4AZIQj
+NVxYHQmoboaJ+Mlg5kni6O7MuKFD+H4YcLyJFuoYasSyLxQdmrtVvkZFwsBgrc8DHSG3hkJ9YTB
M65cEuxdeXWeVAFAID7zRiASFu5qAYjWgNfJ++i8ikgjM6hx2eC9MbvAlaK4M7QNBFL5qaF8DzGa
0B4if6eoWv3C6StR6l3Mi/QHQCKbU+I/xwVcUt/Wo9SzZNnF41SYRvJkifMO6rAmv6hIaZlKc4gz
f8Ohu77WiZnfo5fBOCCLWVvXlsQMWTM2QVpTFCoaYSzaewSXWsmqCWaVoyhNn00E7hl2dTiNaJOt
3RXb8BD5LNtwqHQiRrzDPD1TSEUQJ8ROyR0Y8qfaol7LmlQQLqCNR5wzxyNnClhnU/CksnI/cg4U
KDAVxo+VsSfkU0v2TtQAtGQqd8U24owH5mplwOMVv2ijoWF4rAsL8C1UYaEVNLwi0+v+tYMmGuXK
i0m9VDYlDeaT16n97Jn3QiFmAXXQTltzimqfUwcrXDlmrJ1EuyfQOS5Se36wtVX4S2f+uvNJi2JZ
vSodIIGJ6XySKKVWm7Er5V1Jf2gMdSIOaOWWPoIUcjZ2L1iBf8UsY0pMIv/w/09kLtZhLRRSZ95t
YKW709NlTa9p1G78mQ5nJvZwmSygOP3OTNC2iifEypNIrmUhKbGwfCzafuDuAihMx15EEUjO+ohv
GnuC+SrLE+sli0ghM5cMBJZpk2ie7megBrCd3Fk8RngRzG6v0p0if7W1u3/FCGNg/7msSJO9Y7X/
cP1J4B/Eph9Jf07MhH7yqDa76Y1dMlHSkqchujHZ52Eq9D/zsY7n4pUiv6XWocqvWvM6AXRbCBkS
OYqr5avhPOk0glnfUI8lopHcwbFMpClwxNT/t5zMwpcxSaTQYGlgau2AdzUkyLFeRgjfevTZMwLe
xAY/EtxGXnmFoyB9k9mD5SASXHN6swAjuc+anYasrk5gDPIEDldoJSI0ZKDGYEfE0j1rxaJd+AV+
GUwa6Di3VHpTg162GVUwO9QiP4sIbpGsZtYBBuatdOVhJC6k1RGyRN+nn6fMR1xvFRV6YfeIOef+
ZGpmMzmwplZ5QXRAxJWMvlObYSLFyxRCxKJl2jsqCHcd9Z1qhRN2gWKYU7TKi8IPfSfuP4ZcfeP0
Yz8tUOXeA8SfmBX8Tgi3H587q0s0pwh3ElYw1E2AgDLAaheuUfdDErW3F7xVJxL99xUTQKp0lIXJ
Gx29rqfR2ZAXfLNd/8mGgcluDANaTiJuWccX7ErtYTOBfqiSu70uADTecTo/G1JxhMGbeVG8QMob
xO1zY7zkf/3MM0la6q4/HMGLptUrvxaXB1HWRqxsl2sw2/tlvWtY4B42WfQFO7LZIUGxkYXMkWTS
//hMDZmQ/fPai9h0EV4q+4keBC7++cuOKBPNvBUdv4TWL9HDOE1nZ1j2oVbaQOvgGHW40if0osOX
fLl2HmQF6I5gpawcxBD2i+TQmkLi6lIMUScBGYkyMeVkE75c1Ct8mNqGViWBWl9FITXTkn34Wb2K
kh4YQodzmyyMYZjS85h7XZ2T4xDXX3wzOGi6OQ8i+3Om4CTMV3PLYWAedxUNJuiDmKQmKlW4yE+y
vItXVFUXpUeVqpPPO+fcLBh/fHEvYuikhzwmBIxw8jrpfaqClcD9GcvsSrms9t/vcwmxSGjrIe29
8dV0bnXJry3Eoqybfh3a5o5/vVmJGkl+PvAviUDDnCmtIKiRUPiHKgrcA1zTdanTZMVwD34Qz1uU
1iUlTdGDrsgqxnY9YKNMF9lNg8/a45BcVGVx9tFlUXOJ420TC0KtbUlOvrHi3B6VD9usOH2+2WeR
MSEswQmlYUybESTIgGo6VgMl3MXIjbH3wGL9yOBjFvJFnz5AeY2SCQTAedCG9TjGXf5z6Pz91D31
Fv+kJHNCLTpFQBhRcIpt11re+JbrWVMfSCZEPSIlvtIGT/qdZvm5d7QSFIIONcrR67jfHp5hr6WF
BOLCZhSK+zWFLnJl+/BY5S3Fx1K+4oL5bG+yuZC/hmohza6mpOnqnlT8EHoi9MRclwzsPMaWR6L+
cIBcITPH9NQyG4p40nqrHk0fvX4YOKJW0yCCeBW3rr/o5YclJWSq55QgLNTGC0JVznnhggx9cf/z
YljTm6W82Z6a0G3ItbEi0thY/ljze2rrH7pYewcS9Yp3R3+z7lLKQLPtFniNzBsvBQ+SaVe9o5Bk
pkOB5KmrAoo8QprpJYZ2ulu5YSiehvOAN7t19874EHkmRON65qswq1YuPYySuHyyqWPrU1YVz3kH
wCXb7THEbR+mYalZjybFKnnbF4BSMC44g77Oxdmzk2NrAHKezojl/5YjqureZ6ueDeEdmXlfxXwC
ZE5Kds7h4/HpgZeiqB+OyAXJYJnwTLXPrljdyIIkpR9Vj73WVhmALXgwUjE7siTnF4ANWPgwkINx
QZfwm1HphsKetMj+g0sL6s0jcpgjLD16nWn2Yv5aoEq9BS8zx79eE/ipFtTedtox2O9FYtGn0+Uc
PIp7y3dUpPPSmZR7uknCnzN5HlXC6xP764gyjh7JBwlbybL6SntdVsLIJc0uk4as1DuoltRI8cIk
35bbayuuXecnmxrwf3Cjt5kF399qF5/5wMeRgCw+nAs5+xWuTEfQdmnPqTBX8U6FCSh9SWNKkD1T
BRS7qpPx5jdEXhjg35IT2eBMGj1bHgWwHZ4sbrrgmQDhtY3Ac5DKrvYH32hLKETvCHaT3nyqQc2P
txuRxFXOjgP07k081OiKQjmEXuYAeKo2qLJPy+rMMpiYn14nbwFu+iqHDUxHE49UDK/CLpZQSYjg
22Vhhjh4q2xiIgN5wmA90r0fZUSJQ9qNc00NLI6XFRYuy9CPxYIaN2JMOzkYsD+0KCeLDDHu66s0
fJjq4cNiibwoUr07dHvMycDwxkkeFcypb6n/SznnBDDlBpOrmdVJOkR2Foz/GqRQ3ORuGf50/tjG
PpE40jLeChis4GzvIigR+GEXMerNKwm1xtyiiOHtpXUJLEIA6S6aJCdskjXrbO0T9N4brrkDsMWh
0BJtvr7+BATjmS18vctu5pH8Val3eMVOzzZ3O4+uW2LBlbNyN/BWYPruElnGHpTgYlKduobDuGaJ
8Kx4D2zOmxbZq7nbdBXr4zoTUwxDKiyZ1p3YBJyzHDCGJTZkCseZyb1lSz2Zj4sPjxDe/pTJXu/F
jIOuHpbhDS+vP+6T9v0kRfrYhQ2cf1/Pj6lEie3/zuyYeOrGOo2ld2sgvhFyaAelGsewi6vFwrMB
Zx/ouwreRB8mqn9JHlYGgcjxEizEUKzIMPW+pZ/SgXT9GQGszHAushfRdClYSVpYlITUXpEt85+K
T5enIoDCjLnIuHgwJTwPMPQD24gBqjiMcYVz9QLvmlI5JRWMNTi7RGXkJum9YtYCxNsEf6J7u5/z
wx1p7h6Emj18i98koj2b2b5CWjWnikap9l2eCkJKER3L8XG+1rV/e/bJDkuXjM7+IKnyaXeXQ3IK
cdtONnN+ywlRn8D970i5GSMo87ggmqzxSYagnxV1zWzA4bpB+kzfxhC1TP61hYFsVijx/GLO9LEA
0FN+V9xz7a/tge7MX0xMFQw4D4g3ttYeYpem4udE4rX/ajgxRuhryoLP6T4SHZy7cVwLNzbCSsCx
KTJtp9IvUVfmIPiGwsYgS+Bsl/RuRur6apFqICyjRsd1E0an2U84N/a0XEkLk24feu4evw0DB2pz
mWzs+h+NagpGrDfDlwuyi4Klz/YPOkeQZf2OoHuqSUKG83t6/psp1W2B+JlNV5qQsJQcKi9F9ISw
4LO3mrgZIs8lh1mYF//ZBUPPBQR0B9OmKA3R/LsS4hy1SHynnjTlvzZmCu0gP+jyLbkXVaLAVewm
d3mQ/5ECM/5PWl1Emmx2rUG+JfxhNmzGgvJ6W01jqNoODbwui8OvLyohYiWAvsgsJkUuVcWt5KlX
o+w3o/MkY+kwxTy8oBpvjpgEaUdRToNvJgllGuZZixePkjrb3I3R2lX0Sommn87VpEMyRqrUE4HY
W9LloXynoV0O3+mkbdh8o9LFDRyzZSLzDttPa3D6DGMNZGxTIN/iUC21z25H624xTNzeqm+BDW8X
5RBkU2ElR2HAml7dbVwFwC5o/NSX95lCCpWDD4bJttyPavy8IxaLMwV88VwWrCAK5hqjHAWFQHhm
yuYlGVjBwi3qxSRXBWoydPbQXE2sCLwInBP6A+UyYUTP5zZ7cq5VxcDwO2SN9d/wlhiX+IIyoq7h
ogY1s3yfRfevCqLs0rbEafa9jdlX9pNlVmVhyElDD4z4Mp9ABralaPLpVc8TPlwcvQMttfT2ZgKK
oLIR4uUydaWGrEnz4a8JR7IKktzDcjAjvaVGiUo8QNfUPRmBfWcnwpNwh0H34YhMwEH83lWJmkcB
862JFT85nJ9588741A+X3llUlVCC7mQ+eA45J3s1BSNXshazSH9eoMZgG1iJ4Jgol79PZUCPAyHi
MeD4un8XpCce7eamzlgmrYukS0oFMluDFCtbFGZUGvac2by34mGK77+TbDeA/R81YWMgxFoJwnIC
0m7mgpoMfGpk1aoc7sYSJTnhxgs9J3T3bkizpOSYSS19ICFkBjyROkqLOtCNLbsclcsGStwTRbw/
6Z/8Wj9kqWwRsd21NWZNcfCItko7xP9FkUPeE6NoHH1egeEGCDTGaHHj4plqPmrmKvaCmau/BKXO
NnfkobMfU9bLBV1b67pCktIWQIhzTJxVT4EFU6yn6hAJwzT5UwowC5YAD/ARmW0DpJ51hkIfcZ5j
dwFnTbQnYoaN+NglqLhnwt2ZKZ4JjWrUhm8Tu9iususFlKCXP/eCWKDAs88VQ5Z5zz7jnxnPcdt9
cFqE0BMkm1qVCMmql72pjL8hOImJzGmFv3u1Ts4VmlmOT1Q1AhBIXGV5nQvs+C23Uo62Cj+5ovSg
mdWzroAUv90opbpEcgf5QuZJeBSBYtOdsb1BOsXJ+ZBfMoNABmClwWxHEdGkrAYq3+wCcUellhBH
f4UQD6lPz+yKVfb8SDSWDMb3ZWKGbr4sMJlPmrAfdc0Cwod2jtXgbHIKV829+Krl8dC+j8/3D8aS
ELLmOXb3GcXUy7q43q89xjORjbmaabsoO3MI0cditgXXSZQXZ6zWgfsRc1te7btH9vBrYnIIKc+X
9tioaBm1I+A9oEbO1Mlr5KF4WkRbe6IZQUcARal2sQd9i3aiZLxcA/Bw3tknCYpAexVAS82i7xS0
RjSaiakGKRDhY5qOdg57RwHdXqxjt14Xh6vMpwCWV9BI751OPz4vnhZcVCByjPjPPAkrnlsvkgWs
rD6ulI9XSvlTvk2IwpUb6cHBpv47SuO2uDgES6hxWg1UBKdCZrhlS/Hj7cRyIjTtFPItVMgOSCRo
TV/g4tom8wsSYVL0hh75Q/a9pOtIRqeAMGXLJAgfEgYKB6o9d4JycoQx/Sp8jyOP2fE48B+5EAQ9
A/+8/TmSm/zzmEqY0eDhrOQgeWSlVu79rmgiWGOEs4ocH7xYGTwK0j/kqAWiFGpUqn0Vch0TMtlk
p9YIbU1WPE5c3uLlAW8v64zZVH7iYco7mQ6T7hLHLlEZOXPmktuty+9pwkrviwwpDn/3G/yTqIEL
Mh8os8mIANMxMpXOtBozGakWAH9mHTqJ+OPOHAhV6LhWfa9qt6Biqdpqa+osZjkwnX6soghO5jSi
rxegeKCJFo7ZmLt50tG333xDJxsyHK+RPEhaqHjjpFUsLhex1L0Rqx9dKU6BbqmKgAlpW5gqVcMJ
S4q1bIUVe9GI4whPEkvR/Ekt2WOuw5Jlvo+h+txWX7o3cQHwUvNWPde+dyaLN1wxjiGC0RXRKIU7
IDWVTSQRkt9UQuapcepOTf4o8aGrKBaFA30Am+yBn8w/j9j6mSz/aRaGD9yxPLBHkYM7p6lZj0EP
lMso5izCdTSwcTUefBonkW4eQWIkhYI2DN8Fxki6uFCQJslI7fNPDtSnRQHjEi2XJ/gpBzjjme7J
eqc8zR5hmMeH0LGjV1GqhY+IW0iJnt0c/v1XDZshg8z43HK80fwHc6azVVTs0tHh0Pm7miMdd74j
Tf5OOkWm6jSLBmlc83uKplnIjOeKKyRa65720hwA5kYEUDh+aO3iGu7owCqgPCkTThiKCngG5v8V
PH9ZtBg54VrZt/uL0XDG4II4fekd1EWZXLSk0rY/racQH226TqCsWIsRpu/rtr4OZVyUxgWPCa7i
XtscykNgit76U+MMQV3s+aopt5KlOom4qlsvT34iWpEhtIRWOJPYUDVVTSpKp0s4EBFr0xfywoIo
x3sztmxpFgl093YCKzE72jvWwoTlQ5sZktx44+ag50a091y0YE6NSzWDr/rnyyAPlt21PR/oKYye
tQRpcPcNBEFxAzY4pB4ZYQgGdWvKN59HsfBRymBEksaz+JxOjDsUmugkN+WAC30U6cyg6mpzEsX3
mNPLh5ntdiSl9Pp9SSrvoeubIFlZD5Sktl7KiSEdqyt/hRojlazQ6dP53CRk3RTD7++XRUTlGHuh
wjQv2Cz3YGNJ1RAtbQeUreuCNdRdcChNXBhjMt0ko0bBpwEDj6ANR2g8g90llJ6LRO0N3U7GSzXS
Wm7B5ll6I28xHkSpyUIn3bdGlbKZBUJW+MOv6j2WCIF5ejW51LfZV8sOz64wZSF5tHJMFbMnjJk5
Z9JLzDu5x09Kkt03SuIzC9ZETH5Dbl9i7hZ1R2PfYfy/2gMze0kZuZ5Mt4TKrQu2oEDqOC7B7rDz
rOWLVzpRY5LXbMKQ1m9AAxIyawmtgwA9uXddR3DXTLqiTpT6hopmKFUgwpHyYukyDjXeoKvGoinp
m6gO1CuUT6tqA7ItAETyXOnT//nkVcCkPJiQRSr8o7CdxITB9ae1HZo8g9XUQ8CSPqla1QOruO9w
tj1b73KzyxIDbio/e8FmWojbZmyP8muQ7jmVtZp5Udx9BG5+xKGfAw7Blslwt5UskoEypEiBERhC
4NGRpyAiTm7Uo/17cXTf2skc6pssSA+7MjUrzyezJm0WwNlftXYLgzx8MXR00QBd39kQZHaWGZnF
4MTtDDg52q5CcdyjxOSb9avy4rgXnvP72BUf4v0pLFdRgwe3nSTDUPFjWAdKPlAeqcBuItFuNh4N
q6+0HlhXe73Beswmb8nEGmR0QUeOkrsIoxIalkOOiecn6FTEAt9Oywv+/ZcMNgCOenm2+nFXWc8X
s2BzljINvee3D1fLJ+18qoIx6fAOFeATgr1uHf56OoD4koXgBG4Bfj980JkGMUvv+1Ij++CCf5hn
zX6fHL0E8t2TIc3F5L5braXJ8gWweSRr9UfIyfTc3Sy2k9jBB4oqP7zlZM9rRoMbW17VBVKpLkoa
SzW5U1+6xqxxR/yYLXXy94zvK2JZd90wkvD9WjCKxe01csL+7Yqv+Z4/aQDGzRfE6dJ7uV+Bf1Br
TKO8VawGPXEz9O9CXCIMMS/XaPkwtcvL3/gJHxb6RL2Sk2tl7R5w95Aw3UMLQ76onWNks4h7OTm7
XHotgF+9bDK2MP5GujL9VZ+dpzyguwxt1BLE6WYV4jN8YIY2V3fjyQ6uiLZVgtgQB1bzR33WpOcz
MbkgXiQx7edGF0edzmG5idWQSetGobdJ+kb0enxxeNtQWKCPvnXh+tUytL3hdnSFUVkQcAjn9RnB
mlFLv6DH3voF3gLnTxBdz5y7UZG1qUPv5yt/2QMdhn/+Eeqep8i7Yh0o4+3d89BYNWfCOKX4YQS6
CXRyBoz/M35jHy0B9i0mQvFe7VVZuD8+2uz/uXkZGSxDCjh8ZzGI/vUzoag7HVMUKLfL4O7nXjHx
zZ9rPbsS4wDSbDPxfYfjb6TycSvyqC+a8S3G+n664ECNe44QyeHnnCvpsB9FDHz2PJL/NH4ejLc1
uU8MhoUVGEIjY7pdlQVqVCHUSTVN6q+VTUo/elKccQmApvR53qkFTfRKAgZckuDGxZJDjwp1rXQ1
RrYZjformWjVHmOFdZ8guBFga9gGS0by57MrnMH8o62XK5aYkZhaFHFu7Jol3fo9j5anxKin0Tvk
rvnQ+zQ/otCX6iRAwceFgLs0IUzed2jCsaK5x54Z3YL+6wO31qg16tN5AJR5f9w4FwOMdtabhJZF
2lVHwk2c7mLnB/xj/JpPhK1Xzeq0Sjy/LJKQ39N2Rh3LlNxOaYge/F8ikW5sOhNMzGNrm89Eulb1
IKZf+dOYTQG+kyS5RUNQ5T3gWXJZNXayI21wZtldkNlOIlCApOtcXQ8PxrNXPd3o657d1gBsT0SD
jtkFh8DhrSK7Pl138Wxpsns5rTT4bYrRccePbXDSzM4dwbcnF3UgSzV4yfuyNS/tMz1WhP1Pzaao
2q96XDktuGkPUo7fqi7UG52ZbMzvNn2vFJ1CAYfsyn0gBVuPoQscY7u16kyao+IK2CNNzU6p3Fb/
ilSxxYbgYijdZm2wr58kNWgkoiZtZKVdTQkjyrrFfYinX6/B6OEB+y2EEMHxYY42ODxSfLS6j1ks
w3mlh3onoht/JOG/8YB/UrCV0QKMjKz+Kf60Ac9Hk084G+HqjN4i2KjG6CQUrL5Anxfr+SqAAZ9E
CZOIJXy5jLDTo1Etyj3LvFvOoQ3Uq1BdeiQhhY/di7uhfFN6FSOXICAzcXMhiuSS4d5KGRDqOD90
yIQVD0EfdgQrCs2RVbVcCJi0xOA5hUtNuIF5AfA2D9wKzis1b+sHBBx+ZkvhkBNrSo6K4f6iMCRh
HFx9kmXm5bYhEqHYJH6xCP7YIv0ZPKcIOs+EUMC5R4kIrKyv1xsYmzP2CblS+eXewiIEnSHWLuSp
SEnWgBOTGNxchYCjSSghBrEOzBf4bBHhMbzNeF9pHEa26ssmvkzTJq8q8015vbWxPpMs02Y88Byl
V/QoWj+lonaTwYexU+Q8000JlKyrLrkTvZclqa7D+cG65SFcDK6NmENvLL6EAkFGey3AIq/vX/09
mHAP5Ejf7THYm1oELgxpo0jPfb6CJcFjSTRkkGWvHCwS/bNtPo3DGCgErQvkNsqgUDhGdDeZ17Mz
CIq5mM0CNx2t+J95ZkS1EfgiLP0EQPZ0rV5S8fxRDmkQ08B/WlpBnbYNi1oIpdY8CD4iwKrKu3AU
qS+7YR/AZAo7jYHoHbjbNaZ6ZWSiHRr/Hb8HzPiFDmr4AK5SEcXRqIrP8l6yylqaV33cmuzCTguo
7cONqeYkbsrwvOAtk2qRY2PA8+6f28XbZtUzvKfpK5MqxdQfExtCILHHYWXZEiRYpVA/cjW3iQzB
iBHPEqQVP0ngkqsLAkpzrRggNDpIYxuAxxrNQP11Ew3kOEcYLihoMQDXRbLQ9U6cLumi2ut+KDtR
aoN87r6n/94Mwti3h5A5ReW8l2G3T6Ooc4KXMsFp2yxD3sFyz7OY5Hg+44+rXOdYRNgBbRZkxau7
FRIJqPzA7N++IOh5UnxTcQsOkmdvZD423CCVK0UBMaRXSR/XsQqBufVM39sK8HyNckM0AvCjZKmh
bpgGVU1cgzDExxWriHzC3hApAA366R5fJioRpCHbOeHx2XXMRZIaisv7dmy/xApIOix6IBNEB0Eq
JOU8JstV4n24nR0P6yfUCFn5vlWYvpZOUpkv9PZeYphBQ6gMGrDeOEUAS9LiZnx4gh846HZTrRxT
gZB6ypUtFzywij8wMQQQQC+B6WrsDWaETdp94CvcrDL5rXnKT5tpjTh5KRXGNjMs1h5i6nTBLHvF
NGSVu2mFD5jRc8/JM7kb9Ri3JPXNxcA40XdTGvtDh4rAfOE5AbAeHXpDz0VtZWbwtLNYtyzo8FtS
I4Sxc3C3S6pNVTVslpQ4rBVS/4oDn7MIlIh4Ch4zlAYOS7ijGfwAtxv1P3teQs6qrNnIhTdSNYQh
W8BXHkA02Z2ySD8zQGudMbCE+lZQ4fRL1PVkf+e6ampMvu0q5+F+hzqk73c1G7AaAlLg/J9bu5EC
wv4+V538HfSpA1fWyefhhyE3zitGxgyJA0CFAX1p6lmatW+ml85xBFZbhR0bW+xQbMcbHv/FZPRv
0ygnxZchI/R7pfbunyop1vsdn24l9kLkrJPxtrWkAXqxTHideU/UX3/vaIEe6CQcrFkLYXFnWYmt
ubH3qrbHE+LTyYhn4kDt/yhMrPjHue+oGXOqNO0coqRiV44dlNgwP4Plo0/rwHHQuoR9Tx+SZgrV
ftV0p3gAAd6+MQaj9RZbs0zkajG8FwIv4jLpl1byvK21H4smC/T/n1MSAMkTaqYqUrUXv9rB47bx
KY3GFi7pX6T6yA2cZD6OoeqLI3GnLuDYikQYFVzJ0jwK2WNzkCTZJmH0tOfivyM1FmJVNJHMdg4J
G1aMPTtGYUY7d2E0zTvh63DqyaVY9FMsa/jamJlexeZnnofCAnr3I9jnVbFHi3cQB0D5+yp6ZPyE
Cf2yNyR9yGRAw4LPk7dGebmrcNkjEkM6Zxc8FHxQE0ixo5ZBQOw29NXvCMXmCxh1xZXCkAMQHPXv
EOpaFDiIGL4vuQUC678nNRPH4EomdCW8r1EOusMvepwEnsDHDsCjdV0ggUvh3nChszqlLYFGvbG0
fB8t17V1d+BGLyWMmwZuHMgYUvK0kMyGtjQBuY7PaE58Kd/OOtr2AgYRtq/ZNCRz6kqqeiHtGYFn
t3h0qURYw2QG8EP/asxJw7E5gIUUwNp4wiIBQm42WxhPlyJXBhkpq5FDTiZD/1S3306KfTDxfokL
E3XAAU6xSchR0aJagBRvm4WQ0CHWb0qNHUu0exa7bW5kRMijIJZKEwanp8IiPXu66dBUbgzPdY27
XbeWPlClCgZLc3bwTBrrxUljpPXKUzLsYOjs+RYxi9iDFNKJHKqKkx5+6VMMWsN9GMCefeDL9ZEm
tdSDPpRKDM8JvQKuO2ySSVHDyFrwFhvRVXrhreNiJJRxs8GO2dWeGmiovHUGeY82pGCgytn/wrxI
Bo2p5CHXXxTEOHMn02a3bu1NQZjSiSIn+wIXwLDB9f6Gz85roYw1QF5adDKYivsnRqSGFBYb4usP
uz5EYcatM/oWk5zgofSy4OeobDkolexTohKaWrP0Az5xpwhw4APcgl5/8mdGovYh28aC5OhJ5igX
ibaCSfbEZ07sxiSc5Bw3A1dg/A2rdCvwZyakHPAH4eGY94taKTgQw2ruFWbsUqrn4HtgDcqwqVT3
WKyoyIro5IFLq6No8LeMPIB/Wh4RIKZKV9BRnyvB/vzSmGjF0RPKi4kMJO1WMR31tLNWw6/WwJUU
bsKXjywW1w73NiFbENjT50mab1esYQzuWD0KwfLSVb0PaKekytuQ4KEVzZOt64O4irHJ2DF4XG1d
CEnu/3K022qhpandzk8tUq4xA0YDYaQlS3Ozyl8Ktve4P8I6J34fOD/Gi+FQUf4EbbIoDHQhqr+b
86NgaaaGi/fhNDkjwOYqwjNSQ7KiJRmXj+CoBDwy8JQFvfavnPyCKv8+eUuBjpFpNDL//DSjlopO
9hG1/gDEiWZgUp8CO0VBg+UJYieav0g7YWTCM7BsEMaCfjXmLuAVS/jeRcwa7YE3Ze37yUdaONjJ
zhppbpk+ZRW1WVJHpgaLZohoXr0yrjqDoPYOKg7qPal26PXeU8lk+ICSWSlD2fhKMW89qQA7Haix
Lbl3Gu85RPenxbOonmR53G3U77kOk9+r9yGZH2g1OlqdjdLQergdZ9FZLrchbKpGE64VYn4RRlJf
470IFHEYuPiUxKClxvs5u3RKFh3hLNMfrd2H2PLBOQSpa1qc8W9PMaGastdMmU1Qwy6hNq9qVDjJ
7OX1IZKWcGDct4Ds6CxZvIK25rf3d6k9VrV96t7JIR/w53qPVUOM8uE4oc/l/yMPaWb2CnPS+3p5
NBedL4ltSq9B0CVMijdjrMa6w+WrV6HbM1YXQnC+b0ks0umRpT+IaqWVdDFccQ8eqwA3PpBwMoNh
YILhoX69atReRsJ2tt3efoJf3ilYGOZdZxi2u7f4pWhFHMdPdvClJ3jPmTvKU06N/549g6GzGFKy
b9lReswD02QnayUVH+/JP/ignuGrVL05a9VYuoNd3B5mPhGUOf5TPEkYH344No4SbiL4z6eTHXbk
ZmrQeXy4ydlm8at1lOHxeQ2jRW60m7KeCbgYSu0hw6X12wzOO4InAYQLtIGXrNrfILDO91jHRMUK
jYnKgxRkDWdp08yeLH/LA7mFrBR+XZIIYcXczPSoUZACYkOsZvt4w4ToQSXEZUF08GRvlg/pA/on
Imx6/Xh3LfD1kY7anFAIRWDfefesQRde9CpINmkqeT3mXdKc+MGQ0688pNQW+aTrVeLEH3HMj02x
4NXzIRjUiR4QjNhif+4XP8lhNPq1+4XcFCn6SVs+dGU8n10sd5dRXH4DIbvCDwd4nMQqGD2nZsoO
ZDprXSYGEN3EHaKINEOEaYjavCgquKvryFPUd5wAVBF8UWADIAVP5DpUKADhVfjE4SqfCyvf7HMy
oCICcwPJ2Bt+O2BcQ5B6AYdJL3UNm75rFAoL+3k82O6stOoayoGgc2HOKG6N39Uuj+3wY2eYIr/6
P/LDFj8+fN/AXicDbYgUUHKyw/WdtsHbZ0Uvd9y2u7MlnvI/3pC6nllxtD3qm8769A8Wm7JRsED7
HMNyNtexFlFgr+Rz3YmoCw9ZbV1Gbg1ZdMugly2iwrS/qkLHy1eaUJ4s5gJ4kSK4mUKU0NiS7iNP
apoVuXQtcO+CQEvVuiMsq5hBpZMPr0wGzzFMvYDW82ZrA+vEpGGdUDWf/iEDa1ftK0gjjBACeJTg
7i+hMDZEvKvjogda02bbWWSqWZwKcOfTBlu2feNa97RFWZB5I3DSzIA75aJOlAAZjnvsuuM2FwaD
VxAvkzSboZ2J66nLguxYbkKGGfH/klj3gd2ZLZ7/TxDTbjWdRR2CCwEIMsTQxlaFr8nzCrvHl3TT
XDkQY59G0Nq53xwtGomq1CiBj8eFEtN6I5FbxMjtZ2wiC68Ioxurj0DNS3pAFGTaXVz67pIlCo0N
Y6nT/DrDHMtftdP/auA5l+Ny6VJXaaNihyw+nWWLzgxMJEJs0hbAZ+pXNffy9fbA4ttaK9Q8LtLM
kNpOXhGi0Vunm2xuwJ7r0JjlyUENqeI/d3diI7qLIZelUdcbSXfihOm852Bg/8H2s8jgzuUjNl5D
c5LsoiSHWret5Vio5fp6YNHlmM1o9b6coYo4poEaaQGdUKsLXcWti4rbW+FfjRGKxKgVvr2HLBra
5v3PqF/nRbMfr0BsqfBK4Z60W5I/M/RrGumDy+0ILy2zStpLgkuQGWAEa1+LDjYx2DMlsTl7Lq+f
xS0Zz2UhfUOKJpiG2U2K5MNyzfy0C5u1P7ddNzfHVg+XjUg3yMABjmyXmmjgLdBTQf+poYQ48ExZ
KyDn/3sNlxiuN0WHohZjYHEhyOj7F878uvP66sPLB8dI2Lm6XDtp2OBr1WmEbLilZmd51V0moey7
LAEC/ofzn+vbyyTU+0wlSPXqHikLdA+FMqGgiJjKqLkdSiwmJIlRstk+tzAAqw6YOyetApEf30+G
PaKeHh9UtC5t9mOERvmUXUNeQQtJ68uBxGZoGo1mrHblGQeXelbKaC2CVYcr6P4tt7iIZdMIPzYU
xOj/dqTuyzKwrtGg6kiWpO4368X1sW3iCNf1ut0j4an5ATWxj3X4lRSXWKfXC/DjjcYoV3TtrCze
J3GQ8YOd55FULIQHEq8ZvY6+s7lOiSPykPrBdRJVFCSFDUcqN2FzsMM32HO1F6jSk3MSndLlHRab
+ZLQCG/fRDFbnOWU0n/z3dnxAmTL6Agn1HxqkPlIw9BitmZdGceQ4YCmnB1S14nnPXlnzVPtuunT
zTDcZjP9QDkJsqOHa33uXc5WYfiqHDcgep7lb8FrwpUOrofrcfHYPnzx4Nu8PYhcBRPagePC2kAg
gc7Af6K4JKUJpZsmzM7dTWtOguCfL3xY8fhxjAiziFFSjm1uW0096mYRUnMEJScQ10SAmueW9R4r
smx0z8vTsUkTHjESuejcKRWCIxQ59is19yJvq9/QicVvCG/fjlJHm3Yd8el/QtXTHwIzUndKRt1G
q+VLERp7Mblv+046hZ1ueEIj0+FbijPF4tKmOfaUZ81ZK/nxHZdg9Um6hc3dV+aVkXVV8maG1YJz
Ajrca7m8NUJ394rrDGzyeQlTAKUSVvxtqjuwCnGvsHPowj+wshDNheysRLNCGUQsRcjQkfdIZMM9
oUrJTTRT6ZJ0Z5oHIgagENaQpnVVXp3EmNsk62rdsR0jVO/XJygGi2N4iCeSLzTRSYEpGsZsUGqL
/LcZOuKpB2tch7uY59FmoNtRzNoggeu+GZBB+eKwToUJFNHrEqQWt5SAapVE/8wsP2y4EkoLWSLI
c3aVvTnWoTut/vBD4/N8uE6Mnr9sqv+4YePY4tpxigsYYl5NVMvaOecYu4uSDlpNcR8jMTw1fcdX
TH51sb1wFQPvP/YZ05PazM8/IgONa2V4CvxrSvI5PR44FxGerUNh2Xc0xX+G5+vuHeQ/+AzaKIx5
FT/4SwTu1AwUm+XOgmieIGRUcCEvgDg2OtZ8CUWWqNC+6yBQ7AlKLnM6wIARKv1h7FKxuCzewxX1
YfOsN+jXqjSVfJ8hpukIZz+cc1hSECwMtL80Cs4hJuTNKu+bx5usUFAU/IqsrGzNyGgUexqTU8VF
2CDuDxO/oYuPxSdLxjuUptJe3aroVZJv1hebsihRRXahYwtW+Gpxp/LeBaZlfc8QP/Hya9FPZYK2
btZuWd881wVa6+ne/3RgTEAlzGqGyzAtmVrgn7cLIDfC4KAdWSC5LLcGF+yd0fXH8Rjtjy/KgHnv
rkcC188LEKLiEGc3bsS3FGCYqhekygDOAJnzF7J33lHouYd/Ta7mbQmMEYv/iPxzXoG9kda3YL2D
ZyroYFBa2EmgNLrLC2blbtVz4YfCW6GFI0ndjowEFL8w6+zf5HHtv2L1eoZH624Hz5TGMfLOxVng
gjctmBJ2VNxFhS/7aiz8dMelQlDXk9tf89suLLkKW3B2yjfslamnm4SYLghEXtHMYBIZ8gifpbBm
JAWQZ6hGjzPKLJ9ZPMz2CQLLt9C8kpeENBqv3MB1Ou6adfsaum5odAh8NxQNmwIra7yTxv7WA8D1
7IzZxNM00erg+z0lt8a6ARAR0rEyX4k3WvEoP32O66ju7mpZK2FQ8MdGfC0+tQCs3XaLohYMvtUl
spY9prWE9qO4QBbet1rbAezoeAbPuK4/57rFkP61sRlgqsFhKli8xyuZfvIXPmgr/yv4UZ/Xh0Xq
5MuItIMZgLMENWRIk+HiBM4ZchX8oeZ2wSrUs2j6N7BkGbg1ZzkxhSPenYj357KFhWU2FZMuL8rK
0PVMjASN3cBGpn2ZQDhP0DkCAvvJkQGkwuKfPmgXCniizOA4oipf2JmQzo0IDeYQXA7WfgxX2pGT
FvFhzbJkWnqJRosDG7D7df2Pv/LPWIyYr9EPNl/rYqx5SXiT18CVpBfbxxkrYqGy4ifq32Wqdn+p
dNOmc61qqiscWRpp7NsnFqDC/w3sjEblh0yvYp6jFefg8HaZJsPGrv4nqPtSVWBwc6dsiwbbi5AG
glZE6r5orltOV9qcmIpvTiRwHzVyo4hNHji+96R42uvg3o5VKd3hDDPY3iSAZOv3L9DPzxMIFySz
8lnaJRL5MkQ+t+VjHIC6G0j0LZXWKiy53BuxPBTBBylfMV81Q4RxnfpT+yDXSaAKlRIQMCc7SrQX
e8+5+/JOgCOJVlHONqRL3wX/xJzBwkQ/JG9Wjc09fDYC3YcBeMgA8UuNPiosAHhCgRexCrokDlEW
7ZQtI3HaECi+AMNP4pASKyXbwMa7LZX3CngxySvj0nLpbIR126lgRhY/F+3Kr7laXiClFlm35h9s
YmjRq7kjY+xuls9bmZ4In04vA/tQ/ULg5nlWn5cfyHgm6v4E4ukW0znFXRAlujReLCspvIumS19x
D3sssKSS9xsHEs8ARrabm3EqYzgmDInr0HzSvNrnYMa7rkhoJB2cYv2d/7i/NXiUFXWhmGR7rWMj
c5YOa+QpNMUZC2phFnYC1BuCiEMh4jIOq4E5GPARO1PyusEPqXwypYlpqnD1ZKizAk+XvhWPyiBL
gJ+Bn/s/SLVn/IL7wtovufM/VG4AlHpidPbhZDwBKjqSnZ2oFk682aSsIW57XYxzIsOE4KFcwHbn
LdZAnnPlUCYl2llxZkjDSB1pcGxXgx/YU2bSD+pNDwZNS0ohhCscWEi8e7F+SNlBnsTsr6uO0gMO
r8p0Rbcr6B2zJMuKD/8GojG9WdhmDni91HBakubEt68nltRz6pQGZKxz4MvqEvFr1l4+ShfRbV/v
av3iVuMHAvh2Dk/runnZWDqVa/BERdhyCZAJAZQp+uw8LWDQ4QouWjBNMKmDFaf8tmfh6wrQMDa/
2TjZfa/VRDxmL5cWXObLTTz7e4ccXkEjTX3t05qLWIXegzITcipe//caxcCw01Q5AnGTSjRuGTfT
Z9RRfJLszjpXww5amLccsP/o29XGXYz3swm+F/LAVG/PgqnMibvsSnyUlTcSvGv8wJvbgUbgrz6Z
Gdm3nObXcbnIbYMGZN0may40qEgezr/oA48Z4fvILctTW2Z8krMgCym3YQZ5aWQyOyX+76vmK+SW
kWQxKOjdvqLJMmcCFrd1tJlRqZpKHA6KipGjzFq+Zx4SkTnxpdmquiZ3LmNmpc+RHF1eL7Se/3O4
M2Gtuq5zAfvnzikpOn5yxULBoVXLCySBJ0dbMUXve0rQW+7gZMV8vUV4os5ws0nXrC4VFRuDiZ//
ld84B4wuc9BrcvupTfcvhi3YPQq4tyQ7IgJD01ivcvgOUhedYW45jYKYFPou0miOj0H6CwOHExkF
XuqswwSpw7pKQpzdtpTQ0/VRKHVTag5u6Z1vjVKm5jloHgyXH9EhfvJIn7nmT8jJgvbTON/HVifp
T0pFkw0WpwOefRP9gjauEtaJ8JBYAN3lvDXRGFxN3KcFvN2eT2eL6fdU7LcC/iT2U+DZBHvtyidA
/hxnHHg8usLtNANxEjWla3ZczoT9jnFE/M0fdKL3w/SM6aP8HTd1IINOH8IhWxZolL49fdRU372Q
S4ioQVekjTV/tEVqWatqsGwt3K1tQqyMI/rdaSRw1cP7Wp3/KUV+1GKVQmuHG68Z6bopHdfGyP+h
2xR6oCFFzUVOOpYGvYOXCAHdbsAyofGLcRO0TKeyZWaomd5kaBYuZeYncTL0HSLBTAtfu/rpTwJG
JAd0sO3gSaCqOmHsSUlO3sx4ihdBF9gwi69Yv4QDTS+8pK50i/MjTKAYbcTYBBeQWLxmEYhYQzws
3iY7xpOfW702OhHxTJkv8Td03Gkk8L/k1OYDcyqyADimLIc6TDIEy3Vs7d25uZ1tJmulEJT5hdJA
E8kYkKWwDW1p9+J0p4eN8iIjfl0lz24d3hthfyPH9szZuK+fHFpS50I0mrPqNWnYNNifbsb71fjl
A8qbOh4e9JMiIYnWBAvahS0TWNt1WeARQZreg/eRJpXqoMqsU3491+OtZXDyFIkAjT5fcGB98T7S
RrGFxwq9KHhoIAhpLmFIWNG/4lW6X7dIT0A1Ly6NqZwwYZRJbi8/OsYfTjSj2ijgI3JeYXpU2Frm
PahpS4TaW7JJlyJlLff6eCH5l1WwmK/Lhw+GxVgJw+Mezq8//758ZTg5FccfPnv/SlFPKjdiV9VI
KID4/qhUhiCyeM+LnQLxPsiFkNoz4Pf+w2fBmXWyQWYk0kklf7z4CjwKVBQ+Vc+0LeUHaYOL4QpF
s+TCmnzqFr2L40Z7i0SbddwiNjxMaIA4HaMZpzX6QTYx4KUOiarKezD/3iNk1eTrSB0e/4mTCLQ7
uRTcLaGhb4rBCfGyMSf0Np45lDJIkORbp2QbWGzcMcPFGI9k7eMNbksg9PIT3AuKC4ob+LnwgHo6
LA2aMCGflr6vtBYF4PgjUasKJRCwYujaQBGJnPuqKNQa8G8ZH5Cffu6Eph29gake3TVB4nySIir/
qrxRah+i7rXgVSLZdXVKtBXnQHjHAOF7YdmdahdsdUujJwrEm8u9eLf2r7a/TAPnLHzEqaMNJt5E
qe68R1gu56CRR+Rzx4RyR+ibJiroEmx1Z5anqSZ5F8jgcBiC/pfY4WaqRj61nd7mJaJxaK3r8eT2
meaQ4h7zM/dGl4CXihs4EWXugsPv/Jwyst313ZX3wl9TPaM+S4IoEQTvCt35qNDF/ZQ7tsvYQc3D
wYQ0w7SLGepNjyop9VDKcTzfAoNGk3ZhRXN2GpUEhZpq+QKe41ZQfDWgo08brdOsvLhhDSpn1Z8g
LkxEXzO3GT+9l0s4cZZWq4XCWA5HfcuJ70aQ93EahrrtFEMRjmp51uRfLqQN5Gk2LM31OsfirIgm
wpriDU9LBP8RoMcahTIkFl7up4PMG36lJygTPaXtkHOzI0zwrTLC0imDODQfJfxHtePLxfbaArz0
Aj2qiWB3CQpYJTDd6DHavsCWRKvUrWDr+KBecP0EJX0xqLTg3ZxYTRoHjpFXSNu/HGsQgQmj4Dii
XPGZYNdr9WZYQsfzXRhluaSSSevGs7mLcMF8tGvRND2WyV5/pNAbjo9B886b1imKtDWF8mTyOvRS
T7GmZbK0Y4Q5un9bt3iGbddBfJj80aquNj36iIsdd8ZJgmXw9w/JwJHUcZAAJEk/D1WZ6uXLRXqU
HUcE9ZY8WR6rA+xeW/MT6J3RZGpMYzPmsp73tmg0YGL8aivV+CHTnCA+vm3akJ03fPBkbDdnXttI
5Ykm8FqfvDnzFAWuODkCSHL7FpmhcpaxmZ6Y+nm+d5LSyb3oMe4xL5KO81ijQouoJMKzcX//3czB
396FyCaiyHSWVam/xC03FN1lLXE0yJcF5/yGAGn5gaozg1KBUSnhiqXdfqkrOdUab3CUP6so0iZ4
hRcvytbIpDd1y7CYlnB4Ve7y2/+BnHokpCzauv4HqzOXULIZiPpPFKWaOm5SAxfpOwC7be4HZi4j
jPKtHEybZ5aN1BEXUFCw5xHLHemiwyO9wfdm94tKE5gDraQmD3vLK/fvyQRI6BZ0ta0Y8IsHEaNA
5R6tCfsP6mEySoYK6qU5hnC6hlUE2gmO8KqzO53jWxokIc6zIm7JsoMmVhmSdAu7ef7HroSKpO3C
/O3dUDPohAhOTbekZXYLM6HgKaf8UOnah4/iYaCXzm+xlkBCcN+xUaQKgC+uD6WuPxo/pZWS+TyU
G/V8/2iOl8ukU1MxlLc/kEDh21uiPP9bEK6ts2KuAQSG2iWE3YxHFPVpXTa909WxlA58dYH4DI4Y
UfF+SEtK2H1JRt7Z4GIvbntfLf8eR800YNluDwCRMgF4NE1yLOliz6ysidMrKOuCJ3UE7wLaCign
Nys1wzHqfq5K0go6+9UrpWuQZkjqGhGmHSkGybVnt86/pToXh2DKJfFPIioAq1h2LYDN8cxlipB1
HGHbqn2Y41d6eVYU1T9eBHDgvPXw2oCE8hCSi7WFSqW+Uo0PEQWXwTuxoZcmeP3qJJrtcbUv0XHD
geXcF69ZTI0jexmOHVgv6xJHiAH7tF8itegEwgFaT2kYziN6kQhxdhOxv6AkSTVlq4mdZq+VSKfQ
H5BAnCgbUI9G0aDWcmsrIx+Q3JYEVoQTiuT7/FZ/GVvos4/vXpQMMEH3Jk++SMHbTY5J/hEm0RYO
eb2qhOYrn9KB/CHUGl4O2Wd9ZosISBUu+KgmK0U8Homge32iBmnOZD30BmRWK/Qgpd89j2+mNGn7
lbcjk0KhGrFKuCpBrfUhj5hbhY234fTyFVnJuhWkqEsrUzL1/I1z/RsajIsx5AGrSvsmBRxuRMgp
4iM/YQDxKdKp+1ZwNrN9TAE7r9T622XnEKsxTTO/dlVslIqoJo+iulgtYjRLYJBbZLteblDF6dRU
B1kl1tROWmu4YxODrBqKKqvqvcwCP5F8QgwBDrH8mCw/FxI9m3G5B5d6zkoX8Qbb2P1B3ydncvzM
OI54mLT3HXpjpbVPyacfYYJ8Qd4dQgNX4NYFYUkLtSiO9LOhk5iL6npcv9H9+wHdlmGbrTRViMU4
b6+Uq51A0Ic2u5i4l0uMbQ+naeDgmnVtBS2+rK8/hpiraQHNOtflk6M6Rp3iXCiiUefN9haxUh6G
tf0pTh4iqrtAMpMH+9YC1734+3PJJ6CE5MooT6yMKs1LSMWN6rO0hSizUVjejgaLkofOON6vDBPz
qm2ps5u4110qdNlSjDi4Gfc/P8pZ8KdFoCob1iTR+hvDpcVCkoa1XRXgaY13Cz7tnFyNzD3DvIdu
Q4L+2r8pH5TLHdNLcV8i2d2bo2Td/BhTYSQB69L4vX6s5GFnHOCqDRDwFI0K/tPg/QsVJExHkR6F
CuNt6EzucNDdMuAJYlrpcnYkUIqBJ+e+uzCXYu8l9DCd4BMIqYH5P04ctI71cT8BIOS8z1Mn78Al
gfvEq4f9aXszpalcoNoEUS5TdtNZdv8I7PzEZQWwTGnUcQJAEOUUusubzekGqsNKQZlBiyfwXxWn
3Hts2uKivNQ4+HAjSd1jqt/HFsWwzt7Az9zb4yw44/OgGpvHkI9CbfYAwYnd9DYlJ0g3Uk1rQMnx
8fmSMk98ilTtwdtUTwOa0w/VCsiUbrjOd6gp2BdRyawVVg6il6fpkOkL543WeZnBWK1biXzOShqq
s+jGxblm9+QP2Zp4k0wreyGNW55u56vKYincV/6qknTA0Qmi4flIamIKsdAVrXLc8k2e4b+kwjAQ
e5bgEoT/dIjtlHVNhHgxfL8W96z6qfyljgTM2oZeGei2Lh2XkFaXDFxm8J07v3B0SnDqnwNYauBA
FcW6qvP6PE9iLQkGJPiU1+csXriEbTeVvpCzd+IYCR2SRqy9GsML7C2ybqHUOIvebCjSB9GWCDVo
a7swYbn+FWStholA2549KQE6tTn4mARgHLRLezi0ZX/n+6jnphlXzdUxHIfCayteecd2pGHZxDq5
Z6z7YyLonv4fdF/gcVY7cFkBfVYDEvJuf41gXrq5ULAlKv5BhFA+5ibtliHSaJfwwuLHHVV8wOCy
DPqZ3MVabfRqqNBmE6G/KsT18NBcB1NyOPSMXXKOgN6fdwyuVshKnJUIAsS3UDEv0/7tBWKSNLMN
tBNCR4J2ITrdephb9tdkkF20bOCTNdASpvnzYkHgNsDNT0rGgH+AticzbKWz38fptFa/jIAYoJ2F
NsbQWZVzb5rafpXwPQCwb+rxot/+quqs9nOF30Pkap/7375U047Sb9gbJLfJvYZsLBhCSdicBqQG
+QJMy1IR9xlPtB0NdKktj+SCmThGkxfki9X+94X+Ry9cL0EX//mocB04/Y1VfYq1qAYpVVmTunH2
HBpvem7/yUYTV900J4kSUS3iEzhrub/4szEkr884b35d9lRA9reSOy0+FKr1NaL00T5BS67VSVRq
sh0cgNt5f1g4KDI+J6JEYMJSTKsCZcVU/oNpzaYGY6eto30r8OyrAQQTYg63VjKqQdRNWuDaTju3
xjxHz2Bf4xZABIGj1nRR496L4fNWugZD7cSeDAataUWr2LSGtiMA1r1y7VboSmxaNBDxPx0n8YUa
y6lMLS/664+Y05IMH56/3DqAZd6jQ9SPnyFM2PTmxdCxZVmK24Ez7sAqaqS7/UzKNIEDkVhvmdew
Jj7DgrGCuDzYQVfADlfwoaxmiv7m4JICDs+uczYqYkW0BCkBAwC10uuSBkM9aiLsdQhKEFmy4Ivz
npdS/eHreJTzpUtcIin9WB96Y/EoLPE60CwWUremjNjOEMz7SSC9yraY1xNe+g5cnr9NPIdzguiU
Bw1QIMsQMa7RGzPDtQiR06x2qSuVeYLCXUfvie/IrZI5Hd4hxHCkaDX1oFVQbnPR0nmSmRGcRg4O
6TTIADuUHctsmx5C6ILWzHcwPBQmrZrX80JYb73mUGXVtdetvO1F2nMSboRwBc5ZVQEBvKnUCzz7
iVJ/xKUzU8jusk+cqJYhWWL41t+FZ/j8VJeh3/lp1Ofji5D47KyY+ji+SN4VZl4yjw7in1Qc7jer
ZtJo5/gSo9Ow5Jt9AZo6Bz+mqHf1clxWB1s4Tcg2UKs91gORl6XX5uEjA5qAZbpEwXzMsKXup87N
T9tg53vK0rsIuW7hgz5BeCzYang5k5vMQdPe+cjGNo1/sOr44jJsOYx0nej2PMLXNQPfNpqaJ/yj
g4ns2xW/1Wsqwuf8+hIhA8deycUSvZIw2+gnF2BV2MWN9Kn7o4fYtP5TqoIcNFfeuJ3W2rDMhDVL
KvRxUybC2p077E2tIB7oS/RGeSPQNW0PlpHcmudeOb0wVv+HFWxVFcmkLOHEqMaxBMDSk5wsEsCA
5Ed2ZTTwHC3rIrtGe4ZYf/1nVeIqbWsLwuDZ3L2/AwFiVLnfKYSMjVpB00lFNoovghaA0pZP/bLP
lCymgP9zXtrEXoc8iIfn2gVrEG+jl0p6KPqZVURASCJkgfUNWvCm9swbesJy/daRQFgiCJuHlKb9
We8fh43leCYwwetU/PS8DcWzr3nIwEPnF3KTyULSOUaZIRDkbfeUozoNalnbIibMQt/BJ3BZtJuK
2CxAxBa+GTPfvbcLTB8eOitELb3r3CO6gHh2ytpP6K5ETjlIFLkfAoyCOa38I3mY2NbRTI4S60qj
ssbbHA/XU3zojRX6nj9/X1gmDHOZ70NXC25JANKW+BrZyzLygOI2CdBjItWpDPDC+xejhltg3PP5
C9ThY2QCIA75BH/gCh7OoJulXi14X+kgDwwdgHmfyiHj/8Tw33tXY0XPAcomhCeYeGlRMivb9QuM
OEU0myl+wnlKqrbH1iHf3q3shNTVRcNVeqRl7ecvzWyQM12p6QWNnBiP+ESVsUhBufQp9UnRXwBC
s3aYrXWnAkEfaBMsopJbMaDJk0cGUm7MN2kSWqxtNJ5SfmU99lAYPdZ+MOrNuMcjF97BdYK3g11p
wIBD4lVkb+a+96WIcEzZjdz+EInp6+nV41zxYW9OD2/sR6dPU0h5o2zWxPqwD8xUh3jTw/lprz3z
VG5exa8bcjSDiUM0yd+265oP3WB+3E+LJT5VPXgYH7x4B/t+o98hSZIc7YqcotGU4gO2JOXOxpQ2
x8vm1hcM6qD2qauz6ntYbDUmkLO973i60/6ko1DyEj9PJ1GeSzLF5FYM4tgDF7yNhVrCJwMs2c8t
YHX9AgvG6ehIa6rDMTjA8n3fWtHJoJ+icRcYHY0/s7GeGlfqiBT5qOw5y2TblQbdxicCfkj18rRG
m/AT4TcgYQcgvNqcl5Ej9RfFDqqsWfxyVl7VOp0TOfWr3lAz8soj6U2uSLGFgHrnBld6XhDYp5ge
SlcjKkOgRjM85dxd6OCFpvFraZYudhHWwRKeY3fPkck8Z8P3eRzmRjaCWkK/Vih2M6EmxEBBUaz1
7vU2wP7fBj62XXvKYv+u9c0jOcB65XJ2AdNacUkz6msxCm8cMz8qY6zY0SFu+oCEBwApOCgEyJY5
gt04aRIHIj89dWLbO3Kr1ZoA7Ga52ar6ymCR+/bvTH2gZOdw52ruYTA782Jxw2rol3NQFFB/JKWA
1lSi3hDqGqtJIcKfBVis05HLrxygvOOsijM3kxeDPaz51fzmyxuLEx08Tw5o6nc3figvShyQdh/r
nCLvKZ69MkcaliwUEqmmZVYrhCQDKNGJc0/keBHu+3WSoXidIUHtkBpAY49BViIgUPxn7jxe5ZEK
JBFv8Icdgyy0eBeLYMh+mfy6a10MkIaKkoiyr0CGS+z9RoyKxUBkeg/ujyzhhvg00PoAliuzjbuH
zIWXPDAJU3Vxuv4tCp+edoDYja8cCU0xd/z7FFUPgXeyhxDdk+o3jQlUQbvnRy5dBkoCVykSq1/u
2iBoa40MQ/fHjEgEXlzduf356REsuVlYVb46mpVJInfRbsSBWCpf0b0Oo412WZmMgL8C6c4yaGZq
ITHX7xUIkR6JFrQnJpkuimkPN7ebmY2BqGMkcu65KOCgRfPQIHW/wr/lHSQ4C9vzqjq6Nu5XHVKq
EwCqTAlSysuFbw9khCywj5hiZjXQN0t2mOFODDLs+XwIyirlSc/lR85pK303vqe4OPGZ5J1x9+iR
8/5ewKMWn/h2k6YgVZPXQ51G9CZHNw+VyZyD2F0rq4BFxnLg4+53eoRIr8oTd+IzDSRoNor04Npg
VL3R9Za5t77U/1lJjLiCbumXnSWtJGPlCkAO/k4Av0JewB+82Wc0AArDUKyTF0RhGEF4lPjIwVp8
DpzDnZvj8FjkV4JrpxzRfYZvL9qcMMXRwVPdlPW5ASu1dxaFUifQS/flupfJr1+acI7AjaltXTKl
xwbERfwBDKUaOWACgdA3QR4ACtCcFyfGBcvMJrIE6COlSadqTlqhpc5h02GpAnWTIdVLt3wVHUjo
1GOCcNVKXlTLVwp+vFha5IxmxHvXk9X6NH7bixB/d7mM3p1VJS6WSOgVxko6tt0KgLxN0Y0ulXqi
R5PsKXVGNRxAlYB585sIEdc5lsSjd+GrBqMmaQFrvpUdk4Ge7qwjp3jfull4ZbbgcjnLZY8t+jS4
9/BRoELOb48lT3XxTWxTCkuG1LcnX8jF+ueMQ10yYNtBXv3sjc943BRGi8xzBay75WVlel/B8nhR
NlEiuCRTPdJv5KAa4P625BtrfNbv9s8Jsy5qJb3zGxHBF+psIurhCKZ1FQmzbS0+Mj9x/upZ6zg5
TWW4USnekzrEADwiT8oUiSkZ6s8jlOw18kN5e1KQRHdyFsBqWyn4oxYKNtK9euGJ7XuAOpJyAGU0
PytZNoVSPDPZWUHbzqSfc0lKlmf6wbr9k/EG2rHeWBcc84NCtFVMAjl2ttcyxQChNI1QauLCiNre
NGdJfxCzsuJhH6gQWazf6MMQAEj/mhuKzXudqq+Bie2K2YsqQ63P+/OqPWjx8mfrn+o4EqVzFilY
zmxc2NUJOIXuDHWb87LuQNGiQSH3eonDAulP/0ATWgWTEr2X0Itgp/U+fAsK8Si3rN64g+YLVMF7
Tf/PxA6QTyItKoxA3n0MFnv8H82N1Gk1aMuko0tAz67hfUXbfyK8Eh5e3ntH3LIJSxNAygACAGIr
TqQMPWwSb6itr4gxsTOVXl9eodvVUi88dVfI0yZEh8Kr/41wQxj+JjIj77oovNWoJ6LtHTSrWLRw
S1bykEi2FYQPwWx3YVeoL400EWwQxmAUiP2pkSHAgw3apevXXGoTfUPG+BG5H3rLjW7syCT6AhA5
NNMBrKrtlX4stlOFOEl749dQg7GbZ8S3D+VO6WqU5lJeXFhkv8o5raIrPooBhJJ/GZKDTkyP2d+A
YUlvFAGs5mh8D5sRaqeVZLumEGkws+dqQ++/ze1OZ9Iyud935wWRAFLpJ1ZMSrFqcfsD7rqupNxP
CfAXqBSNsQ2xr9kWVRucUha/gTAtVNvlEHamM22tqUlVEiNdYASu2vH7l3MvxZ2oNrJwDwy6T0TO
ESAT+3X41c67EeTBh+PVAFaxDI+CWDxsFxG5oQlcFhJrVNX7VAG+Yow2ADhROOqq/aYWTI0TqOJI
PdedwO/gbfn2o4rjKnj62mKEyRvQfnfHPc5oRIxCYZs7PMmYNaAUuL5A+UJUPHCJSePo1iU4NaZm
mR2BuhxPqdqIK2xHdvU634Q6jvot863zPC7DzxYZDH2Zw+Na9rO0q4hlAWide0ZDHWKzn/ChHnvL
hCgIY+p/8kEF1vx9oGY7a5gsCxDOQejjNAMr3E1YOAqyBys+kuKiP5FHD+J9T122WriV7tTTlRxK
Xq0J61XldM8w2JvzkUNZ9EXEvtnAD0r5KrxumwR4W6Upde2Evej07WpptVhDY408u/iccOmf1kG9
yT0dD8SfFiXlnb9ScFaZQvv/kwGcHVVAhZ6L2/spnlUuUBx/arFvpCDYLwqh/plfBNv6Bav2S6EC
6q24JQ+pDiqdmHD2a7EqiFg19rHQGAq3cJ6SiVGpQrf71UnDpzdNJ5WNaKtn37sdsm2DnmLoY5mP
mTFK6zsH7wV2L0DGvIu1sOrGIC+UCYC57WKmjNgjDCIGII2EhwPCt6jRXopCJNrQaTeRW2gHN9LT
y/q+AVDGTTZ0mw2idFpu7G6jzZM95w4J4svPErxP36L0ck/ieOiek/RDCWQYgbJ9EROmirFgsvDx
gpdG+V4+HbH8ESoEVGS0xnOGc5xidsTOcNh2paMIsBHUopIRQcXSL5Rep5T/lgDcRf2PJzcHwNPd
VgQ2NsxenB36xXQoGKKBWf/tKSkxLkThKaOyvLsAIAS+0mtw9lIZGJsoy2lGC3GHJuHK+TqP2qFg
b3uax6RWb8Xpa2xK/s5Bcxh+S+8GnqQoNiJOkycTbcoUbvUDvKLaFbmEDavcaIcEYIdhXpOzslVJ
XnbrbzwjUPHpV66RFJKEmMti4ksD5C9TCf4VAEN57Z4ItYlf09vdUyp5nNuV3/AMbUTptargDMCn
lO5Z3vZ//qw4gvMn8uRExHRW9Oq62QYj8Eo4MsY5SkyS94OiZBlAPT8FlJUWs6vXD6T8hby3VDUN
VDqoZ9uG6YWEaK1DFV9X9lStAu5tPYOd31gow53SDRE8ReVNWxJBErZK+UrXWtaupKZykAbfvPSC
35CNnFpRlK+7CXnE1tx3J2L8oS51FTnO32Oe0gF0QrzhGp4hteiZlbu/CHOJecuOy8wL2eEJBa9V
iV47Bnkls2nhS2tPXeVznSZKkw4QxPRIaM3G/Gd11etV1HnOt/crVSu9cS5VXqL0KHt1U8qFFTAX
sidIu8MfKTFAt+1DF2sSHus3UAy6YqrZzTFQPo058z6V75r/Z8FkeGa3mBep98oJGD5aqCEo0cgv
bD35gknXiSfaTT0L56SLY/GRm+yvSd0UW/eRaNO0x/b/eIWk3TKAaoh8DgPSe8u7udqY2ZKoc59r
5IqVtsWqXJNGUFcp0/j0DiNJMuOUAN0aJX4fMPhkPBqbbMXgmS30cNluOJKZ0h0f9rUPU7WmTzjJ
wP86ddK7cyaUVlAr2+hG8ijX5o/MR4TDyV9DFAfjjhK+QA0QDvy6YVkEhp+7PcWZ+p2LFlBrPaMM
U310VwclNGsyefNJi8We3f8KGVRRtE18kVXKEqP1MZazUK8K+ApKY6eEXuC6NzDqfcF6gs9RbG5T
f1kV3FT4KCUDGXDVg+Za2oUQOWMR+zmD+JAgy4NHwUwIKaxSAfSByIdN1/MDiXuhmRfsyV+87WSK
O61AXDXXtdHe/aAg8kNHwqXx0GnLjvi5UwQqa7TWF6gGiqmUXB6Dn6Gcqlobn1AiK+9EhUnyzyOK
lFGfExkA/sWwg/1Jf+i1YU17BSLFMa01M4JujlLjxtpkaoD04XhmoMKtCq5kXqD/FWgesGFvThhO
jCWOcGMtx8Aa+eROIlKVNG0HvHFMyMQSL4yPOJAK5wwVTu/Lv2d33Rvq+SOFXltex+6yS7M/GD4L
/3DgWol6CT99WXwK+XEN0lW/aLf3VJUpuQjRT9HXU3/seTBnWbacROrajr23bFTwp1/oRz+SG2ux
p7iQhQlLvtcuErmleIAPZhEsKd6Agj97opVlfyMO66K8RdMhOIi267hQvGZSRq8sAPPq0e6nhTvU
uF5yRGWAIieeaMf/LSdakw4QfSpIAJt0pyTafxbdYjBqHf4LX26h99JJLGuQCeaz/xhKcDjwNUrx
Q55yDUA82yysALajnJtid934S41fHyPQFgypV04QsknJoR4DHF66N9FhsY72P+TlNDYmOaaLgy8B
uTXt6iZ08TWfSn4p5xLAztsBNwPiowgypMr+7BsNCnSozZViRT/C9NA/0mY1pU9coFXbWgoi58N2
8fSRRsa3SQfoLCoFctid+oAfVb2f2THyBoCn5katz5UAnAOKPr1v4eE4QtYNMykinnUeomBfr9pt
FDEae45mua6GbMuWYi3p7VlHQ3oFQM5aCTRdTIfbs3DAbDKtxn4L2adGMKdevwNZu4R0/G7NvsPt
hwk0KRviq54dK7RtvTqxJ3dBjISsjLrkKdFvrPKyk2v4No9ie9GV2fG0EPlPKmMAz6oE8UQl7plp
6ivbyqRjp7AeiilPz3YD4QbChLFuow7IyUQak2REp/BoqXOIHOLUXc971qi9ah09EL17PTozY50u
OBDVbBjNbH9eSPPeM1F5d3cnGKH7yF3VlncnozdPr4/bypOf5hkKR7Ab0pcVwa9vE/jeb4LZOHw7
84K0sFgq2NqYsJthTm0ZKjXXMqIClgln9XZ4gBpA4ifzsO6cvuuyZfGpIMo3ZR2oR/Y8wKVNpduv
7AYUVyYZEkAO/iizdl3J4ZiJY5NgyNJ36Ny+qjsPvtshV3G5rG7MkCRwQym6wNgnabyOJD45S35K
1TUHLB4+WKAl1Xz1STTKU7CSU0AzizD020lpqQ6ZXRV2xPEgZFy1/sOhh6Ii3WKILGkKyaPeJQOz
Ulv13nb/0ekQxRTmLqHspEfqS6e4zOhn9C3AIGjxETVx5SX53wFUrzvRlbKrNNlayWWAIMZntSCg
/NQJg4E2L6Xtb304JZqc1IMLJu7//1a80WxBtkvT0mZ8Z74Hwqx9IOGlS7U6IPQXDPEoihM3uV+r
Eh0M6K3EtiDclqWphFGcnOEoIsrTZFEvTRMuzaSbEH494aMEQjXfY2/t6i8Cz59GKE96Znr53ZMD
xLcCqkU/0VeE3CRA5Um5T7OxNyhTAsPGi4HsuHc5XP5hdwptkWKp4y0tLjjKtI1I/z7mW9u0KbgR
/l4tKIaJdKzHGz2mjfWJTra3fXt/IatIidAGbkAaorAOY8YPOP0yEUUXRhlEPsXhjK7CBrAN3mOB
y+7toxOwAbV32jzRBALOA7/5usQDQrQURqHoQQu0Hs3zFVO6K47O3sVgGCCPvZW9ZJpZRlCIt9WW
+X6s97KfgBAQy8ytjtZkri1bspZ/gGUBHo6Rb/x3wJEw861oaJUkYqpaEH8HqFS/OwWWWLFzuCOp
Btxvu+SpGILyUGSeiOn171tyfZMzQb4V71aVGY+KWAZcsq3sPNVLQlfks+Su4VIp5Rwd3vTQ7/KA
eXIE/R8A+d7vbwLP54SGaUT+LhxSKD99EUYUUAdyRNKEVc9rDwovUnMnmjMOGXrEzFOsTLNZOtn+
hPAPgY8GVcY/oVrAQfeBaRLbo6XF0OluatmDfNjMs9qH9q3ZunfsuH9Kga9MzsBplM+clxzfCTg0
w7CvK/qBBt4wZr2pMSUYQLa2O3dZp2ul0aiGMUrIysSXZzCmfZXDGHMJ50pfVHboax3OqqFc09cj
ynpw34mzQ0Zr5Sx8GuK/7E7e/NZWnhtkLbwsaMLo64PLuIYLYAgbPwmUDQXjR7M7NhDY/v+W5Zqu
SzoXHJ26YnwJ5P73hIV1SDsRJU++OED7gcPDuffCzwyInZfOfwavNhpC0qllBfbM3EIcqpKQhACu
+FQeiZ8Mi0ZEWlTBFmcak8JYe0ClCOlIqpcA7P8XPJkzpoZgKju81Qs0pkVYiyazjZDl9py+Vsvu
H7YT7rrG7W3pz2H5EDwqdvxOcJCYE/MnPgPVIAEV3JPCMM5qYR27d4k41ThTV6aAERekV5GvSwX0
fSG0vSmZIVhnZ2QzAO830MxbVgS++lrK1eg+Kt0jL0pwFQpnOcHMiDpUSFhGjLsjlsc+NSpC+8jz
gqr2tu1jzknzKQ6A2FkaOxbxTkI3Lbi7DRtUWu6pnPjuFYQd5VJXs6Rj4b+ep8pGJedZhNua2Eyv
79sFqYTrUlJ7z6WTttiOwHLccOG0jvowQc2aVhJbMFD8WYWM9LnmflA3IqA+14nbnZKezFwhTEml
yzPfNtbCEO4GaqKXXiWgGgpg0Wfq8dVEBRutBIw3Y2LIfFbuBSL2n16n+B8G1GnNcDNIsm35//aM
Jcflz/ValwuGL4SrUx/tUf4UVqavjZI8ohKxzARKVPMyP/Tbx2zdZI2iNSl4kLjX73fMA9AuM5VX
5nVtpNeLTE8rYZVYR3cEyLXcYFZLc5LjjaX3D6exJS9Z+uoQW+faPHiqker2hcoOGUWUpZqyn4YK
JBezXNSowvNuCZQZYv06ndJOUg5UzHcAmSkggN5lET4UrrqWb14PIv+5lucvH8lUGLt3QRChjwos
rPziMxGceD93338ZxETI9ijktnXwhiTgYvLg9JGeIDu3GKlMf9ZBaJvrtoC6ByXBzoF7FAqYfy+j
c4ri5ugsxu6lW0eBSpaaifaYj4371EGQWJHl80yR7AHgjYJKSUsKWxILnMMFpwYYd4Em5DInPRdq
s2LHv0SdZzb5HzvCeUAgcaw8P8wXtGOt99bq/RN7ABJBxl+Lj0CfOp6fq50Bw9uPR46VfYgAZBoI
kymodvwgiiwBppJFM4njIWzlfXJumKFxBPWwZ7IDOSJcNubVgVM6mmhETDyLKpklDvG/5YzfWQy1
FQw126BHBd3ifU+E+6VsOcA7fgiKogwyA7Q4WttYgvcby4lSgh99KxQqxpF+2zfcLfUhfwoX3MiD
IDhtpkukdv7aF+ozP/bqv93sF83En/blHUNdoz13LaDTLcZVgxhmyYCLnqZjMWNvOsmMvD9l0OL0
vWIfXLYoq9511dCnPBQid62tQd4UXkL26/4iO/lwbcM8IaX4XGp1HEM09/4REm74ckFvq1MYngEt
gKaL1Fhfx4xX9SOvcP7CWnTVBLnk1MyzyVYwZUu4BKFw1BEZt9rxhFmYD2E1Q09CmZBWCb9rxhtF
GERZD4LVDHCuuIWuQFW+K7TY3Wk6YbOOOaeO4VAFvxW1J7Ub5FBpUR1m1xM/uvzqVRxD0oqY1B07
9vws7jd1WoCBUt1S40S0kV1OsY8vSQb72wffRXYXuIoygIDonxEObHWfGDhs0p0lVleRhA17C3NN
Xbjbz6e1kJwwdK+0fl+zPOltOCnQQtP5AiizaL7UoVAxlknhf9auYFDe3ItAPIB8ACmG941qw6P7
6n+ZZWp1ftJTDzWyUOeT/KWyEqEQC9C3YNNgsSsS0xNMHMkl2hKT2vN4eWuNBvc7gpBYXkfqx5xE
9T5xYs2s6Oipt/3ilVnJx4NHtfnBWtvQzEoInT31STTVD8uThmRBP1QY0SKYcqwaIQxxT6+fdsGb
V1SX1nddcZ9bqODTQQq0Iiv6N4P+g+GyB1bpSbT75kQuJ/IwiyPwwfxH5fPFZZXbfimjAen4L/+q
P9J07elU4TOMOeQ6BQy/GE077Etl6c98ExVDzUDtBQM/ePJN5ocyd/NLeKD0JtfJZNF/fzDsMKke
D0e9afnJ57YBZTrJjJ7SDKZnyqMqsf3dXqGS1U3PxCuObn2YFtuyDKxOLtc0xOmrYT3xBe2NSO+4
A6Z/cvdV6Wbf19xNnBzm6D6FqSeyHvuZEhlMwKT35a0hobTSKZAq7w9NOeHixC9gUGpAetEpDHfh
G4NHJBUGL4Y54eIQWtXnU/J7CoB+4wOozBsaQSbyLBANb8+kMKiRyLS6w3qCl0RWkkbRpwtMQMVt
IChVGYeTGyx7pL3IlNphN4BTy4pP4Rn7jzgG/SrouoygosxaxDIGA+/T09IEzhOv86vCS5SWpiqG
Bna58p3+RoMP9C74YXGrgQwfq6njyNwvPrOmGjblzWL1u6eAqBPSwJYGzAJXTc/S17005BAKWAiG
K2M9pcoVM6hfwAUQ5MNVscluuL9m1/U3q2S6kea5eT77p2VsHS9S5glHjpdVbYOrI9RuDBr1k9jY
LSuy14XGzAvu+nCuvJl1xyIhpd72s6+uo1cfIiOgY/zCE9eksOv5+uBzg8GjTlTXFfpcK4umyD3+
kIqNM6rAGSz1FWOAMNg04VpEf/mOsiLMJydsDszwMDFP0wgq10GHQsHbAjq6RrlSi+iOAEnry9cr
XNVRWf7Ztz+S0SSzQ4W7O84FJoIi4Rd5ObGRfWWdiFZSgQc1cTziPeZpMi1eSJdQJ3VrzJmoYxNu
wuqxysKfVrg5VxHX94TDVP8fVuUb2YOe0lUMOnTxKe+8CW0xgq9gEn6BxfoT6g2i18a7TdUh5tQ1
9RYu8XwiG15BlgEC/oDBU8BOJjynfx1UPvfjuJEb1kxm7VWRH6LcgH1b0Q3dO9bb9UGByOa36aGA
jfd3MfwBclWD1DsSGrpg+/zCXd37cT6LG7Iks4QOWpa6NgoTOsvKEUxUY0/34AG6x7GTYugIb3vw
u1pIRUqQrTGuC4DYcwBLphUgXxfjJ6gPaLHSV8ybxJEEvKHo/lpnaLYSNG6el8wb1/E9Pr9JrVp5
1r2SK3z3IFfqsRPOhirfLY8nzcWMhOE1mfh0pSyMBypK4IfmVyNoOGZvmFxEPE8Ji0eD+e/9X3c/
ZhiLbZ/XHhCzFjK2RgymlYDpuUXvM8Hlr9TlOeglzutecGUSAhZQxYbyh2/ztBNk2fCrbYGLaWMo
br3BWanItAK4K0fmP5+hf6MgPEk8QqBcBSVWRdWF+KP4vc0HbiO9O6Lto2ikjQEBBCkTMAxU59kV
1rVfPCHEgB78ytNT1U/smyYXFwcoz4vdWxl64h/lOHjn05Ycx7ZHUVDmg8M12Ykf0wUCHIQrudXH
qkKq3CIF4UDHMs2lnPkhfAgsHwFcbedF+gicKU9jOVivp/XgfbQ4NWm4vHOC0CwxqZreZthTyE7T
K1L0BQNmNOW2QTRaVMBEXs7dIyN9URnDSQfUMOI7eIeLSUA0gJIpqcqcCFoqGNrU3HxKbRtrHUuW
V6xQ/WpgEBwoHurJzwE7+LtBCoNsAW05QJN59FMU7vOQ7LZihJB6JOvr/DNDymaFzjOKKTi9idV5
G5fbiEL6MwCE/iIB54v5u1IOka1f024hP+0OWzEwArJX1MF+tKzwPi7AenN6OLAmOI7fUxR4hTpS
UwFhlZO0bsBNBqm1vC8zSZC2A+G6kbMrHAJaFebvdrUMoaD8pWNPRksodOz1NZkbCZrJhsrzXsca
fjiwakDo4F6GI7t+ZfWH9X2WUvuLJtq5uh8To1rAUu25Q94WD+yd+Q9MjBqVIaWXmK9nNQcH5/Za
WKMm+TXcVicjCGcZkG8L18Ay+sBqJxlj+eydICpDiDFMBv0fxGzcMHGByf+h/Z9LGRbeeKyyosRg
9Wrsdow6maUXIsIlSDJDIZVFWLqOQd9jtPTHUUnmeYHc5MbyG3WN5tp/t+uxD3L7RKAj9KJnFH1q
lqmDTYdfYv34kI5PY1PAEbrXcPki9DDQqKXSQG7Q2EqP4JwRaVCPZFmZ1kz0bYIDbM39MGLs7Y6X
1V5iwj7tuOQnFxgjpO7YKRxdb5iMrJBErMS/Y2tXuP7WeXbumpNs/yCWmqlVcF8yHHd8PjAcHlHd
g+kx+1Qqsq51gxMjHT2/cO+cvMB8pJKGiEg6Hk6u+2HCR2t5+lAmqDs1JwXMPB4E1OMpqIG/Q73l
wYHzoRQvya3E7YgkhrnRft+YnaV4j8+yahqt2jzpc9xGivY88GKd6IcvvedDCaMuh2PwOWE1gVzW
WauWoK7yyZppRf7f40d0XBxTjrW/xZzAmuWNa769nZFqpMi9hyLCD/2YU4BCpsDq5OhatSprofUm
L+MA3kB3gd54z5AGW+msFoQTbNRDjPzYhyfxxfDvE6mTfJE7czGCdKOE7jRI85L3ZCcGTpb0z8I/
Ezh3tmXzHcGgtPHbxYRfeDGYxE6tQlkqh0dWpea0M8H0aT12tHk58Y/B6RpH+TLsue1uhMKtkFiA
WfearoP2fCTqCtPnErtAN51D6aT1pfcGW4PTi5uHlzU4qDLjHc7HAlmz8hE/vKwSBH9WTb0jIZ6R
K7LcVuTsSMr9iwysp2renIb4MY8R0M2t0SeIigoCkJh0m/+cErkUdLrGDdUsyluf8KFcQ1NG4KlF
68LewAjzsJaLuPr7AnTKOZN+WqfT989c/CVq2n/iX/75WTDLmhs3srWoThL4zTArSn2JL13xQjWW
RyHyk21X/LT1Q3YWgKMncW+dJobW41ShedbdMGhASkcmWOEOhE/dhZJhpNQIIQQpViPgsD+mHuAF
X1WGlZv5DmrCy2tadYiG+VvEEuVeaRiTb+0fU5Z/5fpipUoveGhqQZbEZad9Qv/kcamuFX/R3TPo
pQEG1IZooF02S1WR9bsbwq7972CVyxp1UVOU1Z9sNcWNgpupdmfNqDs405f2+L6DfTLh5W2DSGdM
Hs4oGn4OXOM3PJzNiXNpyI8nFFDim1qJDJ/PJU/IvqOa7OasGNRf8qL51My9JF+ApjPrZqy94vJR
0vvtQRAYPw+SMKDvPhAZkM7tIVdHHGGBsedrSigWPcth6JC4bKkspElgpEt122IOOuVNaJziESgL
ddob2aLNSJ0X4R/rKR+HzwQmOhBI9eK/ovyloxVxudVM6JYDAujUFsAXSlrhnf5lllj2uI/zEtgg
ZmGkZHxL3qWO1IaSGM/EAOATsVz4VO6jMPSpYyk7HcRw5ZJmMwB+8vevWh73hdvXm/7fntuicoX1
pEiGKmPTWE6AjpUoQ+sIitrsu3Jys5jTqHFU5uwc9Z9+bhR4FbvjCBR/YwrpYB4h+InwI1rXhto7
hq1T8z7yUR1b16PXQLFvxaXj+1yr8pcoz9OSVVfnyVHvn71cy8hiWiu41Bg459VC0nip3ze/ZasV
G8QliIDBoyGOLpKEELrr3zxUR58ZA3MXQ97UT3xZXcXZVsNWVvp+B+Xm8NgMfBUspNEfvopmFvIS
csgs8Djoelv0hjnQRzmTW4IipP6ktsVN+DnslovKSCo2s8yI8cFRgGoOwJsOctwU4/xdxwfL8O3f
ec4Y9rySe6eJbarD8mWckv7AfkX70hac3kauJ6sOzpHlAqqwBPyHGIS+eBh6Zl5E2XSAYMtX3sv9
jiuiRMtDNuGDMSa6roGZ7bP6zJiTDXJt4uOUa1y4m7vbq846hoZ7nVHe9IIcf/EOvV6oFMTHWEIM
7P3VyYOgKj6kF7oGbGmE3KvyC6UNdZsH/HrIj+uhNSAD08WfMlVeypsa+oXprvaD3M6j7kGhcY5p
AagYT/GmO2CHkRnnoZPO7dPfPHeKNjOADdfqexUXExGQz6sOLl2bxwkI7e+bBTw8wURyM12FoOLM
In8W8sIpaZbLCqr76V4UvqI+2Ve/9V8wJqIpAb3hvawPgnihxefzUEoaaaGUbQL42nKYliYSJJ25
H6R4SZMb32wW1TR9KUGFJ8DBBVG9uAUVgxRqJk9l3ghBs2J5Ov5X4eXagiLL1ZhSrqfth4CvGKC1
AfQYTt6ZAnYFDzCuW63vfaCLaCigF0YMBv+abRXY/YYm/Y1A/OopsCEl7boHu7XAG99VPhS2Iv3Z
S9Jc6umL9vESXBvjXO/N0RDPOSlrZFwgwUuc7UI4FHreDFc+Xy+5C67kkxge8uttMcc0ga3yZWR4
DHyHlbR+rvrePvBBLmFLgXL4yyaAuohDVwFZzGZrid9DdHsf4aTQxPrqLdl0kJgMOuhecvDbLB6X
ASOoECL4rnP1pvHHpK2cGsBPI/LzDHhK6eIl9nViytbXgvWQ9Q7LUu1Q2er5DKuTaXTavcvMPZU8
zmA5tF8O8AZDaOE2eclhhvd6BNglqTvY9hsWYkrVW5/tvqzI8+B4kegVeJYK2UCZu0OwhCBx98wR
yV0QK5XCCoQ2aTMxV+IOL+BNR3YdLCqKqLnd9VZNRG8IGaSEm7O6yh9hh3kwNDHJj9io/Erw8Bft
e2mncIvHU89N6eK/vRud9j/1WYBm/8TgaksfhwMs+NfqRTgi/tuhAXbBYRg1Nx94y4Ue0rTXj2hU
c88UklNbWUAs8VLuDtu6RH8qVgEhLQfMLyF9YDSdX4+U7AGqPVStFbZgzypm6MPgVosU93nwpnXn
raWGtbdHZ/0wON445PKesh70L1C88oHtXWr1/ayRGacVj34tcKqNmNUYiUtBeOYrmk37HnCCkCiZ
5JJ0ihY1k3gF66IIVM/AKpP9FYdM23NzKCNEzXVDT4fKXiOdh9HmCnKHYdo1jiE0qEONffAFXe2S
pc5q35PSoYahNnZ3Czzs79VpoLKzEtEH8KyPH5IZvuAtIdi8CzI0ldfnJ8QGJG7YKV9yY6o6ZBSD
VOlbUVC2ofcpAV2ZvpJzoFVeaQR+A0fNOuw4zypGYIY43DI4PY2tWDOw52Jr3pptyOQf91ShORM8
qB7FwLWOniWFuYJjtnhkKSr8q2niT3B5sPpIliX/msusjVXN0OAsTXwUj31yUScKdKjvG3SnI7ID
9uxumOh0JtZOMlKGVKpyiaXIIA3TYYi5RLk2AxBnkxklkTmm+md63xr06X+oPyTS5t/LfpP1+j0d
F4H9Xh5/fbMVS420kBUj+eKTNIJjrfY/UUeui5B6Ouefc62ZhJkvJlKoGDecmjynAAjeHnt2eKL2
/4L9+h4/LbrxNguIfE+fNxpstieutGES2EZjoNzzwq6YFQm02OwJPtvw8USS8wa6z/bEWXqglAUp
xEqVsymK/im7/BEHifehRooFcREGg45M9Aucqw2mp5qTmGK3nbxiINoRhzXe4JtOANAmdZwbirJW
LaXjOQLb3zgK70ZfEbhov7WVEe3KRj7D+QOIrIfZ4yb0cEEGFNs11KxlTz/2/Jthm1c1ro0Cxqzd
OM0qR0TPCHiy8s6i3I/LbK1yKQ4mhpuzYcj0zJRNNtzOkPHD/nXOJgWZAbdCDAQKHlw1dByqISY7
BYCkXeiAhmBAp0qz28oCnthsh6Ux9eDGKZLFnL37BJedeA/d0LXFiJwPzEg9/MkoTr/UC/Vlcnog
kAW2GcjRBxnkjcCakhEGWXdP/Az8rH8tKGkC8eyDKHjhATNiltAqhezXVCw7NPJt2/1biqG+Ipfv
KynHZhKWdRZ3G4fsFN2KG1UMkhysZDXWQWrZXhBh+fwxeVFvDuABxJk7H6grP2Em/TDMAQnzN45W
9TRFcTvt1N3b5/UQAV50PZhzKKIiavcYOoKeRJlxRAEaTHVi8AuqrNLzRm7oStM1e7JKUXUMN3TV
fZR0ol+eH5w7C9tWNYaFDGcz/U/J7DEqIRH24I2QFWxgenrZ9L+PqV5xqcGFKWiTec/MMDOmlx2w
rOI0y8mdWbrpHd6C3bphG/Eg7RpqCZSYtSn5Iwg8Dlrwdt2F7UFWm8ZpQjun+x7F/wAwT8ONc5FU
00XXwBZgYs4RB/AuKiuA38dUQlm3mhWWSH5JTbezrmfaYvEAcoejvOmjrMfO/3A1epGLqo7H2iSK
e7GvAqK1hDRtn/Lz/o104XGk5Dwn0ktuBWVg7NNG4LVUnbgq19c8yYP9+MDU7bA1qcdfO9KMNj+S
W21VuqFEGfR8cTobrk8XH2qR8Q6s+T0H7cA2uYO8KSvfcF/NxYPkwZ2A3/dhdN/VXAzNjnIBR5TL
doq25iBLUtONECAoiUHz+CPWX8Azd1k7XKeqqOa3MpuYZbiKp4+9j+Rv4KCqA3rnt8Nk9ec3Z89C
jlBSqkfh53JnZkh1EUph2Mz3LC/Ui5Dq9Nlc5N9KMI12ua9mUTo9jeCs2b353HnhffbGm9Cufyts
hIytndCgiDJ+nlWCITIQPsxGaRtTzamSVw7b8T+zktGCT6Ezo4ytF9LzdmD2AxgwumghTfBqrwLf
u4NDoRvrkft7sFGhD5BQHiB/sUnbF4eqVBk+6n+yXaJXTcuxLZxvwHpsD3KVbTV2N0cHWsBG9qs6
lUJnhkmkU01BwMNTMoDT91ZEU9SmLFP6kpHidryBGzsAQE2g6QnYY4XDBWP5O8j+HbTtf+RpqwLO
04nmIZs22uFm5dEzLGC9jC2AJpsl+sZ6l6T+RBFhgH/R2epkkOGG5IA0Hk9sDCS7QaHzNm2JlUOw
bJ/ZIMccJXhQR4qv63v+QyVcrox3LTSNO4Dy0tyRzM4Vd/e/BPJDmWDy3mjMgHgZPhqb8VDuuUrU
CQwr/mbUD+sRtn2sbBi/9JyIvE72vVYLC8ONAYyfdrJSqkMMWh8Jhcx8rh6p5yDQk8gUGW8pa3Xh
/HRXNKqXJo3IpI6vkUWTO5vJCeuM8oMwUH3Lqdf1zZQLZlm4lXEfnQySPgtUcQb+ANS97fizJHmy
Nt9AnmUXw1/IGxQ0J277b5CZEmFcZgSyCCYz4DtTr2htzD1vxb2cYN5HChNmXqOpbo9gaqWOUU0W
lPNLTnasIln2lQBNE0k6yxYrA+Rq+XnsyWc5dEEci+zl54iI8qxwUXyzVaHX32xtRxXci1B7Iwxs
o39eMeLGMfHrzaAv/GX7KpZa5ZJBvkzkmJS1moEdveLUYRZwtXtjf9N82xz/RlMTZk4F1ocH0A6D
bGcgVljdi9WuzK2g2qTazMkGSoMy22GBUgHDQlkqasbJJMUugytZkfdtrDKDK+RqNam67hMlD9N4
/boCyE3eL3CCmY7n+7tGLcSnA+WCckvPZ3uKMvuCCb6hYz0SA2YqJBRJCWRNizqkzu4RknsC8dkR
XlRl/jSwZyKWZMehGYg4H/FH8HPAnoUGVsbICWe2dR7iW6BhohLHaGsXwA7bIhxfxRSA4Epw3DkW
plOAjKtAFADT/+ZyFRX5Qbns8jASk+2ujb03lHXN4rfwkuOVqkDSz8zX0+bD3yrhbFCCciti7l8f
gtz3OS34fWOFdcXykWaTYu+QWbC0zqR+bab6gcWk6NKomXbnlmi8MZY4Aie5or9DG2Z23Jswh91v
2HZWNtZmgdv0e3p8lEjPlkT1ogTND/Y82APNvGTrZq6kzOdNgp3HomKSq3M0Xbxv1Gl4LbtIEaCG
PARrTIUpAjxsoDnSi4VeLp59B1X5ZekVfqA9dG4H+Azahmoov4+cEH1VYFCEKPo0kvd0xfICUtvK
I4Q/iP7gcSZTxMjGGDTNK7Zjj7/qPYXJTxGXhdBrUQJ+tNvDrXejnmlKSQqHxoJuzO3aveN8bRHk
y5SOPbOgRkTbfAdHXV8Mh19bEFgMATwK3K1lvzRkpneiMXmm7eIbWuSaJcPp7OrJZrcUb9iyAZVL
nUW4OBFUkrGOl2LV1fxV9ud4rMbNwGqKNJKDnqnU+tM+uwYH2gRFx4iBKkJexL+GhtfY+Mmq8eSO
pZV0lkpgDmkwmeeXZYBIFJXNeSmgcRQ0nKeCbHgHHyZLnuH5UWkYxGczSjbAhT6wF8nP/hgME5v1
t0ZtowvGMBjxyDNnTJNIEeIX0PGzswMHfeyTxiY6MoqFvWwQDCuYGPNqw7KltEj2iqcDZa+aFEWy
PSMVdH26hyoISxZ/oThwoMzLe6c2MnzXUia4HW3fJ+JujGMHXPR+GFiuT4y2hKqUMJm50YIV+8un
AHlRxhiXVMlkLhDdlfyqO2jgTXIwgXFcmHYLmsp0nERM2i92vpjgyBIDX1UkrISQFriNgHHImEit
1C982h3btohy3QIMIynZnUCCTl9UUfJo/n5fhol6QpE3g2AIntwFi8nqTSrWRkftI0XYnu1KRWgc
l5quxteV9YkN1z6Z4OWT39dN4jttRPj48as52CWXMY5xtxZluD7h1ljUnrTTocEdJiY+cDsbg9//
DkluOV4CBZxxBG7NwrYQitvb3nKQIKjq5nWavIbZOsdJ2unDHSLlw/A3V2NjI2700LS/TRt7/eNl
CwLOxsOSU1LAG1tQxAbb8H8e81TWxL7pVJUH9d87R0hJgJU6c/LPyZHP+v/CRKsmBilrLmYBaIA+
8W/WCqpQIIU8O8uO1WdrULpn489IFlK+pYe1FZINn++bb3LDmF3SQSIFkbelfqCilImYGn59Ifjj
AAdgzJhko0cxZNnBoTNgjdnSOC4TBTZpfK7A7tcAti7dN+KMToytGuoWMrXxo1nGgdyrqN9h6fci
i5Tk6XC5BzZWkUawWloOBrd4PSc/R+A93AoUjzpfjnrSTbnUK/ul7ZDHXDGKY87o0GoN0dpQWbhQ
BTtRuO/7n6B63GCXab2XuR/jxFqYiKcFp9hk2Q/TmE7VLYirEE1dD04lRCC9dVl2IlRTgpfb/nQH
XqZPpK8KKcpR6/94Gb5CBR8Nc+pTFKAE5uRHOYBm1memwpHfGuLKKEqAGk4bJd/iPQcLzwnWpAsV
7k+4AkERwfFsxhD9mLWVZPBRPu7od4pFmDfEmHuxxUHVhe7rPXCXHmfBQ+9FQ4LIQdESfQwmtLQs
RB3uK9yw3SmOnrAw9sbzvHQ6Y7f0j9lseYckN1QtP1TRvq2En3C/DOWReBe30pjBEbqYzDC6byXj
MBxPoFwfaxHRdXmgvV+QjwoY5hbA6WeSpmXpFtJGFKvnWs/BxHrOQ8XzO+B+u2vT4O9pN+txMsqs
gBOBfeKZawv9gsNTLxTMddP4hmdjUDmb0GDWMI0KPRjJQpGuwsCsrfiUdotIF8xjsCwM9hHREKgZ
JXMKvC56xkMIwoyAblmuIVfpgWUGYSCznCL1D0NI+aJaIhdzWJ1rl6Q26/EHFXsKTu3GJ1qQKryZ
nM4RyygCz8EqeOp+bWKujVhxnc1zTV3NU2f3Ery7qek8PYwRieAZ1UoQx9rLkuG2w4hW0lq5LCeu
HxyBEez2+qPyt5zlwZr7cDWuPelo3KLA5ztT3098rEdYDbk5ys0z6+D4bxOHJBfUbMcOpsOTn5w1
dmlbHeM6QLu05OAbDo8ZHPEMC3GQ5KtTTQRQo03maA5HNS/+7DpzthCBKmZj6zpF7a94UMmRFDyQ
cPJWFNCEERNYcp2HR1erEc+B53rk2ISV5EqpBOQEwSUS1COEWW+WAFDYB5NPPRYcZ1WV2n+dDfoc
kDXpAgn8ZXndEOBBvFPE4OZa3Fx+YQP7JdOWxzRyA0JGeqqNj+Zl0zNIkt2vemffXt+WqXBBC+TL
mYJcH1X227d4NYR+oqfxZvM7cT+Kkv+ui+MBzxrWv0BoMFBH0EE4qFQKHssEZ5EVz2zAxh3/gjT8
/pXGc48DN2VPyJGgKIVX0GkpnQ7ygnYfEUc/Bmz1D8lO6i1X5zsnx0dYvO5jqXWgshElWWR6BFaW
RVSNa9AzC6piCSqT5DWQyRxgmQ+8iarODPGP/3rGPCx8ywmPOjjhKpJ/4CuGBbjUkhsnSLvzrl2b
+DZMyIFdrdTlYaLbuYDgODx6oCIX3PWCTAzSOQ3TGI4cnDozMc3vy2guVVDGymK6q5qSdOkOYojQ
xn7Y32ZbDUwwWXpYO8o9ex6/YqD0SbYtEUWA6ZlZrMdwiBUS9bn9u6N8PmjhWz61hIMWAMOdlf9q
RvEl4hKnlWYnSgXE8+IlU9+SutuvN3xU8SwIE/8tfiu0Sssl3wdDgEBXZluUg/6ipuNtBgQ5LnVw
tgsi972aoJiQmOD5e0YWQ0i4cRR5GMZrZM3stDcYC5UjHjjHn924POitQm/CHpn0rpNz14QOnq8G
5FdEqPwNH963xaI0LxU2iWGdxUgytP37PppDUlOa6DnFYTZHK9Ib3oCAJotj3ch9uJuY/tXq5OuX
k7GTBfw7j78S0wHLjSWhShRgEuOnNFbeLPfSIcH3ydlwEdy7lJtqBGldJhkiiOD1Gpp2BrI+FQyV
3JhGapSY3dpHFIx/mFn5KL9fiG2rWHyHndXuOx4JwRBFd9MwiZIQPejIPKyYv9E1Hog0R0ZUoSI3
0hm8VRXIwV9XGJo/2ho1WW6XuQxTz1AkBNvE57rj/8umd+90e2xa+1EtZ2srpcebEI+MxKgb9wZV
I6n85V8/Ia7sPbQSNkdWJJMmw7umtbwU3IMiulwWtqks+qGv3wHFPrpZA0trVHTm1O+9oz3LGicM
A21KAnuyYDXlWiAOq3xF67Chr/NVAKUcXBjOPkpgKOGocCWFxo8dNDBoDlj6y3GwdK6YoEWeXrnV
wLExgk7+/gug1yckFILmbgorJglMLEwIssBB3wkTUUVftNRGYGzbzp/LBtyLe+YCXFNA3FaoIsyz
OYPySmlzfSOg9ln/TFMwA8xPSSKsh+Rb5jUMO5NXbTL8bP5FMeo1c+p5L3VmsjtKsIw05/UHZH9v
YVbprsH+GJAGALueHuZzekMW5PPIWY5ERJydJty7jqqxvzkIrR76+cZ17d/WjnDG5/GjNMBCDm2t
9QR/k/nwV+ehJSsf9ntpJxYQ3Jc8bkg9kSUSK6FgNsTWD0xRxqvmBWQsrBILNFAUbnlA95TEZ/05
qftLQIgHSYyHjuOSHKZI4pq1VUFafjjbmsXi4QGfxXsZP4ea8SeymDI8L9lRPKx8bN8UzF4ZYqd5
3CFYvOB7+suJOT9hIgcXt1rMaoY35OG9VAJGKy24PUiIzU4FBBAEXOtBah2ySi3M5JFwdXGLUpvj
QKnAZi1ulqr94sLLlkkiQZbijSG/I+8BwG7THLRMKZmdXwKacpK8IS9UQRQJnk2i+W/prnuRlqmp
MGJNiMSTczFrqnoiLmEpmF0nK9LfxKVNh40ayEKhwXsgycjEomUGBepqrrUhFZpD7rdEVmQN82ol
PZJir54yaTLmGPSH9CNEkqbfsxeDR+GJ9xIvc4c4mLY3DgLQL5wSN2P3P0+iThxvHIpY8CHFZaiG
oaaeYjpF/Wup4Z/JfFSaTFhe8SNMr/w94Q4JwUpYTSbwIJj7uYxPGGa3eWKMSefv+JmMHLCoYa+q
nu6bHDakkX4w8yeyi7V88qc92KkeflyOBkox+Cj7NLYmH+I1VIU9eCspuFqyhd6jjjIzRJry8+dh
tT8WjUCcUoGLOsZM2xKa5Ir5FOYEgn1JHPRv87iDp0KF31Mwzu0IgNhhgigqNf2nRhuFJH0XJalN
viSP2Sjy4TryS/2MtnyZPIk9Sm3FwP8GF5JEPym9+6ojfKSz+m1equ3w1N5DR6WKWKCNfdBbkW0V
0FepuPNoU5VkiceRMTtX6njo3VIq4o3RI0jzL7+c0TemBolcc8FVyww/nd/NKB+pLhLZK1+rSfpG
S74hs9GwWeDzNDsn+nLIo3VyY14t/0FJryp8DUbnbvknv6l+yHXml5rlM9ZVZDjO4q6NXRyaLr/s
uR+ZlBfTa9rZAnY0fPJPSZtHb2U9hwMuX6S0pwwtsxjGMBDz98KqS6AxQ4aXRiyfUGe8vDDbNulr
gX8mXwc4AFL89stPFz9cKlt25wh6BE0MbNsh0Sz7wyeWF3Y+UWtR/PQ2wI89yQEEbZrM/oyhNUGZ
hLmIGTnral3Ng1uFWyyPK+T2vwtoTjiLiOoQWBq2DXx0MfcFrr85R6Sm+skNHw5EEG9iAqiacvPJ
fy5Fc6eV5rWSkGbS/bAI1YlS5j3cxm5YogtLoM40N8g4tod5oareD5celBVEjxASjtnUGoGH5m/j
eGJ144UnufQWsusoohPCZMK/lmUEjB1H7dpbV6aYCam4ip35ymiT75EmLwZ/bdSINxISHDi51mm+
vwuwa5Mqe/kCFUp4uHVwqhMGBZcISxAMpF5wspFDGiNuG4KmVzhyxPgEJvphusHC2zUNZrQ7DJmJ
0NEuPJ2/uNyMwbGLpV1xDaFOb/chqRXHBaBLCZ7ZUOItU2Su15uAvWAh9kqHs/WYxzJNa67tGn1E
MSNMgCQ6NHieVIhxbYhZN/xLVfAsh5lpYwKfJhNBa6noMZG7YD9ebscD/JtDo5I6RyXpusL2olx7
ONfE0Iqeqg/9mpvP7PZAw8mrXyJTaFw+LluMDj9Cr+kjv1nJjFjmKG24shWTEowP4LYGhi3yvAQJ
Ii963t1dBfC/zLElOufyhJtahOmquV+LcnKvKRtmRwHZ8M+6kRSGOfQkM7TWYCIrjJna8xwC4+Y4
NVjtgvS6c0X7d9avX/Q2q+9Ra6Y8qEvBeA33VS7d/2yzcO4DXA7DuA6eCl+OnJ3ovHWr0y51ojxz
+u0PBdEhhJgvGUf1q4pbyIAAc9OTA+NFW0RN4J/SzYXfDIa+/3GP/nUfWNG6nLmvtgRJYPhUUjIC
Y0PPtlk6i2c+KT/1HnHHcuibfYE/hsy0CdmiyosMDK8p8smtYhOdy5RgJeDiA3w4WqEZeixkKXBQ
Y4Pkj/cZgOhcQSMPVJ0VT7TrwmO/L9AVNUMqznwq5xx0hgMvcvsF9Ed1f0/UaWtNP3WzuTHlIf4u
ElAW3qZsX3x4wNwAJn7ETBz6F1Q4D4UktOPy5/IvAtU3D+WnuDoX9T8aFFtpdfYcxFacePNTGiRY
7hIyCZzj7bk+qm5gCcUJR6O5Ue9/6FSVsF3rFg8NtMOYegiGaXZ/UqRGLVjg6RWmEx9RHyM0pOK6
JzyDfZ4mYHGD4OuI73ReQaG9t8seO1sbqPoRdyHy7I0eXCeV9WZ8JsIQFZL7yW0mJwJy16j+FaP+
MeHfHSq/HHi9cKaW81wE+7JjbEo8EMvp6yKW0idYtJ76nr5XtURQkfq4QykOSYgqJ8h65g7ksfKv
ls4SQni34QTpp9Ds4wy1RQzZrP0P7PfEQFgKg9JqQ+rwl4l5hD5b8kZ0PWEuGAAcr0wqL6NK5f5x
cHavkZ7+B1P74GmxwWGq/9QN94I+aUuIfdT+E0fDOLfIK1Ms8etAnV8tc1ze5IQGLZw3ZizUnY/9
VezjKCOIYG88gsTdCjGPfwhIntotPrnmdo7GL1pmcp3S8lfXAauPDNvRpxyBUxM7gCvfiR9B6vwg
EG2Rs1xO8NqWE7cMg5EN6s2yLfgjZeYjgZP3+0thjfZzlfy8V3/qTUicdHVb3SX+fdx6LAxzt2oU
hMRmVECPDNyNWU4Ks7/My3kQGedzEQwww6busl1aSC4vLNFFd5j5U87ZoI7nZSqXTQB5gqfj3Cgc
duluhwEYrXdAfxE5FaKaOKGWwmlXqBwE+oBRkI3SVgJzlZE9ancYWdPmfsNKOIu56JR7P8EvDx2n
N0ii8l4Zc/39N8m//HTc3Wz4KwFd3/Ste6XLtyYs7nbaMQkPvRNUDVImguCAHjCG40cdbC3gpgZW
7QEDcv9l8zMgZ2+k9GjwbiHH7aeF0mYnEaHl3LzxHjZ2mxD08WWeTO0A9lA5+vu67rAL+PLIEcmB
Vau2c9fS8PePK90RkhxXgvesFf1j/34t5Oub85wXgnz5sieWenR9Ip9aDdJgKY6BdEiI0B/kOAyu
wCy8BjiQVT8IfFh+ymlvJ6oWQCTplOgGA32calDBxMn/RohcGZvwAgaSTKd8Gk4/8A7Ke7o3KU9i
aueXrqYxGaOTUyI9bMZ+R/vKQBEwjMWCM5AaKu8QkOsNkZiATfvCOLkEtyxykN+UonSGE25EXCa+
dOGET0tI0F8z0S5rosxIl4gRupw1BEV0UrfIiakaACnDlVEbHEPWsBWUEp9e2uttGCH/CmrV9OvU
9XTOKsuUK2cjsWntE14kCWZHD5AWtZKFaOjmaeNIA01eNh8ncvHmO+8vecdC9iBllYIw+pj1fA0s
X9INKug5LGHD0Q7IXU2P3sF5Qrxp28Ey047HlIWWQXfYCV3ShiGE+uJzgG6v5OtrSiLH2/kH8tiN
Ag0gef93dGTJItD7ByJIWT2IBja2Lw8240fIm9viP0Jo8QK/W53du+CdUoCzQ+0fMcxlH484VU5S
bIE5r90CX003qTDtiP2Bqrw0+YG8fsuh2wVflQh7Fi3iEEWI+viggtLUmc+3TTL52uarYyUa3qOI
hyqk1GaN3uzBxOY1ULcaUHOvITsRfevJDq7NlGu0Fv8Ve+5YouHIrw8q1Tg8bikaTzJoLLCQwlYK
owBrHPnLEzTpXVtqExdcKMIHaSDfJW05TJwkiP+B9R6RXtWtKu5bUN+RxoCElMrGVMuDwjxHwO2Z
lVagzhJ8CgU3mCzPjbTAQirUrpb9bmf165YI8qjmUx1xMbCGpaDNXPjIfBWAlCkt9pfoK5byp+3i
k6kUCX966rlimmXKwE3fwQ9gDvq9uUZmoLqQMxJAQqyHA+9fjY+RhpJQbnqOAuNKXf6GGZ/8Pcpa
kHkniDchw8N++z1SkSfoN6jlzU3GZMhZd+npPQNUIX4idQEaHrehRDxq/79idSkhpjAOJCT8zCNa
W9f9EPaVSs4upCqexEEpkEI0wsZs3wGRttEQIoMVyh1p9o7IqjEw4cVfAzV6iDN/egiacmgVdlB4
e1EiEJPFRoo+O0EVqLYdjlzoD/9lnj8BFbWwLQi8WF2jNZnDAxZNJLqrerJIv7RyROe8lHIKk15V
g5iw4FeXhAMXO2sVunswTYJTB84Kf4bgYbcU1IJv5GurkLmuxS5NdpSA98dSni+cHW2VexyxVoi8
0GP0jQ8+pS4x+cMKmzBhM8EIl0UlAPWEPAvKEJw4EEo6nsTbQmR4i03LTxQMNDb6g2qmUDI+T0n+
3jglzjIuh8+e61VnU8IYkRx8lDi++lW2iUFUMFzbGX/0guYDynQeXyG0BGCb7NsMLSTHtCiDKtqn
N5Ec8oCSz4TJ/IRY8R6qV1J3o6ai5qc1BWIoBSofj5SbAtkeIewmG+nk0D1fq9BHH/Nbnwwx8S7T
a4BrXgZm/MAFFmWGXxQuBu2RDHq00AGTkI17r50yHL/0Ut/3mB5LDr1UeI19+kPJDs81TsnaBJBv
ld+yK4lVsaGmFxbKswa1cv8HFz1mUC5VN/vBJBi46zWoQPa7R+XQcskJ2S0W2wO5P1Lw3ERf/k77
I1hwThe2Ps/nit+pbcu6XPtEEklViAoyxpP285PKRRBB2okmX8VkMC1vNzo1RVsvishO0U5bJPbt
SQllI0tOpjuehrwsWiBx5NAFRsxeShfa34KRpUV+25CiCWut3VdWamgzwzXeo9I0/s3n/1Bktdhf
CYxv11RvRyzvM0ij6ik+hvKsQFh9joO5gAAMU0sUamF2PVUIKqeVCaMOJbfpN4w6DNRy4ZMibtr/
gzQuMKWdigcYQVfD59jCw+scZAcbqjtBm1TiThHBvpj7FuwfyOah91Ooxe7xl+2cNKWdbgi6ApUv
A1I6QGELIJSorcuDdsPbO9EmlQPIdcuDcHyAvd2GHJjwM/48tISwZNxp46lUMk9wVjdcWOWy1lCk
MeyLBaatOGjzmsJD4KEsYGo9rWVQfoIONmFfJo+O1P0p/DAbi1tzJWXn8nx8BhkLCudi7t5YpBJW
1UWh5TNMS/XzTly8zKuNuAjCOy7bZvgfKbIUBSJ/Ub0yrTYLIAjrwQbGIPZubfPFjnnwsXC7FImH
INhn6OS65LD1UVfUDLUNY7rdSXd8Y7VmRUs4wQH2lLTimlEXL+4cboLrnMDvalOyeaPYx7KlN8BV
TYOK4CyuJ+nPm00oYqi40pm/0TnT4KOh1nxOXxwFnFRLmOCZj6312MChxT/05PQ6+n4jK0lTdJj9
5qySbXPmnHrNvUyk+Eb+v9Jx+PfduvpcJnwRpQjPKZQp9r6PyezyqJ6Sqi9OuKFFdUDNdRTEMhln
pKYHdlpKFzOXz8gYpzPbxGuUdSFwFCDMQxgV9pk7e9JKGxKVgOM0b56WPlDnnHljZHrpXe59T3uT
qvD4mKocJZPa72fbtzyzTcsI8yPE1srLARqYNN2tJ0VYzl2Q50lp3ZplRW47WEyO6hh11l2qw1A+
PFdcETB29o8o7KbRjLgjQ9atd1O2ppO03N1NrXoWi1mkbSexV1hKDjLFyPkuKKbCutup1iGzossD
QG3EGEJrwEYQIWvZ8icrOsipQo5zb4EAMSYntPd5SZUz0goXAcqQHS3s6a6jqYrzyahb8xB42CfS
P6469HAbUABJ3Wcse7sWZSySEy9Lw/6EfxqoUf1lmvzV4Y2LdMvf3WLTVO5gAzHtQk/5v+vYmBEB
XEvuyiUjVb3UhmjOnC9NYxY9jCC6R0k5vNaUdhM3XmiOe1X623L1qw4HM+4lmePWTeRKSOXlOPxL
T+esAly80bkoR4N86tECt579K/mLRymJfBHNk+OvgVzgFea3iDmmqOVYNWFBseGEvcDqpoIILKYz
Qb2R2335me9L6SgK/et0y9FMS3IIWE3qpP3zHYd5iG+kJ44McEmwpAfvyUPNIPggz6Hj1ItcNytr
hyqAmUaOEYa5KBIxxgyLK8cp+PWJBKp7Shfh21699o1oY+2qWTwFy60kARCdetJRqms55B15rJ1J
Wk2mMjdPK+knF3Bd7JufvCPioUD75pxoJ0xGAS15ormawRW/b3dG/vnQz10rn1uuBDtOqort3nyq
6wedh09ORwl90I5mRdYMbciONf1NELK33OkGQmLFvoG8NWbsA+u7XVAq2MYp1/FRsBITPXMrF43v
QNfrkbAsRQy8VX8aj1EM/sx3DIxuPbh1p7Wk9iY+s2dIi2/nNJ+VK0iC9pb16E7Uv5+NcPFwW9FL
lApWVdSh1bVHdOv9vpUcBlsbKRhD9NSylWhKnd21AaaGZTJSzl4LgoVGYMP0u8O+J3comEON/FDI
sCkoh2gXQH9fgaTrkxsE2xtQY6/Bg0Lyc/t1hKJUc+4QrhGLGtKu+3dQ8/GmbP3FbCmIWH3yZWoG
GkuHVEGQz1tv0Y/z1db8JEksL4Ca5pSe35xd0dodEFlEIfq9XAM3++tgRMa55fcYQBqgJiEKZU6B
Oot0QjbtIgbV8rcZboLGXGawiHIL4asc5PnmPk8RbomNEpNJfPcu5WgelSELH2KuFJ1XCoXVoNMc
XwWmjKr2xqH8sp5p5s3dd1kMIEfJx3JSOFNu0wRCFbYrM/wknIky0/X9o8tQbkf2ypO6bAEVsK/U
/b6Or8HDx2bNCUi4lWWt5R09JZF/jfcE5LwfbrZ9qBNRlXFOEam2lq5bR+XwRNtwib9kDPTUZ5ud
kN2e4cqDSu4CCqlx/t47iqifYdHzNPHAFg+zpNFKxu5J+2MGXCE0QpM+bUGpXdnR6Y5a8M/PZPBL
9zI522v3R4rFOToudqiAWpijLI4WXiPB2mCQHz545zEO2TSPyIfANY57n89/Cet45EJXXDZu6KNp
+BOcCK5gdRkr6EjHgpBn6AFrB17W4Q/2FYsxXnpbzluOjdBAhxfrr9wIHY1sCr3bTgjM73pXaf0N
vtm9qytWWW0QLY9lY/9fv3dyj1EeveBfjC3rGyPFzSnL/RVOhI9vNfKfFruR1pCDNBJT0mCZuKar
1PrAF1362zaCsz9JABj1N6SM40Mn4CREXSCe8sB1WM9Om+KljA+uP+zD0S3iTEVWXLvt1LQ8hcKR
ef0lpvWxymUltOJX20o/KzSYTbwT2w1YZFpt9qoq1gMG8XoI0IHFNzrrXq89gH09qAoei8Tqrqtm
AZB+/irrn9AwZFfHNDERwl/bG5eqLT+0dqOzTMpq2gb7WvFmS0FKDKL0OSsruom5poVL2UmSGXNW
/u00CPYpb0BMlJG5y9Yxjn8/wXgZwUmVleRnzoHcXv12MWK8GMttbo+e9KHJoxqZ4Qe/+LpO8doH
t6oN48oLrxuMr3NsOkJu8YiysHP5H+9cxnO0T+JzNHZ5VWb9N3g8iq0UCn8uzHooOxJd/kmmZfzF
0hThakOYxkLcCdTSqWczNK87Opbnw4MXHAmlIr0z268brS7iYyyN118tT86Yu5EBbNmvvt9k3/Qj
NdREtx2qX7fg7h26kuQqZdYmjqiU5XLpzLeClrFdB2w01kUwKQEaKm770gQce6NfD+iQNtLYTTHh
hInwCNYX6V0PUKm9FdPCAjPUq1bHj2VLfobIYHYoylPf5Ib3SJcnB949f5f74PK2dZ9cCHMu4FS4
++q+dKN4aY0ubJWcD7lsYBeAO62bZLS/OMrNG3VIWrzsZeSTekDltYhi7LPED04bQsDrSfk+jSQy
ZeGyPy7XM2XaTm9S300UHmrq8D9ffkhRCb/UYulT7uCDce3g8oocXjOHoFeeI+LcBH/b1qjpZVtD
lGxgTfX9309gECRU0Ee+yaMwASTbaG8kO6dHXJ+iXp0GW7P2kaFsdipCARMtCMTu23b4lwgDpnJV
A15fuaAsivba4UtmJnqYU/gMdEFQvL87Rl4+d8dj4726WI2OcYtiw+A5DcDRFZ143TUN32kXjlaA
6KnQ1RNESyd9DJvKxg6jWPfUCkp+WwD/t+EURcWeJaa4mJCPWu4QUQheUivqAiHT75JGtzcEuSM4
lY36OLfhP6Oc8ony3NWviu5VIYJfkMf2FgvLqwNwo5XL7zpQrEg0U1PCmR9CiWHOBAyC70tU8M3c
a0wmoGhg1eEawJfdok6KX2VFcLv86ug7+wjiW7r12VUsDxNSmoVDBbWJyKKg/FnAPrmfIFpQjwRM
NoZeu/M39fRoPJ52YZdIjdaaPCM5kdJstYqClGUj/Pf3i9k805jvrx3Mr+ILkezL9ap4gGr4Fk/b
6bABcBvjXhBxhF0DtFAfUSCp+2auKkGgPeFBFPjH9BGGPauj4OsX+wEx10aaBl9fTEbHjPjorarK
wksB0rkexnXW4ffg+I5aV+1OZ/JRNty0E8QC2bkdTnGt23gCpW17gXQ1IvnYJHFwtMxrScYBE7w/
hjuayF6hSj8wLb37pbwxrRXIN+mPEdSWbS42WR5yfcMxs0O7Jyv13VhiuUwlCR5Mz5gVTh8OLdaK
pvQtPTmnRBVbcdyEGeSwftGG8rkEDU9f8XXuG4Ye6NMSUpBQutEkAVdd+HYlHkfBNQYALLxlG/yM
ieKZzZvLFi24r4P5tE9HEXQOuPeNLJCScZoOCg6i/f34dKykgYyrM38Y3XMehw4hxRUS/kAStWdF
N9ID1oe6Hn44zPTqU4u47h57jDkHsqAWKTIgalr7ziLktq1NjDojBnLyX/LOF10nAlBYKuVV1Qgt
GPXT/Gr5bpLtUXQvhox3Q9AUMjjHEucARVFAoklRPIgWkkWVZFu3LfI6dvQOGJmDbMnIbyX91v9j
0DuUloAn4Q/zm2SEWfnw+Zf+ovfM0nfaMSGStkt4INepVNFkwUXtT6DpjwxQr4pDU0DaET/3rGuE
qgFMWtrz2OW+Q6S+K1TPxWl3sFgCsYyWPtSAvSrMEzFHgSSyGFMhNQ1qaZOtBzghexXRI1Jj18xw
uVHaHbFp7INmGY+881Hm5Cni7+bWTKm9s5QgIi4S4j7YUVM/WZbWwQtdmSPUlfaumTLH5hFGlQdW
GQI/sXxQatCI3Mjw0hodh/ZU1lSb6YTbpq99yypKF9qofqk0je/U0tNUKZ/O8uynNwxrjHbn8MLF
8A+TUAxe3Ta2GZ79Yo4VGpWxpAsWixosmMMWfp/2aYMxsQjCTkhUtOUckpJCYJQxYaAGHFiPs+oC
p/K68hQc9ZrfNY5VBvtUXnXLlVSyc3dTdEpErDEbr4qcgkydxNlirwJ6/Rc2uCq4Dk8w2mVXfwRj
XLCOVOJsV5DRfG2XwJ4MES3EI5gnxa6uh6z8T6v5brKCzJ1W1VCr+DcMDgoyfQg+yPomw3Aqw+tf
iVVjXA8u4JQwcKaSMLS84DHt492WC7+zAewE0kglrNIdjz48/vEEp73RJHj/3aWnLQA2wsQhKVSJ
3WTu4zMqvD3tLh9ASXQ+cs3hbABDMxAn1hqQC+3C9gQPCarJrGntQf+ifqiVDrK9GomN/GpF6eg6
PuJ5pbI2sY/h8Y7dRQzbupy975le00jyHdV99gxUktkpYnl18RhxleLRXGT+WSfaVhvaB+JAI8HH
fbH1A/ggGDZbxq8VfzFdmt3e3CbYaxlojx4ogxo7z9OyU373iWfbZldpKOaGwU87z+9BL0SiZ4EB
vOUz1KzhAlZU3aAdkQ9Z0hEJI1FF/CiQnJrjcUH9r3mbvnuM/2F6CsLsYMlrQxsf2pHwMdfEtk9K
84tIevy29jNwcJg7FRgUuziAIwbKqIF5V2G5XJ43iF3ULGjK9xSKYyEHYqptw4LN0pPuLrqRUhxl
Vok66+ljKsWr3dpzIcXNms3XRFu95hu3+KVQdJG/B4hMS8YU+EtC6d/CHKue6lCKkogyAdkDpq9m
/u2q3bI4MDgNPBP7f48MxiPRHjtJovp4ItdIzMjGEI1CnGvOk+LBHbBduet0zKzXLHzzyA2/98Sr
yLZFKic+84qkwVE4jWpZJqN1ElA8pGZb3D70hMXP17VS6EFcR+5y7StvjW1IPPEol5eR8o0M/V7d
zeIvTJG9WSVv8y3jvdcUfko2JSEmsDPFnepZXknSG+7+TmJ1sgsGt4grVd1LWirlNyID3/cj7Sh3
5tXZZt2SwESmWNLBiBgNUNghBAixvLjZs3eNiMQ53t4f3LCRlNCRJZfaqwqwj9zpw7mAfLwgwOyu
hyaHdSthkTpm+YG7w7wFxZklUia1fu04Rq8c9uL2HHSB8VmL9Xsimx17qvQqK5X14JCDMSSSryuh
umdkULnvw4jwbQ7YjmrLw7P/myQ8srDDvLI9PJNJdS6Pa7nLDc7q44WZ2h7X3GLXoX5a4OPc2bzL
xEwYC2V674JnIU9mZxBEUUEhNvloIw9LIoJ6E1tsSRHeWjkFlszi/Pia8ul7DLmuXYqf23tvQeic
irzJwghS/tnWhWtPiiiMxvId9gwbgIC5buwcNZ+yVBQzfAvg2ONo7DzUb3qanUxFYEo2HEi9KxT5
GkuNtoTnDihpBBE5rirufbc5+HUImL0PZbMpmQqJobBjBuNXNHo253OTXjCqWr+AlvMtq5KeAJFr
Zvlanziy0vdkFh9uyZMp/7qkjlCUNsSWrtcbHjNMJ6imrv03ZrYEApXnquw2V04U2RuZYpuwwZVT
HLKjgdijTgVG31NbIn7EXmanw58WpoXMDT8wmhPkxR4N08lCrgrBLfjwavmU6kRl5lwgu6c0nANM
bdXZILQpjjsy5BIPqQceje64LFKWChynXmhOZ71O+jxJUoB/LTKsPYa9AMEW290ZqEwTB/hQloXo
x5Ro7QNMj5tHZeCPGR5DNqdz85QRCXZroJo1mVkpTFy21Zy699d/U+GO8JSYr5O5zyvzHqeqOAc7
544I66ZdJ4uaXjRCkTD4HZann6R3PknGKq9/DQoRFloG4MwEOKuo5FOhOKhn+YwLz8F9AKT2AtFN
9nEBm/nABAzjSmq478zy9f6JTFEMfIecCpXRc9O/CUgVehOwj+BDR3FY5sfP66ldvbb1i2fzmJF4
bv0qPAOzI3G3gOJ3NkrBGWRvCMnFeOxQPvivvy/MgcGhhU1daspVLZVQ45vtxP+/jGB56n1D/QZu
dzxjBoW8JFPx9MDFJJYQg0pmC2d6TxRkgEuhFRYj235dOqlGBB6OknLB/WWRhGf2VuVF3WUrC6Zm
yBARiGbD1OO0doOq76z8YuzNsK6sPjiI3Wa9aD75bfCZRGzavMxy2ApnRaysyxUVX81+fcA+WF0y
7hgS0B5wY3+U4PAatyWQGNQU+AIoVqa8FN9vhK6KWIX/CGMoTR/2TKiyW8R6/fG48po5uu6eKXiZ
BEhj4cPKWW9LCkuXwK5MGV/+fVM7NyQCKSqAb8a4dtmW5AeSExQ9fvWMwe3qOAJi5PgsGtyjAk6q
SkQQvE5rPm2p6w3RoRjcKNjGCpxc6qSE6UD6j80y+8UfE67Wtod91m4Haj2NOmb8OQIFbK8kD1QG
fNKLAscfWIMC1hb9VjilGiFA/GJ6ALvxmJQrUC3DctodDsk9YrvClMmYxMQt/83zOLEtsjsp1FkU
j2+Pou61xED+ooctIHS5SxUw54En3bAlz6d+y4WDs3HjUoEV/v5E6hO+hMGjd1qqRvfrPv6HUT9M
cQReStFCuBfFL5qystUNeo8eXLUERyjSpZrXpCnrFwGOciec9W+AxRu5pH21nFJhvCAQaHW1LX51
gAhLGsnY5+cSgzYscMdO6B+c4GPLsA/5Ed6FSPa1Dzj0Mm6JdQQJlsVx/da+jTaRlr/BhJ9Domvp
Ufv+mR0uyvQ4yp8IeCmRHXjN4dW6s44jlIRwPxzKes92tiWeaKBGMj2cmxOYmWGMN7l3NvwS9fGe
OTrbYf2/BuTSmoiKzny5Aq5JLnZBVkPM9LtGtcxamZBgW8DmS4BoR2QCO8SMOerK9KWvAUkQZT53
FJcASBGmm8kAZSBY3I6lMZx+A6UPmMOg6Iqe/v95xBczWMIW6yO+MAwqvRtIwXP9UNP7p+630cK3
7076ioHBevIEEhFQbgKe1QrTWXNNsWMUAdBKAFM3PN0kC/pbupMKL0DLmtOwVNDHtu7eeyHWfNzx
crZDfAlsYdXm/tZH5zM8GkGSUWqAIjyqJS20BdxIizvmcBxpJRdIRdQuvvepApqO5s5WZ3cRRAgk
1Twu55yiqHbQ3yBFg8sB2sqTdiUiS3PhCktu4AQSQkWV0ftUqBejRXHPd4gLBj1QyAquZcO6O1y/
8tgLmQijzVTXe64rG3bj8/RXsKqUVQqIDjj3LU4Nty5Tfbg6obskNgkJrhrM9N+xhgqwtwcCSmgD
JWG+/ITWnJLEmZjQLMj/JT9RC4RADazUTriizzxtXuycHUy82rtX0qD8G4lhH1EMdjgyDZjWUUEd
5BioMtZ9LjlpGjl1bwShAZ21HpMRJ8Zad6gKVGTu2OnEq0yv/pLLccRfV85S6nDDoQndgSRuoMAf
5nCVDhrsIwLMTjs8vxT03q6wq2AD7BvE07K4Gc2S32D5XJiByvx75JWDy8JzXdjBoAveqOsvkzZ+
3N3jFRwy8MbfUx6hZTqZb16Qt+N56E8M+YKZ3qLtRmzMBLg/7NNALgsU2NP0BBFYAccgm5UjSUW9
vGzO95VMvw9NXuMsk3ZfUQFZV+VKRaC7bxyOhFGO5fRQNNvQ7FxGSO2Pwliyg2Qi3UGO6/j6x9Ev
phvw+lraCS8uXccwWcye+S07Ex+4LJXMmGyAR/c1Oyabxr3xDmPhIBJVQxfC+1ni8GAM2Mkugjqk
Dz9YCRTUc5rtg7fmOdDQCCLmxuWkxypVjwOFFtLc3oxwsdsAJ4HgD0E5+J4ixudnSL7UG+AITWtb
e6xRW0dXlSUMoRDHvgjPS6hANu62qJgd8D8M8JBWyHVd+NOwHnEdTvtWgbqaYjgL5pK+XXnrvQhX
qFxBq7KdKyfYYYW7e/xl1rlVnr0KkIncaVmlJBS62QnV9E41lopBqj9TOAptOBNzvekwe9HhXObM
42S8qaKoc9WM2UmVd/MFGQh2AYPJpLKiAHBNQ50fBrYjmWvDyEPol1RoJ9kEUnJ5Z21O4bYhIKOr
YCO2W8PVunaOwSrUAQxKb7O/R1PscveckiWOnLC26JVWUE0RpcDhDlWCQHuIAQjCQ42zkSMYpH50
dQppZd/pqMU/WHkpsK/zqJHGhivycO9kXHKTj8ppdBraEWU3F7ETC2UUOwoFHNdgulv8fOC3UL5A
cy/EfBAXI2hZlwnjQLrKKCTCL0cFanXzcljfFnjBrHZVwGlsNdavZcvdqUYWbPgr/IRmpGXIdfqS
iRJG/gh253sKbEdVMVJFfjJB62FGJvFmZtoOptpoywMXev+LNsrnbr9FjXP2PFEGSoHUR3X5J01G
mTN91nxntFUorsWjzeNgz0lkdgtQts4nP1Wwdw1qZbY3oZDdX9B/1twE1npwL41lRfaKsqiHDKhn
oQeP57nZSDZ8EZ7oNCPuXIsHv07qD/Ugauh9AQOOjeCWPbajAa7CcHFpyExMIJx8itMX1yRBwsAn
jVznjQT6tF2sGfvJmXI2kJ3Vh1zqG9j9ln8bq1+LloaR+2yPrJoKniMxsn4IKB7EGoBFRUbpHSeI
kh6qkcclXIiDGxHehTiL3uWo9vK6FD3Vo8E60fGMRzKju9Vkw18SZhxw/aLYw20FUD+qjrZudsE1
li42GLq79TWLFFlkbytiYf7YzKdOIIoXvvZJWQEzaxidQSa6l0E/vEeBKh90uVVFZ0B4VIsuhATi
6F9S5b8aJLgR/OKedQVIEx2sHc+WSyvk7s+/uMIDfuUAR5hUxLmxndw8q53LsL3d7Z+aAfvZrnWs
BrToEQmH5QK4jUzb1eNQ9Lhk/6bp4MCqhNh3ZpHqA3fBE7mOguG1feFG80E85+stjT6s/aVPer3T
1kfgfbrFfxwQFAWcYOnEf3qm6V0R7S1fApVfQf4+H66EWfbso+txyQxTebVU18Wka/anC7EZuh5z
qVwTtSD0aY6gXNPSr7+uMBg+xSKnZkJo+SeMf1wFP6E4VBlWLU8v33Nq+d3xN/C1mt4nsgZABcID
SInMdtNt2BHD/BBgvD3zT+sEWz/cU3u9UehUAtU4Gy3CxkPSAGGrpXvXyIXatChrLHgSuGmAVEOz
8KEzfNZwvpmXLIMNwoBMbfcG1fsKVwRy5O/yRvVkinNkOFmBPFFfkjQDF0Nby1i/1S3WyUhMg9ha
WQ4Tq9KCrB1K59rFcPJCfwtLut/mUDnJBH5AYuyLsEb9ob3XZgreiuoFMKyUfpcY65fmeEObkvgO
SSBF3kZgldq9YSHWfOwyRf/hsH7eoMHhb2qUzzRSlvoiDip//ADno0DwWSJx/z5xnxEQBR4GJds1
4dKKQsrmtpdE9X6UFyNMaqQLDwEmlspDnlFnP1sRigoO8j5+A931XP6HQxh1tC8BlVGgsqvQ+1xE
Mc2IfvoXnUQMb7a1iUgfGMKoy4zMZGdgcmSonc0NsZgDKOxQpkHjthZoZeIE31iqZekL3x+2jWem
RNLy8HY3ESwRyylnXvvS52TnQ21jfX2IlZk0GjxLEfA6pMCg5P42rllTJAj9r5l5tWnKkXzmGjGz
bsDvH5GBGhVaWGGhulvWaQHnl8s61NIinCb0oIehch2EIgdqzKjfFyLvuzqdHpXVXCed5jGh8ZI9
bGWxbZ8wK8bQY0bKUH0fkofyILbqu/X/22OM66mDQf2tSlkrpY6thhaAuVwKTP7DNjHUggx3WqRK
2XGPqOkq8C2u+UWQMd0x0zk7PDVt8nYSeM6I0o9qUhEUj5sBk3zfTv1lWzck+n23RpiVsnnjxrao
TQBP6Qqm7UZCRU0Ga3VuVgK5C39JMK5vPk0LL0WVZU0/MTzP2vS6IIIJFslWOs6DwL7Atw4TI+ih
Gnb+xDDtSHbHoVOrv/dfqw/Iev4uO1E/z4BN1d75dBwNUP0OCRm+3OKI2RfkYpOgjFoumyimErUe
uc0NM4jDx8044qzFzdj45R9q9aeQFMs8X1Y7tPIulXWOBkjXNhSFnprZdTM42/k7TEFmAv28NKl9
3uVp3fNKHeIic/DvL+pbSkVSlK3dEO+xE5UeQyu/NMSFWr3RHpLBd4OpRNZZiW/XN17LJhVLYohn
W2gdeoSNgKX2RcDQXBqiEuUyASPvvGXSZU6kPCcy8QK6byS8RqMXAYN06kypuDWiBnXo5zzAzMnT
C3JuSgifKL1mtWPx1vWE/+P1S11K74xgElxtSmSrM8/CQLpC9JbMojEL2xgmWwjPW8SQwqSCnJfa
pweAYWt7gs47MkEREyZRH5vB/mDWmB4oCe9Z4oRmYO89XSlU5hLVZb0SL4lODVbr0VjAAhQBsuML
cX143lkr9y+OEb3VZAH+xNKG+dpk4eonXIbhFTCSbnG7AFSekdDmwHn02L5ruuPL96Qe9nr76jiP
IRw9DGXo2zx3VdokVcy9KaL8jiy9JiPpr8kQeTm45TomQpzrjie3FEZA+I2JJTO5paFRJzpWg3uk
IQPZ/BUeVjDliMicFz1j+9KQ2DwcXf1VK2Xm0AK3LdK3qk2RB8VizWDSC8l9xIqkMUrzw0hffhIB
0zU9i4TduLgPgdFmXy1fx0D0WXI7kImwt4SGrMj8jQ2b3Fki5Asa1ylQVqefcAbVbzUgYlU9Pb4a
ZBv4ZydJyXQMJcsmWkjZWADfWzr1jpnwLZHph/skESzrnl6ylxH9sSiyJNvV4lUrQrmbxv6y/3rg
+9QsPNz/5YQTidCsjW6bhk+CZjUGQ1oTvqcckx3RJyXta24qi0B3yCWA84FsDjR1tDUJrfjPLdeK
OgcQc4lGyvA4vz7KQCuBsYGMvkhiiTg8+XmSHjXPxMmbrpqXWE8TxEeNoXiBC4hKqBptv6rVFJSe
gwLm1mobr6li+M38zcXlFfCpBJu/fXUCBQ3Ui4NiTizySy3wkxOZIWhH+vyEWc0x/6I7X0ZufkTC
DbuGYi/RtednSrfUMTneDtZZlG3k0A1yGeySmaKUrvs8kxQ2Ujp750aMV1utX9l+/s2gYjCHqs/4
M4WjYxYBXkG9KjQCkU5XvNY9eJeNTiw7WJ+VrPBdIPR3kKrDJF8meZBztjULoF6gdRDcuaON9PdR
saRV9KBfwDdjhSihjOVlkVGhyX7Y5C+8w8HezEPQ09msT5ulPqF6ydPi1NuIsWlZLilOfoQ07DcF
jA9l+Y9A6HvCQBmLuXuWRg5u/TOjJR2vKHCrNfic0hVT6wR7BgEW/cxtpx5cUjOLsx9uQVvZvfwL
rkUxyexqd7e+h9mA7b3ubs8SUTx21fJ5wWTwI6ShsXbvi6uRh8Wc75su1lO8dZHJu8eSyXcQ4Vm1
S72zlUegBmC9REEPhkqh9mz8G+mJ4YDIRArV7n68chZnH+S1dQ+iVTQv5dvZ9ASe58RtdNVItG9V
tr/irhILDlhVdeD4OzZ2dU6844+AWXuR9+/tFvfjfkJ18B+ufZW14PaDQsxh9QPyZHVMell+iklA
8bgOfi4f/0p7XdpSWrTGTyCgJqwOH5utvUPNiAy6yv99ekJgV4/j6oGw6W3McpDH5DL0cGSZvi9P
/ozwqgC95P7feDATguJSe/q35ivrXVRZOtakC4qYyu/FYvZcgUveGa79za/ucc+ExbKrLEwcuDpD
Y82koMh8H9eBbzRvCjqWAIcxOIWG1amrLc3xwOz5NOLOy6Ch0V2pIP2M4xn1mjywEL0ukE3jREyW
fgW28md8udcGR/XW1pTXn2HTin+k5pv5i6zC3sW/dyCBRn5Y0s1fgWZbsf4evf5gIeESwzJHVIM9
cNC5Fxi7sisFFTIYzhgwabbDjP6KcEf1JMSC+iOqsW2Ewk0IqbHwASvUIImZobrfXX4qsP47yWsV
Rs2/ekbNlcS7raDQe2lOcasf3xoe8Ei/Dhv3N9mHz0JaiDqz27MJro4OxTO2VqBXSbvh9Y0gkvXt
biy97Q8jWZwMNigittrC1vlfFvM+ycGqfviy+eP/pV5ZAW7O0as+NDuC4TWvVIUnYDpc9FuBHwnP
Qnf945Vb5yOq6b39mLN25oXJl8SSgJdLvRPCcvRtvXhWpR2pECdOfXlUC5OsGTdaQm/VsPJHLt4D
zsI0nmakRL0NSAyk47ZlU4GcPAkEvgOww3U5d8so7jPb2J5bMbG88Y7ZNYR5BUa0UcbrR16vRR9p
uM0+WRgCSeOFRNBl9zaJOvty3tR31q5fsyKNI6P2kzHYNP85Mkx7j/Ef237O8AO8VQEmlhwsaKsv
JSKxAe6u+zQQveIosBcssbsE6nbxs92RLTE6tvTtkOJdkEu2ltXfk3NxyPyJr4+9vXD1Vptvewt5
mGiixr+sNyC8wMRfaqIxD0Qs8p6itLfP21DDKDHT9sGLv439mX66E+ACIf/0hGzxMQhAaVNaUBKc
aAtrv/ykJYsm/uV8yoV6m5jBXgclC9r1kTL38EXrOT5bxAcFvqc/Yi04uAPJYhLCyyPCJQ2bIL7E
DEDwfuUAxPA+cWrwLqSyiEueSFP3JZdZ0+/gutL+wyi+c/mGfbw8e+OXJmx7uR6U9tvxZS3F4dxy
EWOUWVgGLSnasQYbdUPOPzG/1TabJ9kSCrUcx/PyhzO0Aw+uwJX2MjQROPXiPdQSCZo3fmZWGtcL
H5KFBD6upmR1hvWs+v9GpGKNqeLlPzFalAiNMwvhfjf6p8ocPyMxoSR0Oh6wYyuHwsK62DP24ij7
429Fviy1wjCxmP264bmAFqjIgBj1bctqGksYW4PT/HHlnVTvs2jtbXhOaFRwmieRG8bvztJCZOyT
ibT6yxaogcrCm/pqWce4THQUIWYfa/gEDc2oGRXk+AZWrLXWol1sv2p111rKGzLcsMr7xDopvy0T
6XTXtC6IkRKQ1MCCSu3Lp1XwuzV/29XjMgvKqeDPGgN5NglMnSsQsCGT/5BLyT/bcpYYE1ZBF2Fa
ysXRhpuTKCGebLJApd4ivUkVACDuRcygp71vSdjrNAFiSzpzRXcioyptmnLjF3f34y8E0CsTSgiR
JUBkzrLTHKV69fhgHgLhTSBXVeY8V3K3cj+ZRODegIS8m4IPQzbBCmQM1vQgzOsWCZLT3cTmi4AC
5O7PY/JmFnXj1HP1sEIrJeybGpdeo0qeQu3386usXMI8Hr871gvwYKq3N2kzeudVEk8GzzUT4L3u
dggfiRJZ8q8mVNqBG484iIbllZGURyfVYoD2RsysOMJQuF2NIwYSjBjG6byJN5FlOwDECeXUq9NF
JAy4DVGnTI1c3I+cGwqAogL3yYolQWiD5MgeBlrImDf+Zd7rwJciPMSy/jse5qEPpHqm3BcdSl5n
eSZbegDxFYNva0aw0WJUb/9AZ8Buz/8B2TjA/lfl3ffih125mQ5JRVIGvqNWS5Kr0Kj+VjgsGvCw
Edtx2gV7F+Lq6AEPtuG6HWdHMtLfBmyQxF2vxbp2mv2cTh7Ij6BYSTYPqYWpyuHdvQShn1pR7i7+
rfXhzHVUmCdb//+JiHp8vkPmAHLcN91yjUkI93JepAdwg2g//PUEi3hAsaXm7KlkqHJ+AMBDeRFY
I1OIe+bbFKtoXlFiwa/cYeWcrBHTbAVUXhQue0w6f7t0Zo9V6EtkDBfBJG089CUGHnteGfOn7K0H
LUHDLzmBTjWaLyL8Plk3aIzgCpptADgxWAoBsP/Xq0AqZpPW8CQi8k2gDEVdgKzHRSqMPvx9m7s2
Lm2DKUhJqcab91Xon15famLgs0rLM/ZXSy+KxLxTzrJETIIiI8wwaHEWI2HDyPXNpwTqIdxHq+KS
x8q5LrpWSwrkNd/33q175Dag0utwOmk0uPKZ2OnUu/alkaKstq2Vi5k5U59TIkNbt1NtNq9Rksk9
twuPCkRM2dLcxNA1SpMyy77+hEIMCJNtGRk6Rda+NHNQ1oZw8MGWHVPOnZTVoMl2jsOEb54pYIoI
YvLUBGEUo3jkB4TKQd87O8khNHkQKJoglMgX9X+0JKgR95QSi9olPNkE4vMwYJHO/gLR97RqkRW7
XKB+Qo3t1LOos3W/iJ0OKv1b2At+zOMCH21nF6Kdpo9E2s10lKSnVZ6LBpw+as/Gc8vwdrMar7Jr
UOiZt4zxrZToyfn3RMmevTmylgFs83kmILMtG45+/vuZRsmzG9B2bkbX0xpAGmljrX0egTiNlb4S
FrmtLOplaPB8BuZv3J9xaoMV8g7lcPM5zIsXnBmAd1QpAJJ3aKET7gMyq1F1Yj/EWUPXl54iPn5N
LM2cJdNM8GroftnmOzOEZ7L8VMRSD7p//fnqQxxZ+ipctHkC01UNYLuAFvNGcjKXJfAOjRiF0D0c
FsBC88Wy6gojsoMzEdJKgLeAm381GhVgsilQeZzjTqG0vbEaxhbExFNCFepKHJcOHkbRQFpLWuvW
HVCkqsOQYraJ0sLeZJVMHwG0nFcQPXwLGYZBhk9wZJXE1ckVFVZWIbdFgAZ486soAXmw52btqkYD
e2v8bJsmsH0RasNEQS5whbzK5xCrEbv7IuEGs1oTRGa94QjR+DX5U/RvwFvMuNsEKdcBciFFUbJc
+oUEi5JuIJgGs5cviCHVDoTCk3sJec0JrFDJkvYwoQENig/ZMClNG328nB7j0a4UVzo65Gy6wNj0
O+63b5UslZB8dxjlhMbjKJboFTSicrkbQaPL4CdP88ISVmlDTljDB8TXTKB1RKyNRkBxqsRlXZy3
XIoAC9lgZzr1DdGsoOFRCjQvvC9hTSMru5PeMC/iZ89fFHfJA3duidjd+Z7at5MuuLLfAil47oT5
WD/da8mUD9po7348ryJI8YR9m30rP6BqD/PqgUikeqQp855fHx+BnWiL7BKrxarRBhDzeINBC7+S
PnzxVGea1Q+irPD69nrf2fE22sowwQA56SL7jK84FVq0gpZnmlYMaFVK05sGrpMd5kMdI1Tohxj5
AnUpZdxKFVX06f2UbTp0d7gsqO/8XaGGFAYIvytbKqwCwM1wU0tisOm5oG69jg8Eso2dZAhWbbkS
KQ5IRf+JjpAahTS1Xp75Ba5f+faDPr3dT1Nj+s3W0Y0JQMesBWeqT/pe1Kp1eLrj18GMI4NwFcOp
Eff5r6JjA6PEpQe5gcEuu0bBTVHLaYGo8Pg7rUK5c1NuMxkIiSL6WXzKiKw5Qjd8rZ0zUbWxA8xI
qr5Bp3738ABLJ2OW6WifjMXiHJZFrDYqL3J3XncMf+aowDLAx6c3VO3xVtaeKLpBn2IIE0LvSCoe
REJwzVUbtynfCE9OPSJlmXcYalJ1SChRNM7Opye2WgEH0+Ary660fRD+Cbdr2p8WFbvQKJjoxg5A
WPLZw5l99R5e0oKz7neE+bbbQDHC68k9wI0cpOh5oINL+SnhUIGhrLCZdKbyrzctHvL6nyzii/Ml
JBswNPtVyB37SYmw9kR/pSvPyrp60azRqqCEwUlLqr92IWEWAUCnBtVDvYqyqMoRQ9YFZ1pxB8+P
P4fWmA/uNYSa/yYr+Sz76Dt39eV+JVDYbIowTWYPcu3LIBcYxh6u/R+NJ1TqWYQMH+RD3LgXz/34
VCXmX5omIGWMyoOHgulECsamwEM4su70pWufq9BFv816Hs4g8XXAiiQ2sMfeUULUfoYsWixnza1y
qqIeWEZEMHUmfFZsirEEPYR2X9O0m2LIbB6JtgD0sI211XPdaj6U+x7aeSEp0yV8jLjKb8hRuFiH
7onB8W+Laqz/PdpyF8gXf7a76kgoxyocIh97PiwJTCoWSf9V5CypuVS1aiBZfjNxIdgj/uHM++Ht
E5g5FF2aL4bwBPedL8GSuipX/xzdj2hvadZfFGUCPY1rthpUYvYd0IGPWB/JpZ6i2hDXXZkIEMZ3
y3tzlRqf7YCAEVcnfC+N2gGC4KGX8mgKIE1mbg2ZqgDRPqAF7JJiZtOAq0yz+3W5TlnRPTSXELPY
XrfM2npUr24UlGg26JqqoijXHNu+DpXU+Ku9zxZuTv5ufLlW/f+Vh97Ukl2N2A6HhU96QlC4W6Bp
XIYaDv71osEmr3qHytyxpCBS+M+lv2H93bu7zjKNmN+GDnOruEd8TDHJgEOv3PuZ44T5mFIFvhbD
a0bMd9L9o28CQpFYKzvck/V+0keVJd8e9QknACevuqt4Wtxiex7qHzX4p3Wh3WOdaHabx5Or3SNq
FXgRAVAg1cgfhWC2UM6KaeoEmkKOr2LNRwvlWB6ms7EDphW/CN26/AUby6vjhVuF/RekkRYRR77Z
hCziXbarJCXIvePVzXrcMdnslnXGSFtc1tZi0Vr7tnHkjFsTH+pJk3Pg6WU+K8zLRaiI/V9JpRBp
alurQ4FBR3ZbSD14j5awIIGdqEDXtUp2IVbSe5fGM5ixx0WdLU8HdVi8Tok4v0kJ2jx4s61L+PSw
rhflYz6ZjxPxNSfB47khtv/giiN53EC6wjextvEeUkMeJY36QtT9QJtLhY5W5UGoGd6+b8P/jg5C
8ZjmLdKUOckMXnJGIHSXZB1Hw5OcgMtqrlbiAYRZt+3IccLJJFpZRKew/xBYPyHw3XS/g9BGWfsx
5Q41DDz8tzdCeZlJowwvuMFk7RElwtNu/UhYrNz8SLiowrKFx/VYePGXulloWvXapNDsYsjrgMR2
UA2NGdaLQ6QtoSb4T/awBwLq5pLwJU97KOhluOUf36EjOxUxOTVjL3KtL5WCD8COp+oBaZdzizPG
dPCCWkIi/lAALDDvYjTJMWfC6aoLtYwhtw9tXNvIjXHD/1eUy4HOEoozALxqq1c7oGc8I5zThLFM
sm7Gzflefc8C5ZwnsIzfKlkEezL5RUNHeBniMJ64CdNh+bQ0oktWGsQvis3XuIqyC3KEG4Wgg8+q
P6w/yE/DIZm+ZnQaR4P7eCuVVABhuPTaLxW/2kCk5sco05wObrhNqytYuRTwWOHQFkC3iYjym5Zw
7NtavFlvCvecKertWJNWI7D21FZpDpSib0v74MNDvz5cIcxyT7B851CS86NyAz9cTOUw+bIS6bkD
3sQoEonhjILBjMXYD6a/KaOPqVMFd07M3e42Cuz72j+eJuH/HVauivQDPRnlKCsH+IssTTFstmE7
ycPmaxn4LKnU/gRZu6z2KAnH836EtOoCnzXS2d+IR8TPxpstkPvE00vNzkU8wy//X4Do/yxFTupI
cQ6QkxZbB0JZ9/2WtpP2+ePTLHRN8YSU/lvg5VG7+eIMiV4jPC8xtLiBAnvQjtpBQ+mX8d+7AoT7
/dnnwSIf5OaEPXHZkH13bLG+lTJQY3VOg/lT+xpbWuVxm09nNX9qxxVzqxigN2MuX38ST1IyywxB
tUKrzaWxQhtmZGtcb/7uIrcdTx2H5PFKwDYmrymIzmUUUa+0WAR/SrN6yiwoOqsca0qwZbNp19kZ
ZJatVKkgvRal9BXjh2JXFhNoEFYffzFfdIIClz+LmvthOzPq8ZibWCSGBm6atwZK6JMehKtifP4e
zCEH3Uv+prvdhW+1Td8u2HtrpWAGaRPw5r95fesGoLv3Fjg29H+zw4kKrKm7h5B3NliqIG+Kzcbx
oBSkJ9JP8tiNjb38wBC/JLkMhmxDKAceyd35/0ZuQf393XTseCvdnILOtkxRGokFW7vO+eO4IOvv
3FOPEnVPxMj/x7nfQ1AQECeOoTyI7mXigBDfuNYjDzlNXlxbffMK/4OSlb2H2UhK2EdwedvJkFQk
MRDrNdx+Fkg3yxgJysLN+p6cAcYe2c4c7kLg+nUbCrqLbEHmDGzNm9y9nR+B3PSCCit8muETETz7
bwCyzJV/vZBubJ/r1qEmQiPNwfAlqNUwi4LfR8XgqkxdOBZUJHm8z2Tpem3JY8VzOi+IaAx7PKQd
F4jzCM7CwpaOxIQyCkfGhRkokIY2J2t4coTQDczOn0S/l8bG5qOfzWy6mBgnO53oADBFZVhBY6wv
y63fjkyUSc48ZcfpIdlEDPLOa2gn3i9gtKHWk1cfzwdW4xSlFHCh9XIEXJeOef6BJetK5rhdFvw4
cZPi1guKQxcmPnQKw+sFnh8EAbBePbGHsBzfoWZ9GCTD25FD42KwHLlW/J+rPD0iRhx5EZ0Et0IV
WQzYAUojD3Nn0LxsYsGZbWpZ7w2JQsDPduo4TF9O/2zzxv/AQ0YVvwLxJIPDKivYlYWoL1fUio3l
aCMnSWQ7L9MWDrOeR2jrEumuwoMzDqqWgX3hOKUD5Il20gKcz/aTT5w+vNaAsILtZOn1Y92ZZRi2
CrLaVJq6rOf5zvJVhrV48tfpqc8kzcGad6XeELhhZSE3ucu9BKvz1mvoGzGIa2Q0Sh05C/HyW1Rx
LYZ/ejdbuhRJXT2xyur2Mj6tsaWnBnvDMBvK1nmyjdv53Y6khDeAEIzDvXlelWX0Chbw6UIa4bBK
k/yxGdxCy5les1PhY7YHDHZXL/msmExhH2W/AT6lXgAGr9XZ8zOxSoy4/4Mik801QHlj4iJ4sFH4
tsWlKnjE5GXPzGNOwGilZoGMMhCRHVuSo/l44VK91fDUheJrPe+PBVAPQ8tOtAmx54WpvGP0qXyG
1AwIpZPskEeVLGAt7EC8Lv2imEhZFNRR9Rc0QlXZcXtmp183WQMCZfRtB2hNe2usnGvS+FOksenG
253pWrxATBR9nxXy9NzCsisEnNc6ZjqjXiD35WWVBrILoWX7E8dBK4LjfU4lb8gdADjkPqLurspc
gnVz0h3fNWSM9xGiszP3gyrjkyaOJFokgjZa+L8hBGGPco+mQ99cAz4asm4/DrgliqG8MrwEjzjX
eCqMXG+ebxYMm/0+NPQH0/MQ6YZfLSbyEIO5oembNpSRWJIBP9waJI2ds9gZM61F2s1QijfxQMco
AJvf3PxuhABKOHMzkhIbpBXeH/Z0CqaI2DXGSuzRcpuO5hKWQfS1Q/KWLwAQoXyu9If9WdmWtJ2W
JqOXfVRLUEicaZLn3IhrcaofoNAwQgvAN9Jic0VdQTaduugSNBzaGMOrytHBSz3PQH10a7ZRKDbo
h9xNwkqc9BLl6wpsHINytCySURjQ1fCmi31mO2SkOym0Agl2k7beTBwVsZzIOpI/FGJEMYjzesAk
xxbruriSkEFszuC71TefsJPDXEou6MMhj9YnOak2VwyC2DFOlQOt1pmOs+v8WIOEiPHUCWNELco/
nDcuE3Yu3FICn+RdKGrxmz9colcR+O6/UXbUeTj4tXMeQ948+zBGk8Vuto4RplcuQ2yGgW0u1A6Y
VryH8wkFUuyLePo6/bCCgZBJGkgM2VcdaFenm1dzVxt6Q3IR00vXr5dzYh8iKImnOEcpAzR6eKxp
98uUj3TQOY5n6eP6eCG+Ratpr16yTLQoNnPz6ayrbXCkb8b1JJK8klf+YtNFv08SRi8WPJs/uVUN
lbUiELrRSglA0D92MdLyoYctElolvnRxsdbeEg2wOUebxwA+6uwZ/50hFFd5Vcg/o7spYITn1s0u
ZOW3G+PXW/3CxuA0pDfffXHAZoTEkj9MMl40SHflpMctWIvkRhajDnmAEBi8c94xcnafv2aCUXl3
chCLQzLbn8uNDG+yz0FDE/I9obbWuWJ/ers7v8n9QT5lQBw3LazrYLFtCLM9j5kUTNG4no+c8Twr
Bh/351KNkgfuixQtukG0antis72hpYbZhU1GIRj1klEfdDnrjwtkW7zJdopwql+hARgAy6r1yZbt
C7kCBovY5z17OtjihrpOjehTUj91kCKsehcW//Bq6poPNTpLC6bRq4x9hMVmvqv+xM1OvRoprb24
+OyWWZvwLUdnxtsr15yUom/ol10XViA0legrhj/yM8vDmr6Tns2t7DAhIfoC92fQh55HggfwO4vx
9+0aVQnceIXnQextFKvhVjclVXLzMrYYin/HnEs7KFs0FNoGAtsHJf/pXY5BkcJVd0FpfVwifJt2
5gKnxQVyQkGaK68truSBYFOaUC0kdTC8YApc2+eW9xOKc9Sr1yzuT56uoiKlTE7K6Hc79fHUkTsx
9RtQWF6P8M6QLVKqVTmYcck+TWMHmSdEU1OwsFZblAnAfQ9LjmTsmz/LL3oQmJNilNXqaH392DO6
RBmYgTIM64HxXjYkLdOsZYVYbu0XnovNP3nKS8Jdc0FcnrubV2nEn4fWY4ivgzaVIyKyVWY3QyoS
yc5wREHW++Tqv4EA/2MVTs/bfMChrFnd3V5swqIUlgdXmowFly4xv85a2/Gb1Td0vyPwM5QT7JRj
Pwn5RHtDTYe2vNuTxK40rx3Cnc29MwPul6Qhegcb7icPRoq9E8tHSvYwR9mwRSZ2cwpPHx33tn6F
xf2lyVEbsJidI2M1dZV2KJ/AQPmHPf0zJVt4r2BjIFKCmKYQxVN4xRSbzIYf5WonpW4ZQnTljXKf
cAP1AKoHVtahyzqM1MGs7TR07wZudQ0AEKZqlmLv91WkC+PA4DDCUW2wRZTNcCkwikG1d5fo9CY6
ZixYwtBcetk5OV4O7In56gLqtj5vfqmQSr9Men8tKrY44dmbmNm7PISMKLsmhroowFLToCgpIM/W
/+DKVcstzgUJpITZyMMljSSOXLuoLdV5OeXOldNOVP0l2ecaxbURNvgSFK2g31W89uxtEyYBFwjy
Oh93vVtiFFjcgYmc/fjSAcEceBdv6wOUOuxwd/wfkUFcPM8XXjGlOnqw1bLe55FTrmakyG55Pczl
4IYeezjAzs4mbIXLYfeG/CNgKPHImx5zEFMMBneaxjEF98oyV8wklUP/Q/j8jQHQRZK0l2Wqkj9s
B4aJfQ19isWO94ES50CXfLOyfURCe02zpyrmsrbEPrPQd4FZdAJ3i1ERM07QY0xME7WjnO/3pwZD
bsfwUOhiahF0yuu819CPYr/BMYGn8hsGWimxSI8GFEfflRYqPxIWZRm52m4yQhTytOTAL+M9v394
aq973ymDamIalmvehDwW/IAmzK5qlmlWKx+TOUItuMTkrfMgvJaigmRewvQHxWKFNuVxtq5ILNIE
rYPEyN0bhigqGmIgLr3b+aVgKlPZ3HLzByhqQqOnNNofEpVO2d2BexVS1e80rCAxVLd6lvkLosnh
N1ZzFG09i0TK3BFud2JeD0gbeYBZlD84VUQ/iY14vmd5vFob17j5UEhPFZhLPtXSCyuVRUfj8tBc
5aCg6+bMOrNzyWVyjz6OFjkEnkAmkYU398hbH7pH3+R8TyvqIv4WJ3XBvgkMUsXnm8FtnLuoLvq9
9yayYY7dEPMvDXy6efAEsQHQjJ2Vh0XVOqNQhWdGvG7dLvVdxX3yJW44wk8zqJqfvxmNaQ7yNzPh
3rYaBxj+M7ITS9Fz1a1+YzCzBz3PhVHX6ADNuCJgirgV6clPavkP7NuyiNc6hbKH3M5D4d3yfV07
MraE2nahn+g26ZoDG3F52kS3sem/fK2UCPsKxWmafxrQ824UtdTvq8zKgqV4FtqD2yQL+HsfhLQ5
3iiGjHjfgbkBO46uF1ij2BNk24QWEXQHZHgO1Ww37EEdD2FaEAPptLAFf3rGww6ZtjINkcloejXE
scJ/G+SMbTiVH8s0gvuYJtVSi9zotSN7bJS8AeFYOFBi1SJsWABN+icI5ltYJk1DGfxqBANmeywc
15sS8zmzJLdX449LwLISYLeNXbcR+RP9oc2PSb9H4KuaBmy2U4FbVTMLbLvDunv73kZ9jCTzvVtY
QdjvQsgNe0x4a4NRqWAmJ0B65fRuAh3W8ryqp2Lra5v95N2zUAPIoVYFeHNNK0ahPIiPNgmdQIxz
SXajF6bDLd1e+Byp6INkzUtMQ92ovP6PFA6q9law9UP2HdKtPyAj0XqEnsvYmUmEqkhR7GA8dZ6p
h+DEdsfuBhMsPpVZc9rVbQ3ONxJQ1e/8NINVzgorWo1B+GxzO/PuJI3FOI5hmE67n+WcUmKxn0dR
v1sVBVImPOinaqz/VfEZZRm9B7Rpxf8chnFKs2hh7oSvzgHXpjqiWoewk1u++VgjbLjILViZ8+Y6
UxSR/mrS/JDZFfcqZ30SltkNNo7wb0U/QEBRQJO/qzknTvnz5hBCUNDtqa7bR2rhotzY5yVkZ/66
OjOz9f3XbKMFI/qmikKK2sbIR2msR6Lghw10PCV5jvdXCSStN2KJ/g+HMYVd4NIyKFTfQ1fUTrQJ
C0ee6aAi6knLrZwpr6yO3H5gVxFhAOEUn011poK87FSNtoXGGr8wyMf6kf60/qq+dZyuTzEBi8JT
1LvrbmTqsIpDn/9t1ISKZGil2ZadnvwgOAL7j782LchnUmh7g0cEaAEGTiMvUgstF4wtJxwNbe6s
XASEjgItQtkCQDmN69H3gqGNvSQDdgq7SkUbOC77EBvxnK3rHWidUlnJUkUqJQlv+F0V9EjlZfSS
kw4UygsN+zQfPswXebb3Bb6vayfwzeC/OFAJcYADa36Z1RdEEX91wpd6+Bf0E+FAgBRuAIC7WwfY
NtS52vkUsyk69h7fjwrKP8rXwAdw9P8vg8Mz6oxeJzqiMUmvZQlOz9JXQK9eue7MrOnk1m6Kdoqp
Wu6wKJ1QyNqLgOpQXEmq0yqLw+4zNdLcnSYltKwCASf2vcJjW9KTbi/gqynE00zneuOpB+tJ+4H3
biq0QBnCWPSvs62iM/3B/L7YOxvaCk218VSe6JnHGnxM5BrP3h95gWw4mSPk1uH/MSCgb71hldo4
btruM+YLKo/7E+3/lhnSsUvN3iO6EJneng4aMpbCbT7hkNyYV92E0tVVsP2Wxl+R07uGMOykD+Jx
yu/xux9Bh7qyAboDrKEyEtYflRDbze2SHsKht6tqg+ECvH/q2wqviwuA5xuCSzbVyLI4PoddmwMK
xIokNVRNrxdiJr2GjvGpUHMsiHFpsHnq2X9m5bc7/Peem45KTQFuUOHhLhuo1GBvNSh9+oifQzoG
XozwFt2mnJMQe7Gnc8fJ/NgyvrbO9mPUshHzjjPqHAh8X50K36tjTzwXy4P3qYA8f5Niph14emGi
38jocfPWZo8nO+N+j9O8J8OgRORmtYmlDecdd7FeODgdzVkI4BF5dZLFPbMeYTEcFtFVx6LjRyJC
34L1QK7JyJEPcTcLuNqeT1lufOe77yxolnPfaE7Ldbucft6i32fYbWNBo4Vs5dLDO6n5+xbHlu/j
1KM6zyL9P4XgdQbHhW0CYFm7+R+u+9v+TO5yjY7DbvAXpb0Uw0qdhhviIvQXAgh3HZpoTWEoa76e
ppr8ssqpfXUxOBwUmcFcYKQyYsp2yUneN1ugkOIOXUC2yPidg+diABpYb127s1RaW8SO1lLWerPv
1qcC0Eihn7OUWcrSeKlw89vqXksD0p0qPtwlfj84b6gXGavYMEGrl23KQRCTN5jRffkt8jwEl1v2
5Ujd2Xyi6uP7w3XoaQU36X1mbxvoTqWl1vEwwBkaSLbE4qu5v87XQTa8Im30+VgBgvMH9Lq5IhOS
tfGWByVNd+t7TxRpSdPiHltA+0zlWq4WnCG9bLOZo5e1i3rLR0P96rQS73HL6YbXWnXRMyRJ4AfO
KKm9IiHarFYSciNLVSRVYQsTC9xkLzP3gtlp9h19oWoP3ocy9gI3p7T5PK0oOmJiR6xWgKlruBAA
5Ux48CKr5ZFxg5yFhXVe3OO9of4RB7VqaSboUT3eEbV+LaSGczT/SvY/r64NfDN7WCUZ4lEet+kT
JLQ+JIn2iYXEm3KpnsAdpm/jO28yi3pdizRdXYWNiLsjLE886t68TtEajkE46xbtTrLq1aQMLzSi
/U8J9kTWs19klJRztGLSMxSBs9Et0SKb1m8Pp4n13jL/o3Ih3u9qoZuuEAZNX3RkBLZsWC5n6SKt
11tqPu6qygzLWv00nZ1uszrybhOp3JRjBnylB584W8YwJ11FoYJHNwSy12ZPSJHqk0b9d++bP/51
0Go3W2fQ9qkEu4GwhQnhoTRlAPlO7gj1NGXLUpD8so1TpBFrA3TMuHezHHh6pVNAGRDQLPsuFaCk
tcOENkmZmN0o6xoEoUw4K4KTeQTw5xmATTkCIqMJ2DDUJ4UQiWYNCZaEtDvBHGn8K7tattFbcO/d
tTZ3f/Hsc5VKXNFaLc5ln00vuaNmhIkwhRcvm6pwYXRnYesPaFmXfn4vFRjChmZTJXdqB1EcUJR2
fs4BuGY+4lQhuamGXIZ92pENkk+AJx4sBpfaRW00vQL5eU+x0vtezqRf6N/kvqpR05yuZn1k8OCW
e4N9UNiPIVYZhal3aDRoYUagCXgKEpTya8Hha0rCA2aW51vgNWLHnAGUNZ6N8YUShDnNDvoUnSXf
iKyaGVpMPGRDQoUOiegav+tiNSvIqYJJCukAnRj6htpVefrif9TIF3YelOsKr8v98j2qGKfoMjdu
aQvnyjl/c5hyNbiKNlEvfwv5Q50AHNUZPGNaH4KaChOS9bA6U067Ivj/8vv6n7RK3LQpulYUygpH
gReoME9R7IjnfsbmMNWAme+h6PLYDwGGqiXbk+HE4fRdj17oLjyFwR3JvFtOSkUdr3/7HRqsAzNW
z8losuYU1DJ6y/LG1Sktdhj2rKx7FLTKQO0ERhWMPRsW2gyJ+1X+8zHF1Ce1kcooO/cWf39C5nR+
TePraE6dcMq/ntDA+dBjDh7jO0Nlh6Fh4Im5AdWkJ6pPbPyy8/Bi07yGXiHX6Py0P1AildSOAqiW
y06o0Uw0Igf3w600b0ZFdcIL2h+gJTh3JsTk4l+i4ScaAOAoGBDfldyR26BJES4k8IMaDXVUWt8O
W7PcR4+pXLuN0x/6EkUhsJUfhCdKe/f2Tp96qqSUR9BP2H6Gz75IzaFLczrzR7vJZ+lR7N4Jo74O
qTNmvMbqBQ2DXJIGILOIdFljaGRUto0VGGeEawK47lqsMkIY6+sHB9+Gizj12XX5AgvDVoeGVl0Z
njbQLhl5amqZVsftbf6FpKUxUbgyS+v5UR3D8rKfmLRr7H5p0witLWCAJmxNjeXFQf3j6FrTZhhN
cgDArpVsxKZjSxqJbWopTD4JBlcSn+YpP0ha+n5G07WXVR7m156zWJAvXA7keQGb6koyfw/nxCwZ
VrPzBBmA1zlIwfXpockZRa6vFSMb9jnnwLjqa0fowuGoxZll+FXGatkG7Ruo0WwBROnDh39u1QFp
m1y0uTRNpAmq743kKZ+akR+0L7SyT9ZPNrYsQm1RRk8EA5eqWjOTSomxtdEHgbVlSIB0ap9ZzVOY
f2iT1ehgrGK0jhS5I+MFtOQR1mt5iFhmCA+CZHchDL1BNK7I8+SWQxwhLcWcsL4MR1b/72vWrJfX
PqlBwLvK13NakRg2c9NcKwDEGi6BJQzkDwLPza4qoq1T06c8wP31mo3XnaezuPjpr8Y0VDmAIheC
ts7AOx5+ydlhGmr4gOPsG/MksUQPzr6IMW6y6af32SBJtE4fWOXE7UoGyWuB0hcYTYdaBn7ZgB+a
uobu1nshyqhs8Kg2Lg8jByLNJn6FzEE/2vItP0CyVrEMru3jbzxQO2iDQaNS/xBrgR6hR0NKKNll
d7fGIILCkfS+ETAzisIauBPd1g7DJ+BZqKKHEsNtqJ4m7PNii1i55zquheRU/yLwdJ/pD79Ctx3j
kWsmF8UYuV6vAJQDe3kZ2OJJrM3vEcanv7QToCuNm+EAWLEg6dpAHhAZIGbPRyZWyjP0Rqsa5eB5
F1nVuWnTlyWdr3pQ8V+cfsxLqyPisd18054a3vFkNMAlyUaZEHi05Ajq5D31xKFNsv5pjE2L0QT/
mtchcYBxPOkLFJxIw40tq5G9oZs9paHLJgdbOdILc/sMmiEyDEMLuSzUWOpi1hBkKJn18SHQf2um
zN4r7xwJ0jlm/vxXh+Yjxq48UrjV4IWaLkOyIhfPRoaRgM8718cHO62xs4VwQKgLyEt3haeqBPts
uOEj1hk9qla48o3Fki0Y1fu+Ei6191nlDq3U8XBtMAz49tgePCxhnbe1j+qTltSuJ+3BNPAHo0Fy
8yxvNEhSaNUfOOz7ki5UzA48YsGRxOPp5aUvJkJxVvDububFaIpgvRDxMep8Q9qiJVAUyRKCfuOR
fuKDh0p7lu2pyqErXtbE7qk41859tZhgBq422Xtm3FQUZIlYeOkYgYcwpM80RA6JTGBowr/cjuCj
UwSXU5sgQZvVkCT/kqZXpRba45typI8H4572lr+LuVvqNkZBvDXxcSCFzQl8WA9LMLyjCMX6mxYx
ljGspgJ6WRIF4jx+fa3XfP8GuIDzF2HwE0B/L+EAAZ920XDpkfAzC5vDhgBar6FM9MlSWTqjYSUU
ZY6gfXpMe9IVmyINZrZxN+jzeR2zsAQ1b56SrkBWP0eW+w0oyCUOWSck7Dlfu+l7U8bLHbEwKszN
HBPBrL6zJ3mEiHgyEWR4Y8kCxoPbtfgrOKGxBZmYkpy3rzddsmn/aDFMxjlPwtJQNo2avRHakCxP
FZA4dqbffqQWwZo6rUChNrAFUntDi5AmIY92KnLrXJfMpYN5C8eqs6xDSP/1p0whWFJAEtlYzldY
tJul1rT7yNdEJGxmW8Lla/IGcLH2tjW1hAlczBNEN/s1KWKKK6A4Qm+NUPzFxAOZr/LfFSH57ff/
13Lmrcjb0IlVu7toAUpU0ux8vuxfoWazoLVjgj7odEgaI1ofcx+XXg0Mizrmx50+hRiI/PL/lJ1g
ONEgER3ZI1aqFssn6w4kThm9Y2I2C807wA/wpATRZjUp1pttUSXLi4UMAOm3XLuc1b0xluxq7iz2
EO40YZWlUwHdxXFGrH820Gc6Lp7f4/ZCEDrRsj14RJD0vQXPuwLHHYY08QHN/1E+gfzmUXbBK4nn
/t2MySfsAhznLCL70xeS3q3m+6v9odR4uAgNoub+d0UcVYMFCEnnX5jIhqDbmt4g17FqmV19oImS
uvA7DqP9STbnO5vYyuIzGl7ECB6odmTwDk0p8LXPYH1Ljl0ZOSmor8IQlhDe+AmF/AatnTnqY1WM
bOzfm+q3WHofpPw+G1L89ue5eVIz5LyYBFSVuLu8ZgiY7sIm2Dvnyl+BdnLM1ZX6dCHYOzm/afhr
1Wl75SkomAt2Kzk85AZGAW4xgODQdUELiK8i+/2Jge3VSKbxmzET3erl48PzUJUGYGBJHvKuNzWA
kHxg1aCbCrroRqkYFzinPvRmw1vWF+9Mhd0fQJHXrrplid2kII6pNQFGh0QcfjkHet5bsRJxBp8q
rLQf/WZniwGDG1voPIbd/EGoa28Wyza8x4XFMy4UxsTZDkk3Shb15/GY+dWtrC4QRQNFSQiiTyPi
xOF/h1z6EgQIbsDkuqQh+qqMokwZAjs+ALXC6C8uoZl9LiUXx8IMGff71LAMmDNuH186RYDHVE2l
DWwrYdq6uVtaDpZFzN8+dXtq0B+4H9RVuzuL7CFrVtfybTSS2erLvIJvvV1akFdJtM4V8lYDdgNQ
FfHq0K+BmYO7wEStNYL1iNMw3Q3bbSgL9+WsKN8Ya1vvGHXCnQfTcKntoI9dtclz2C5OZCEqScCr
boh2eKPvyiTGl+TDFz4FypG1/3gyIPZ3ZjbCZ+YnJPEptK6WPn8SqmC6fzJf/kFvqNXSntntrVbI
vWZIgspbg7hn7j6gEwbQKc0An8yi/+b0BKPkwJJtCSD4YNk15yifcd4B0rLGMO1sYuqYkqrSN74q
w3BfpRor7rfRZUbnB6IrzMGHkioQoGdkmUBj1myxYU+cxxMRfIdrLcypjx9B9y9M2NjfpVVrRSmw
VlItg6ejfcjmxUzQi0NBPfS/PyX7LKCzTAGZRzzfdp2b5b3sTL0vsVM6Fw1T/7twZv7kr4/DmcgH
2fVQgdFn9EU3KVhBOqMDC96yzr6qbE5Qg5jqKuYnzb+fAU9DyKRBIZQHJJvjX7VOdgnJBrR1flwC
xNRQ5RtIu+sLat54zrC/CrTLL0TdBx4EHTRyEpW6BOrKfcx9Lcb1iiAfIBMDi9AqZwZqEw0p+6mB
AifKk4QBMGufEcVIRk+b4naJ5S6cuCInPbCtSHVkfMLofajazyFhRT3NjmESISNw3f+o5EERBDL9
XbJiSp/CTXijq8tjlhg7NaPm6yPnEqPYEwEinFwbJct9doZB4ORGbeWeEk8SRtXeENPEt6tjFd0v
Q5h9w8S1fnUxJhiUzVaHva62rPwiRyC5f7qnHtJ58hZzo/x4ayUGyVbxYLnPxPfdtIJz+M5XC9w+
62/Lgju3KbpfBHhflYzGB/CWQyDly9i9RM/2QDNx0kiXsc7QIaABU5oEO9rjaPT55zJMKQmLr2pC
R9gBfMbEC1ESFfb1fcLL0IMcnINj49EN1Im78LGG16atIfv5DFPe0xlvqAraByq+x2LB4SeuVOZC
VNjHfQOcl4mt2pV3tOc2NltT2Mhhb1gzvSQWKC5heSej4kE7QGcHxC95Nt2KKH9dYQRNEU7WJJ3G
EMs75hc6vTuNyV1YLnULBo4CoCe3HRPZYUl98HY5SdAtKFLWxF2KRmLwX0wcEOk4rUjzxfG4y9A0
SjYyVUJmEoTfCctSfQI0M4U52GtRmcUhXtWkMK1NjZoWEUw1yvOWf4CGI4bTt/zVWaCM/39bE7SL
vRQkpUuFF3xcROmTfqmDKZCkLY1xj7guBPFsZkY32cl2BiniO0JHTfrGfBIrHlKVP6fKpLAgxYxI
5mu+z8Z50A+UVXZtt5ghyT9lXwo7bU5aDefsqGAQbDMwXZWuKKZvrgqBiO20lqoobnOyT0fl5ZMz
AaddsPPdqpS28PFpsB7zoqZnZbJPt8ditttwtjnMSf3DRyfxnUu0LYayqlZ6oSdga1JfhywKF5l3
qvelXlue5Ls/a25U0Hz4JDzMOhWuu/zDSsrrL0kZrS7TVVTdezKVpcYlAl9FZ1a8cNr/lfBOjRu3
7HMtSFzY0Gust4J3rNiyD+D1ytqlYNIOP/zLsTrDhbICHUFVTfsRHYZaMMc6AHiv9FqKJx7xsotb
kRcsZ+7SZsktbXHao8alq65BdMsXcpPeA9QGL51IVm+ZsKfCpavTUTsyQajQeiDjHxSkqrB326eg
H4BFhgDtJ/Wxe06a0AlpEdQFbsWc3DrCE+RLrcnENQNBqwxqV759Ujpxi4TNKEExga/aetJ6TSzs
rwQVwPpat1wYWzI4MWVHODlNh/MOtxSbNhmpJ7UyrErkkg1USefk+B94BA19wA79PWe8lmq9BEj+
31ByZXTLOsRv3c/QSgF5QRB1x3XfGswgm20IQHN0JfaS2x0E028LbEHDvL/XQEF8tQQNBZ7N8V8j
qkIdcF/yybMISMU9oshRbr5D1pF/pum7V6352w0RCrCwx0UMUag/MEzDenG0Y7U469+xywXnPams
snuuk58mlnOegT88fwue5qWVkPyhV38xILhERqttSXs91WzbRSTrqjoHMPVsxyCyHNJvRpufQVjt
x8/uu5WDy5s22/0ie1VKupjjVJfaCj541OAAN8OocEz9clxvTVPgj2q/37RBFmH3k8634C7XNyH3
5D7HLpaJoKp02prBnarTX75Zk4Kw581CvAek3R3NXXma5oev64ag2B6aEXWlKJ6/9+irpXNyNIWm
pSIVnPGRh6DE97AWVkCcqdHF93RbQpSiJjBlbYIuUAnu8e0nHSXGqdD1gMb3Rz679CVACmaqZfqc
11mpGvWky3jy8Od/E5DBvk4eaWgxSeZYmq1ZIn7FrSiVH0b+M4YwePrSgwyFvCN372spfDKZojaS
E0y4WoH61OdlDhl0Rwf+9AJ8TvyZGPwf4TDpMOSDOU39nmkdg2TbYnyk/UgZJxqecZp1grDKSW4S
f2AY7vYFx4AQQQPduj+QCzXUcAS6iF0qYngsshXnQFpXk9GJbQiYg4CcLd/r9Tz4I+qgdrnM4y06
mYB8I8Ito/K1nyJJHSZtCeVfSg/Vt4zc5gAP5N5NxvJ2zBvjmfDh2+zNHACsnFWREi8JGGEBo2d5
LfV36kvfSNxH/xCPOmiF2Dv/JCdxzGcMoBd7cue63FLq/vAERKO0lUdNexrvdagxb/eIH65YDh/o
g6O33ctQGqPcVW54ezunLLNEegOLF6SFshTMIAEpH2PHZWCRKcWVgYdluqUygk82AsGZHJii+g99
rNDMTQyzQhmnMUWn+0YIFneVNFZHXdWcNEWnb7yTvBgdti9D4f8DbhKbLmCiccP+AJitYVrDn6cz
KBZD3BwvIOZEg+zAZuVrbsq4nCuAw7iikXZmgVPQYJKtw2jgfQQ6Dzx7J8//nnYMze5bGQ17ZXXF
8PPYWLg51mR5qwu+4hSLgjeuy0kpgmV5aVFk066KoyNItjO9gViJrBUXeC1J7nzGmTz4ip0wTswc
ondPQOFNFhBaFmKouainlCV1CyukPmEm/Bkbp63DiigrEYMLHq5WevoKDr5XG4Ah87bxzmPHSqQE
/Dy01tVWOGfC2+3eVOjAqOd7yLp8v8Pfl6MVIhkDTXHQLhOn3wjfelHuqSVbQlo7Pn8olkoZb/nd
+CXvp1DukKFpoPjzTLRJf4qRcsPtGD7E7M/Jx2K/0y6obA1hemofvdw1s9VL6IJT94NAnk7/KcbD
jcp5rpPEt0JRTHXK2yVf3E1WQqTOidDfWPiimRMcVedQAONH0OZWVDqVkvVi85pFmVIqBNmHaHw/
jIvWJS0rX90MNgWhcXeCx/k2aLwwd66n3e99yfNbhtS6dARWJpCtZJtnnAi0hS17HGEzPxSYAOw5
2Bx10IDmRB5AuW778TdsiWmAjsm1rGjHvN4qoKtF7MiN16dgqBh6Uav7BmxhCmoJXxjWsAPh5MwR
GmjSgxHJzivbJPLzwJFSI6T30Q+aVwjTOgxvjBCwjWu6SFmY8WL+fopyomKQDVEm4aKRxfX1JGPP
71HiSxlGF3ioRnZvOc4gPe3Ne3zEnfJTj0Z+0qWrPVxlI0Imj75N6htGMtBe2lrvUDcChoCZWCjR
D+ld6TjcRZEOV7AKou1dFbnv5NPa3JkxbE58es1ERbjDijzPbWAK52uyJo54oJxU6pUQ0qi2TASb
jo6NbLSj3diM2NvDK25qh8sLa6vT/f4MQYnnhdMOa2549T5kUF4/88Lj4f/V8Vn2F06408aZUlxa
ATe6AYtVM7kLsI88KijhQP28kIzdAcNfIY+SUuLf2ckm4lXnfncLXZSvbInMTtKEd7r4mfqwF4tr
U3ULxPVbj3UJPFsuD8+xtU5pFJ2qI00ljUoO4wJ3nYv9WXwscdD0Fc6wncQnEisOmxXYUTjw4Wb1
ZlHdJz5xAQuuIsUX5RVo0Gp09hZfJoycCsBScYKuJppqEluiHJa6Ed+vec6GLNDg8tsP6HwVOXYy
ExAxuSK51LoLLjjGZtHSz2jgtoijKfzJOm+4tGqmjg5RqWon9Xom8YR6t1ItTFmuFXTe2YcDzO4+
38bS5TV9mEy39ByDDaeseCvnR1eU2wDTEms+t84Mna3ewewTEiLBDRfbtEIXdoATszXkYrh8YEBb
0gOoTo+Iqjvze+QSq86fvwrgMZRdxK7pVnbdRpMCVViIdn6YIuiIBhO4wzlNvdo+2EGPgZVwTlEt
ukwTOoZcLYMkQ1tzf9RON2L5ShSqUDFjtxasuFFUYm7sHyv5H8QIwDzVgnqA0nGTIhZKsjFcZreH
2ID0Q3FBTg9NqMoZXJyKy10XyfUOI3U7+uWhsVxkAfHqvqrT9EfjBvetQkV2o1ecVTb4hn5hskRC
vUN8t8bud2si75J5TwPm0GWacRdDPeFM0j7eq70tEl2reTXVP3ApCXPg7foVd65MKGT6MVbbsPGH
zF35ef6JUJMemLrVAolgeWVlSBfZC9gNLcx6SSaDB9QdoeeNSCVzsQXEEQQi2X2qWei8BC2JnlRP
RmP1Lii4NZefvOKvY8DNWen0OdTVVYb990Vnuy1979R4AWdJQIREX8+ufF9PiwLIQJhQl+8UZsTy
T69Ka2eB0rJJw2igziP2GQFSuTNnfCU5eFyihutKDTIcmPfXayiu8SQdESLzB3Mom4vdIFs8JS5d
u9Cu5Zo0tMH+0P/CKdN1l0od2Pd5wJTv0Fbdkbf4d88RPr6Q8DkxluOMuSfDal7CdTZApdcxSbZF
KlUJmWD7fcUI0h9rv9VnTzhXRKX5lQHN2fiQc00Dw99wCuhs63RLmZnlJqGdGAfftIZezXwFicyb
NPaMg4l37qeKH15KT6UvLLkxrWyygmWCbg2/kpTu0nqECWwtwl6IccXm1v4SunKw3cTx6tnWGvdZ
wo4Fzbxs1kufBOKdOnY3BUmtOSA/TByFdDz6GEcDbKsMKvkSmTnxtDvm2yMT+hS34b307Mv8Mxke
kp1DnKRJ30UNfKjkHXGyLfuBKaDgI5zd/vSUErd+fAZwI6riCHFQkUxKsN0E2AobVDpuuxApWcbH
Ta8ao8ey8GeNp2UWFZeD/PcrQfcAnd38ek3Sb0k2QMI97Q3h/AYweE9/+Nc78rsx4zL7+uJTkD59
89OcsA+20AH4VWQHPm2yQqfam2kwdzJvG/4rFWQBs7QILKFwmCeSZMOfXxJx38WD9WYzVWr+KK/S
RE1ylTFdY5+RHdd1Kj0oFPjCG3rK13YalnO1PpkJTTCH5AGFpW+LCizsDAeEhrIZNa9gRhCdH5s0
hm5zXGtuUYd9S71QzyYsh2jTHQEsmLZcNP7i0nPWWoHhhocAWjlsqhkuoDwyczEIJrMnIFBejFEk
rC3fU3ATiHGMbboA61n35Pm//XJlyz0CdaB02T+5y+iZUSPnCH6PNGqFJeLM83U+eGvIOP6kSFlh
huRVEi3sZp62eFlqQ0G9GTudqemXJqhBHr2N6vBpjl7K1VDPe5iHQ4sEUGgxbgisXpaRPF9zL8Gp
iYSaRdcUS6jRAij9N/7JxhvwJm5smaJ72xA3teWqCkELKNKq20DQNSvJ3P5f4I4g6Z72jvI0sREq
aP+R08iYK7GIwvIZBFcXLtoAJwJmGyZfc37NThldYpRFdmDPqh/1ozCfB6dLmEG3GQI15+GWqgk/
XbdJa6HX3lqNCkukPVmL7bbVLru1ZjoEqawDDoMrKpy9DOTxpI3LbD2FOekdeRocQggDDp0+56lk
cN+WeM3fb0Z+KKzngawY95cJAo82qg2J9LLmP2Yo2sd7TSEL2UfeoBaf0GN71t6ucB9CgMuWuGoF
95935ojF9Ih6tKhtJtogIRGtCkk7xvQTxKroXH3ZYN3iB68x73QIPHgQSVTbCaR/on4NcQObvzW2
TWXmepuk39RQuSY6n5U8Ni7M/HmcS4S89HrMdN9oSzBvLYn5EPqJUzNaGSD3OXU8SKC58VRHf0Y8
QVH6MxbXXkobX++iJzg6L2TbjzyMEtjnK7tG4EEN071OsJ8Vnu+tO1PokjZ5eT09Vje2+5WVLi+i
b9bknxckb+jV+q7qz3BF5WHNI6G3QCsbMrkFZ1fyUSYigr3ULouhLAsNXSYvvGtGM1Ihmzsog5ou
CW7U8HWFuzjqOAD7/hN+ED8TqYjgp+nZMrPqawrRljyAm+L/P9SU94PDhvbm3uyXa4mRRKMq3iNK
Hbcjwmx1HLUvpVDrxiISgHtB0jsAQUOyxcT/JXwfZF7/6xXw7GdlQwbvIb67JqK0/bzlg1Hc3K64
qscsxDKC+H8pmp26wP4sy6SxrImbNULVo2uWU9FVLTi6sBV0wxmBn1DewzoOIqCTZ9iRjSMAMefm
zQ7HHGQxnvT6znCVPG7CNIOSrCbypRo2JLpj3Q11KbvWmhEJ7CKyIsHnRLF27gTpCe6rOSCZtofP
+1v5FFq4Fiau2PVjuAcboiA8eoJlhBK20MCay25iuK+0jA6E7MK4lrQCZiq1JQFJXgnvG9GZjocr
lxj5IIRWSENKNUjfodi7AR1X207bEU18frE/+aItsPZCw97DhyVsGdZJT82tb/Nyxu3prEl0XjkU
Xx66alX539I0k9gXbtHpfYYakJd0wugIV2hz3UfinD4lL2wzf5YJaxiIOgKfUCOlQt1mJU0mA9ZM
k8juX8PphHECuQUUL8fAQisWk+/PJ+yufPfpAWbxZmIeAsVRTyUpPBhPU+QwDeZVlpFANMcnF5US
MYPCx5FiOFV633ZqXj8plN4SO0887GCJaNlT0kKGC17JSe3fw9jkrAxLq4lx5WCBwZSHxhDulhSp
WuqwVYQkN96kpUb+MtlF4DRTXpFasScnpxRs5f3tdGxHne4RSB7yB6ix18xWlJPx7NuL8xc96WVO
DnQZ2BOEuZRhhr8zB0U0cWkQlovCpxKgw0HHqFWtHTJqMEmvja1ui1LPlQkoQ/tzWMh7v2Pz20Q8
rfqFkE1bEE3widTrytBfhWbs1hxmPFKD5MlUSvzGMTnZS78+9Bw49AbI7K52o6xmxxdHmvU8dckA
p3iieAWQJ63ioDGGHpRzaZgwnHdaSiTt8153oQeIBmzgPWrB3wsKE3SaqcwUmuGiTnFSGtucZKRL
TwdVKpeI89NjfTdiAvRcZBCD5PiTkBaDFlCIjXsqgoDl4QRJ9txtArTSAm3KC3gu0mUFYShXw39/
AWiwGza8whuIcg20s3lfS2hDn5/mP/RabpZ94mKjf4+ZXGLVOrXawsAPaSXfE5G0YfKqcKack/fh
0XkPrfVAfWu7JWU1SXwY6F30Vah+PmMtgOGOPWH2Hlq4IWgVt8krNmDc7Al67WsDuuZsFoxgl2jh
YXrL23k8Op7EPMU6MggrTIM4N06lC44X1GTlV3Wq9gyHstlLbXp1yQGHAPcV0DNt4KUNvCxbiSXe
YWzyogJgPYceqFDdvaiyHr6fo5GrFgW39qkqz90Dcv3nln0T6/eXPFFBjcdnCRhtMksc4A1zq8Aw
a5mwCwehtWy0UQtJkk1rFOHkjvvjwuOOWhMv88pVahH9cVL9TRjm9QoSCN3Akf0Nph4jXxw4PLTq
XgXwHVwAQHJHTH0bB5KqD8+GC+Rw1UsMzlr+MfNxV53zJ/J0YZP2F+uDp63GN/z8yVyqGpLAgCy5
Yc280KTIPHcrzxMECx01YV15zSu9V6iFY0sCQ2bb9FENG+ALsKOTCijPM1+aX2tXO/T8KIxVbcWW
VU2hs4ECE6P+hfHnLFv8KG0Mf4wrpl0WBdsxW+HU2Wh6dRwP9VysXfnKmDJA8oAelfdvyZ02m8QL
SLP8jz/oXPRQpN6GobMEb6SmYxWx+P2P6j0zd+gJEC9bYyOxO77VE2cE5R3KoZNgUJGJOOZPhFFy
459uNuMznIXQ39V+h77KNR8BMUS6jLIKU3AJcq8xRtAH7jauDrHCVP1f1J0VOVREp+Qhv8Vob5/1
6DU8SrDzu8nAqXgO0XkwIgLTt46feS/xrEOsdl6CZD7CfCG6+507bOT4dqnsZYrDWbud5aRHIOF+
cbOAqvqZldeAhGO8eZFtzr2RtSm0iIhTiD0jRMwTG0MgbRbAd24atnjxEl9Bl9EA5116PMA7mXif
s8n+ozs8u9UZ2kpILOFoh+XFddtLIeCnHPHAYxvZc8GMyztxaXTChI6eeatHm7trAS/3MosBKLrf
aZhNSC7vv+Re1WQnoxeRjbKpj6yfOTDiryyeIcrUUB2QzsVtJCCnEXjsodcgTEXC+oNzY0rCuzYT
gd8WmQuTTJarwJ/iFhWW3vIQfZz0/71arktt6Q92I34tiXDAg2YtrC3ZXqE2SCPjlIJwPEoTF4r6
t6FO3oXpAUC69ows3PG7Px9WegwikQt5zUX8VtAf9iSInJ2kIUvEXSUf/BhNKlgpEXeFU+gtb7nl
dOVBBBD041ZjGXpIKIIxjl0NEm5jysS2aSEkX6R1tDxXLSrZgPwpYYS4bYMqfzu3lCp4B4WGWHzE
yedFXSdnta1t/XONuf8c1GzBpTQIx5la2p5P2crFl5mrMQXb/KRRPk6WyGrRiFL9WoNd7OYk43pX
TNZiaYj8S7aXmXqkdhP6d7VWqeLtOBHtHrxFPx2gEr9QBZz0Y/3Uy3dbnxMooCKRIFWbsISPyItr
dzxpk3pjF4lpdHA/wf+DwaGLkBa0S1dp+BvJhUodO9l03lpaaVoawXPVcmkTQZXjFbkcA3tNJR6f
T71t9J88ie5VktUT27x5LoZ1a3VC0PH4RmmPfHAkg/+Spq4gS1mPwhI2QLtwLA+1Pox0EySOeqW9
b6EOtnh9f6z0hM9dbaKCl9JSWyNXb5VpJh+dBvYT0CIVPHefH4c3DBlRNuJgxctysSOTXcXDxzVD
plPIvY4o+UggXxvOgmqL78+auIuDcrFoIbC3svPkPsTjS3Gh/gzOzU9AU9swf+Sl0UL7zuCBDBme
hEY0BsNtRO1B8XD6owuq7M25RNmGyPHfW0Z0W8Mc3XaYnUw2YfJ7DxCFauXjYhLFNiZidJCFhFRM
tliq46tDtGp0RXVM2LVGgpXB9JIL1peV8MkLpMLBqSBNNmjsidb15MWEQlaf8WFX037q2rLlG4W1
IVqOlDIz3bNXcH9GZYLdo5dX/rz30ts8hv3t/gBEpGWjCamwNDqyseWMCyc23d4Y7P7RlGDmLVM6
+QtaqAVeIhaevZZEyfAUKS7y5x5727OgshVi885Sb2G7HzTquqa9GIUOFMSXPrdbcfgpNlit2wsE
gVMvejs3ASYtA+ufijQRA+lJvKNoqs2MPgM2DDxrheT/DuHrD7J+vmmF9RvCDokDRXremAU155Um
iwFr76yg5PTDsd1ZQn3nMLPr7IRyLkb/fkz2w1gnamt6VOM/nRKbM+Fpp/DKznhTNpEVzt07OZq7
GYBftqEMRVdUwQgfxwEL9/s8NU7VjuqzVhevEVWN3VGiw6CKUDtiJhy9OgjOarSbWzDdmeuZ0+am
ZPNq6LXEQUsnsEWmyft8/j/RucVAI+phZO0cnqpW+oJiU5t2Lp9LApxqFemalR3Lpq0QDyykliuI
pDBhxdpJHd4SfGy9neufyWPwtgKY5d+K8U422E9COaINHZOZRm5T8+R96YDB2KWqmQFu5tiO95Bo
jCdukBQI8MSFHgf37gizj4ctOHUZ7S/Y/d0jmtFCsx0+rv6wkSifVsLc19JqAza94rqPbZAccvU+
IEYcMDXSc9DzhESwfP3RjlwLsV/CnGa2pxtSPuFsTuEQ+61jaTt7hC2jspngs81DMnlzfHWdPJPx
037/4fjgVvlTnghbIgCkincPFnLCATlEunP0Liv7b8ido/jZuZ9++wTgAuhaUAkLInRc5tH2Wrpw
YOn/0+a+1XxB9gnoustw7FtaVu+3XYmaSup+Z/B7N7WfjE8g0tZBHCpH9kuDIf3eI8Aw7pQS3MS2
s2LHRqf25o6Y9hvmKb909dEnhXs5pchUbDPg0wqvCHTLs8VrQLsOk4ZH6yaxCKmcwGIYCqgx7Jn1
GzJ2AX+P1UOK8Ts4t0VyUi7qkf3YMvCc9OyYrTxJoQMU/YfJ0dWD6CmVnUQOI3T87ogdV3AIVOzK
QUd057idz6X+7Nzzuqf4U48waQkMsnm9/TaOgQBoLGQ7S0SvdEAB5BINEEU06KuZgHngwcZFowRx
NghBwNzGhnVnySeu66VaMMN8qdVUTHKh3jOT4SwpuX9uE86v0x2AHb4GNj9tktrZkZqDXStPDJps
FE/0gqe86SLIdWYYos0wN4YdT8nOCpU/kmIrmFnojNriKOMYRrm0e++8k9VJqkqJBIWBkV3OVK9w
UlR7EnM63iNhbUynlYtdBMODCeaJEUYrhbD9wj4qa9bgGK2AKGd08hXC/pkd+5wKjS1jmBAtUc+P
q6Jc6p5fqM+W4GgMFpJKTW82+GHB1Sfv3A7vqs0Dbw5J8/F8/6nvEWKrTW1nOZlMZeQkTAI+kAoZ
oyUcsIk6iHJVx4LY6ad/u4ioAdw4WWgXF0d8KCtFBUeVqAYBlTgj6atbfIZYMHQsRBrNWPtObPn7
8Pbz5KiF5EfnkFrZsju6fm4S1WwP+AjCsEBrOJjSZX+g/XP2YiXbGwh0L0DV43dUxUZx2Q8+ZcLW
WI5tWnEsu7+48fakyDLzshvuszwn0un6o9hQLUwlOhXXkyVJEFe98msPUwzJuS/y01MpQXBwVLE3
qmdrR80vqO6I9YUd3pkEdmOiIU7mrfmCR3bSYJTe81P7bjmP+WeEymXpg5TwC9e26GAyXMj+yXNu
0OTQE6riIXpAiPKnXpuG0onh02R/4h8L2YctpsSLhyQu2qgXgxpqH3pfyRjFAcQBr5N8PpjgfMOQ
LyGNEwkHPlmokv6yWbH647FUO3Pgzk8r/u0PvGY/IMrbwI+zjg5SId8Daa/T1XrHzUEzT3NQS8ph
cGz/S0aTosQ3g5wSlYnvFK+yaiw7QwLKq9eyDHNLNbwRGbKM+pWqEa5f/bAqKuUnH+IndwiNjmKl
wx0QcTq6D/Ta8G5OBy2SPl6PUhR/vu3qlRMQo6BtsSOVSce2XJVg9ci++KymiIoh3RAom8AfPAka
T3NPGyyKKFUd9rvPmNkh1tFwNyBjh4RZddDd0bMfBCjRcWDPzxjhbwpM7mq4k7fDlLFX70xCr7q5
ye27nWNikD/z1SMmJ4TwvmFFnrTXqffmh31EVFcEi1psh1i/5UpirdH4hBzpF9IWcqrXstOh80Sf
z0e+3EHrHLZMSCnwGhOl1Yak4tq3ai+I1vEpe9IZ0EZeyUri3MkOOUnA6QxRiQnjwSTjgXRub1/C
RuTxf4p1+nptirF97T5fjyM6M+ivDdSz92hjLKL4tZjhzkG5DlFrlPHK/W5VvJPj4RRl1MuV4BfQ
FvDigmBzmJON1mQAM4aZwvlH+y99cF3TxZS243c2JImgdlstjBYLArpcL1sm4ngUl577lIdRXDEr
WPTsEYi0A802W3OsFadY6zrjVe3ge0Op9czs+b8ErOzYOZaHsIarmhD4/b5c1t/tJ0NDupGt4l6o
ZhCshK4koch+A1Tzt0B7iD0H2rG56LqKsCXPG23TZ3ZvyMhB9YVL/k2hBN85c2tKWGcL0WvBs/gn
IBisDNv6PqYra8MHEOIil4rHl8J6Hr0qFsLCVb+8GZsTFw+BH6mjBG6nzhp9bpNkb6BP67uEF85K
4iDePM91AejttNKFsX4x+fKYYRTZ8hMT0U3Idp2FrGrfirfmomm2Hlp91CMA6kaA/Gn6XCDInCwg
6A7s8+kjbGSYmW3LaIyw/eszD9gK5h2akPBAy9ASzmkVk0nuQVCse0NvcGu1R1FVg4oltXM5MxO3
L1EkmDKA8JgqCotgFurvCGxlArrz3ZmOHaGPEMfvyGY+qi8HI6LwurJXWaXOjGSR2xi5awzw6kTV
OjXbntZxL+PpILlT8bbJp9XAPrc49Hg19R6B81C1PMzahVX+W/FrtN4hCBELtCCqRAeco5+ggWqr
xwawYVaiWAfUCJrfph/faZdXrbJwfhmd0b8bnI3R6xn1cKvzPeKKLhKJbI/ObA5yskWSf9tYr3rT
LX0eBKoyvgWVMDljWX5kzvQmLkdc3tJPa1guTwfOBe6zFqoQIqzhVMUmZYGmbj/tZPMXIhub5G4s
zGVh3tcHqrXbcr0uukVKnrapLA9hBnlDt7a3IJIeBHo1+ecRQ1Fa4vfFN1RUXtMrziQffYkC52yO
xMGcMMNIYn1k45KSnlHx++6LMPwPxgx45QZeSAhuceXnDBQBEoIZ3JMNQp8lQ3ReWfRvJdaT/rTW
4CHjZQmvGQUzRNoUQRraK6FqPmoZ6pqxdjEiYcqyFC1Fu7gKXHrKWMhI4QcxKr+u31MiFuUCuvof
53mgFkLt4CuxSSQ17Y5m/zJFLsZEH/1CP0fzgF2kunGzaCLc/Ud/uPSdZE5eJL4B0v1TpiTwyPCl
PWrnKfG+1gGqSNnDWd/Ur1KgqF4DswmQNUyaW7Prc+2Xb8GEOkjllgebpzkpipYJQSZo469lj+Mx
0XzxdsOPDKfaBWowx/Nro4eSYSo1HMPrsav9DAZ52L3p5RKMDz5MAFDu2ee4q9/RucHGGp/K5UwH
ooWrALqx2npcyhrNJi9llr0Cd1AbrZ3nQfOzGLYefrl7e0aMyrHeR53BahqXJfN04ad3a4CZvHI0
Yxk8+db8HhoExAtqqdBW57UOinaQBnGPD+WbrmLY2nRbDa+gSp7guIhwiBFrWZeLaLbAdmWXk1lC
RiR/BkO2jktZ4NxIgypWsJ/vvFmCCYohkH4VJBWywGXolrkutL/yB4DAInCakI+ylejT/5QNTKP/
uruwSuPXwfzZMI7y3Vni1Th9AdTf0P++3zFaO8dgGFAprOHDIT0IHGym+m0QtGNJByxjH82pDfF2
GmbAhrgC86yIjkKFPa6k7tojdCHm7B+vQAPsRksp1XVCaTgtkabNDZjHk2e8IkGT8HJp7l4J4Vtb
I/yfgVMxnn833YfKTdaiRYjkH4FUFUp7v7UkW/WZ30IM5xL6oz9CfhrXJnjIkWHjmYle5Db/XZOs
kzV1gKE4+LRlOGVcpEduT4NFm57OBssCvulZLvuWtEAkrp4IKjIuS6BZIXge5SHNc/ks8fOkEpOh
xzuNmEwws6PUvMsoGJ2I9+VR57qTEmuis06gDM5BFiSBNYGHiPQnay9qFASxNN+XasCc1CbwEoOX
u4xN4AKZPp/vlGWskXFvfuxR1VDlbJEO8qCd3x57FHGmJ92ejSHp78KL8SPDdiFqp61Yfe33fxPS
g4G9yMNzwRALtIbFwGZ9yhrfZTTwyx1u4k0xQN23tWYqk750Qo3woaPxePw/fqVz0VgYb0EEow7F
SsZPPyMcad/UVhHsQuuiDmVu218smcJkc5W13EcQdkswzSu+oruunVAVwIKuBXunujoDSlVtS106
IVqdVMOgnCs3lVR7Ku79v/Hh+sPU3QmqHO4JrnFS1N3Pl1O06SiLGajbakDztFMAhXldPFTFxrvh
hPvU9vsSrlk+NhRgDAdunozaHbvx/NplbPjG1WlZUlsyj3qm86tFz9uQm5g6NqqPOExekRUr/rL+
CzfHG2ACh9yaMPScpj4a6X4ljTesvu8P19tmNLhX1GK7mAQ/lBPcqL8YpZXy+ZyWOS0Xu7Y1JGhe
l1El/GMT8/nNpZjoNMAFN7ToXnVf5kbMxXkdK8PECdRs/9XcdRMxTf2yrZ1cTvYJzl2d0/nzylNh
5wzlcE+1whejh2Qv2LRA7Gvdajv2ejnLks4iNGY+2vOqqTQ5b9WfHPeN1bSIOM8mzwXybmkhFZAw
xKzzw3NdR75vZXfVyP49GzyZzHkoLvC9YC4MysasoMcr1f30Oi3Mzj5mNKoGG5w3VyN49XPDK9Xt
6qke9SKBUQ1UhRGqU9GmL9ATUHS9Bt/ICgbURJttmzFvjnxo+E5wNUZ8yWDDiMaZ1v2qbsXnK9zx
JtS9tmQgstNoI3yIf9rKA7kRsxpUWH1pOZksSOQyq0r/kooZmKhjePYrDKjF0sU+kXsBMllYHB5u
/24b6b2MjU8Gomx9wgCgRn89n0dMELeN0ZMZsIp/0+iHLfXa+ehsIFtDbnFl6Jkz1T7f7NhIvcny
rnFmp48fvE9Jo25j/vB6/zJo8Bm3j9cXBzLf1a+/r9xz7xKow0waSyXZSi2HM9yImmjEAUaLPE99
2VQLsXmvKLW1MJLTBQ8tr2w8g0S4do/Fxn+KXI9T4qILg/dAMlyXTL/MpZdCnv54ws8/OtgDs6yl
pMP6cMQ1/8mE60o/VPlPAniyMUXMj6BSwTh/D4HlwuqlBFJDs3s1/DCnqJOsH6CaxyRF+oV1R20L
nSULHTFXbZXi5+KNKmmL4lpxCPZxSdna+g0VV64QlShgprCgGL8mtUshGFC+s2CdYkEOK7i0SZeQ
nVeDMkKCNFQwPPbjNgjillzC1ItffjBit+hG5z//yiV+5dqQ+dARizanEGU3acK4G1Hrz3rAFJN9
0N4GP45RRchz02MIENuDaJxd2HZJ2szN8AgYWD+/NOfIL+S+YosF4eDkqaHRh5mb7kLn6e0R8N6W
J/sKnaPiRjvriwzHl2TuamsZhSKI+WDXzw8shDMfZodMxcAaMQZ/t5KrTSWx5fnbRsH4roITeehY
KmkN1mdVWeG9Z235kSiEpM/JPxMCCtyk0UU9fhKkp5vhrKpQaQGRSsBP08nFPZ52rHN4fz8fdaHN
cnJ2khz9/1STj95fY67Qgneq9MzD+1+K8IwJI6EKyM/eVERd96uDBWY+ypdvsVGeKgUMG8HXCa7/
jUhZTjqHqmpJ1wDK0Km+iXcPkeWVs8ykEWTnO5pzs42znzHD3cV4bXKtwuP4mfMz1hOrrqFKhPVc
KqN5+Yc5LNZaSZVUAwNY33TVGa+7rT11i/cNIR9vYaQvtxPSlLBeiP09veBjhVAJAxISWYT1HqNv
BuN7sGJfBylHP917dOb15yLzW5nK/8wx7jv+80ezqkE4NM3XjZpht1KHfObbqGUMpMXjtPugL8mJ
U86l9JAiS84wM+eRUQcwZ/hpTF5AGfjzD/IdWnPQbCmZuDHkz7+vv5aphraGPBDm9dxdT+ckoWa1
z5F2WgTnCyC3EBPJkbHdEi4tS1P+RzP9RBIedOnV7p7xODvfOFo+2vAmX4yYXrrC3jBxcF9Vn+JY
cfvJf5AggHi0uwxiTZcbw8pQnCmpih7PH9XsQt7jm4Bx7DfJ7wpHsA93Rp3L+flw0vqAu8IrI5wP
g86wxLw8zLLlo4n0jVro04jCHEdssyB3DlTM35Tzf1z/WeV+krJMQwur+jb3J0hlo6t5ajrv4Qlg
J6DMy2J/HmF4zqfhLNgzbpYHRKjznRCw6/XEw5aWXlCI3MFb1y0lO4Fx4HVkuUiC3+bEEQPB/LU0
ItfOmUrVvaI3TnaBA3nTQp25u+dskjn6nXdCE71SRfKiR/5zu0cyjFdblACRkK+JEI5gyfNAuuqP
4wdzwtSCR6SPKTzkAD0FOBVkw/ACsshYD8M/N24HUoOM7BQ5rbHe08X+S7RI9Tav1USBeaVSOQB6
vXE2roDTgKxc0LJ0iEtxGzDGYgJfwHih0EuwiAlRmJ5QitTvOa+FEwlJeZ98YbrpCJ/hgtBpwwqr
Eq0y7TJisrYVFbIssup6KufZ6Bg7N0f4IApo+LdrT8mokR5tsM6zIhe/0OFWnl4x27IllkQGAprG
D097PWIRF7bhqh1SlYh17NMz9ewJCiua2R/15vpkoHCfTA2lHB8XXA9V8iClDZ4L40ipNoZx9fBI
7ar13y4UE9D7lFd8caR5bisDg77Dj26kUmofXXQshxmaFUG3oh9KoEDFrFNYVGKW6T4706J6CJnk
d0jEko4hs/dxuVJ0UWTr+RqgN+eNeIJw0Pr6QbjRDlZl4KHVxi2s3fOV4fVBIzZG5+ez5l2m9gcL
JyBgIHmx7ipV6a9O+1P2PUAzKqsq22UwACQwa6Y/DemMoB9VRY4tN1RkJUJJdXgHEQukqxlEG4Oj
Nl56QRbgoc2QiiKL9NUREC2tT7NA32uvYo5hHgm86aojXYJLnTcWX8cBXJxyfUwKJeJLgukLB7lm
fwz3gdjpE6FeFrPBBDyNBxK6DOUTmqPUbyhTPmz7T9nzjvm2JAGuXOtxRzLSvtuLBSDKqBJiPtUd
X+NypNDU5CsEjha1v6fCvCtjwB6BAhEySWHMhQ9qh5CxkmqbewpnFxF/gsyhCgi4dlcJ7KhtiYII
jUtsYdVEB7INaEQ+NN7WNw4hcrED6F1d/C+IOM4Ogtgq5ODzrzeA49C+U48g3JBeY2Ucl71IvAY+
mGUitTmedSkVilx816cp8oMrJt3JEzCGYGStIO8ex2LnN6PSPT76SSZ6k9/DPeqP2Z7/fjfUgCp2
fTqv+gXWoUz0NQeYSKtRJsg1Cl+w0YNjOXDlUXOMGno1g2116pg8WLOieJXDh44eE6vMc9ul3L5h
OsU4tG5ZF3SJCrxQm1Tib75TvLeQrrake84vWON+R5+UHtL7nMk+OTn4+GZVmWWvGMJkNzahLkD6
wWbjiPgSELsacahB9oeNV4H+BVgmyi+7AKEgBpIG8HQpHt8LuxHyj3uIFNK4kt1nq5XzyI25yjxz
GMJaHCDHEUAdjU2WwuJLC/bI8Xz8gsvTnUH5EGR6TwlPMlCFysm1vLIBM8CjKlZWjfcrzuIw0jb9
B1QtY4fmX+9cFz16kPTyn5qsu2VbiGf+duHslnGQrCIfHGf3FhGY3WxkGH8AXj9UTuukFRIJl/Xq
UpQ4RbPqoTkjYNumCexsyLWGYkBxHdkDqHGQEaUe6E+FG/993+4/8ZGC0Rtsvnpa+qWu9D4oNlW6
ZYAZGwGETsQMEclDTE59YXvSShwYET9/GTRsO18vNpGdp+7xjloxI6JMh5c1V8YKgttRGrMB76f8
XWCWvkzDMfV3P/hkuaVszCp+0ZeS9bze2mQzvXVdXy/fSXRWNBtJM1yt0ijV4QmK5eKATJowPxGn
BpT1OAM2RfGc0yFpXFNMrb26uISu8ilqfDURjdVa0CSUO7oP3O41SdDZNtDpdy5lep28sV4bQJJh
BqfeKKPxlzpJfroaRUuDYUDqDx4nJ5lbvOPrXgUfrwcQwpLEr6ubJ7Xeh67uCESCyUGTEmEyuPVj
M2lghXSuEkGkCVPAZ+zmSZWcLN7TgDGZvS06lMzINuX1pTiGVh6Bsu4VJTaLbgrRdKzFTVwRnGay
rsvoampVTnFNuOLPPJ0+Op1ZoX99JPuWvUU8C3N5YSmIhAWlWlAmtt4bHeYhI49YrWCBlJ88iC0W
nbhvyCarfJWIPK6jyZYIOrcgReUMSFopIFriuUYs8U9lmGVfWJxbl5hC5EYj0TX9PLJpDoLL/rUk
sAAVazI0MhG+TpWEXAdddDVlrsW+ArCTJSakWpXAxD1OOs4bLPPZQevdVF+AG8Yy2M4pNnZZEZx/
jAf8PCgWHamJF8O8uLamZVrY26b6S639qAc7P+tgSLevTgb69JcT/RI/O/i7Y0hkORFHsD5mLxLs
N9UX4ltbz9ZAlCr5hLsIiaf4t4q7y9s6ZdeybHQDBFpORk6lZ763sWh4RQBbkfyreIoFl6R5dYN+
EiFbZNruivzbDm7RLBVqhM+s+fxIJknDSUZSiIizgJ7SKGBfJJfkufIL47+4OVdg5X8AP6dcYOvG
0y7gaV9+IDpup+zS3bGJo3OC0JPlfE55jSA4hY+kdRuiUNDCoQL2iorWgzAERvuKzvyAvNhyTScO
9D6t0mYOa20K8Vyav7RVXVt8P8bYO1eYRkg/lPxngXPl8OgYV1sHqexqJUjKIW+wPsflrVZikgGP
67yJVqdOTC27RAo3JoatvDdw6INHJlFswvL2gpkH70Xm8hkiXJwRx2YEsb2S9M4NAgmbEap+w06Z
KWfKj1jWUwLJRjigXhubWA7u1g4Q7BsyqdAGKjn4WzZA9UzbzJ8kdDHaIrVYtIZJHIWR2cHoNDYE
OY6gcm8Hf3gAlHWpvB0BFg+Pb+ns416Yhmnammax4E8cP62XQD0N0TsDNl5r8dJeZCrRsvon0uMs
DFmIGsymOw269vBJywLFS1GAbaD3nAqmPcLYZqQI9kk7P9btrJfywTe4WMatUDVqaKd1VnuZq1nk
RPQrN5FYZ7IHNJt+LZY+GGh148JJj81EvZSpOuzKFv/fx7ZUvDE/Im4tTE+j2sdkhsvKBlSG9L7e
ijq+KahaWG+xcaBhe0ox1QVBUejnccVs5onjOAK7EcZdSJTxsJ94bRAv6V9munatg2POZcD/EO66
dmdsCO3GLr5yK2EPSb1KUDkZog6EtDh2uPWF5Zd9tdrHp3582IgxBtcE1nkFsabUyWA5BgGNkrMi
lu6a0ownNLtVJLb3ZIHLTGZhdtfALdNZeKscNTL2Cc2TjBcgGziznkUM6PLkU9S2CbYuhpKar8kp
UGeU0ySxsi+vfoxWjRLaPH6ZztISoU0DXsjE3peUHQw60C8IQOw2iFnz74eLuHB3fsjvQ2PJ3vR7
xSakBVDQkZoK8e7J9scQZhDVLH+IwQltNHS4khnBVeQ/YEkee/4rUSNlVHGUff4O1zQsMLURvgym
cXvWommnjpSkff/UIeMwduyF2DojKc1oj0R2IusBLvfwyIBr2FvQpiuLsqBPvdgfa2y40/ubF2t5
ZdC6ZWwGv1yNbWmFExTwWydFiWBNwRFu9YnJ6rO7dmJ7IbL/VbSr3Xz9DmlMQYjxtkHRTJMKaC2G
aOD0Zs43Q1ouBYxKKLBiyMJgGWPIw3YCcXAWQsQxrHOyiv81uxo3l+I6ZYMxB2rdWk7mQK3EDvLc
8Ghf6XeyK6+RQONv4Vx0dUmjS1AoVqNwsqV/typlvqY5cvkGMdIcwyuH3qaOplPbjRffGFB1Kzk6
T+nbPKFfGFZpEg2ByyDTWpIWPC1fba3EdEunsIlfRrTBsfbD+8Dp2l1DNgwAQZBDATWbD+Tj+0OY
6fN7WQdDwlSNiNKhRDT+6Ga3PBp8ahIshMY1PvHye8xoZXbBIkx9UWxF0OIYEd/1295GP29qX3wz
YzhPodTLg5F3e0LDBHnBGhWrilFucz8g4rTeUmOtOyivEgtxH+dc6cKOEO4Kntie3pcZVjdnZSNJ
D3ikvTNS9GJwYKfJCblVntroUxs3cp7iRG55pwCyq7oZx2CMq472MJ91/LHgue9rW0EiPn3swOC6
pdjHSZcx9GxtnCqb9g1rt4PBoOl2/5GE98cfffhK77RYeSJA/0GzMB9YlkDIzLb3PHQE00BIBt5V
EQ7yH0pq9CT+230RMxyYm7y62BXCZBoORyBS7SPTL7AG83Z4VrmXhnoNgWX4r5MVJeplMGb3+YJD
YfgZ8tg8jPPKx3A0HbAaoaJjZdL6JLu7aVYkCRJ0cz6kOPhHaVnL8Jlolj1ZUJW9aVVKV17ySQZu
ENvzkAPbbRGCGMPNoaK/j6zGNxG7CFNWXJ8wkRmbOkJ8iQHg35tGaUc3k/UYMUX8UkHFcPldmvSj
e5RUsiWJXIou1cY3k3MohF1BLlv4ND4/aA0FqmlPYrnEXwU8REpba0Yo5tzC0EFmF0xEzgHTaHNR
iyslrNKzhB9gqNEh9tnRZpu9laFN8rQ4N0mu1IBY/Y17czrzqV4+rkub+AAf6VMPLyVNh5DDYzu1
aaIfYqNBkhpNFFYjSWN+uG5VB0xFlvSxICpY0emI7Rgp6T3S/unbAaMQ+ev+DjK/i6K6Zl6P4/Xx
NiZcOeqKSWShmWxDu6tGPlAvXzl2xbXE2TmfiyybYSwQcpZcMURWSmPIVvg7p2yb4W3bGavDO3mD
MH0QnAcqfplLzg72rkF7RZa7vwSAgka9cMNnRWFA0kCrvnMQapAkxLdcHIlJvhkgdo1g9Ba3vHqR
9aIVJ+HzdHLbBV9jLRFS0SR6EhPzwOSZuZ8TpDnBvfjs/NmfZ77lWgf5p2wj7Ns8IHmP+tTwsDK1
+trZ3qELWp0bD1o+xBWi6kjTFbg7D/JkC7+SssngRhsdIWNXUXuZ1zVKhrpcYyATiu1yGqysKjBq
FocTkFLkcz9EtK4dWK36IyLOUE32JepA1Ca84HtshuKk2t5831bpmFxZkeqN0m7l4atRWVqFrIeN
X5oyCUrNGBB1Tw548cEsw0jH08IL6ZYvpt8KNVdYjkkCVaDq4PdqEdlL6B7qW3CMi4KtMgVmJvB0
16/FsLXYfU3KVgBGZYxeXm2B4J/Oy/KYrOjY43lAOZXsbgmH/JrG7X17iMkMdsAqn/SnvYhkCFZ6
AhVM360LFuI5lUJwciDBFFAquLhfGe2Q5yqJ2mW4JPff3fZUg0JFToxu0szxOjXJCsZcmhEnPKCE
6Fd/299MUa69AX7dWFavJOcqd9F3RZu8hDTQ+aTzx1MA9ovc9QHTR6Dgfnz948QLd1yPUMn1AVcu
58Z67bK0CeDk8k3VcheouMjGMsRJzw1PPUCjBOw2EOENGsmpndfuVs8y+/0pWIjGQtktuZMTQHHw
AafqERT9BXhbkDCVLX60S+7lzA/19Ig/+BfXGB1gBAOy3hRuQb0wbezw/tAEh22zOA/OIihdEv7A
nfFlTHSRj9bgMh77/lBmp5NulQ/9KkRJLTfGSwksKIdDmHOFil6/LN9muFm+4v6+FSIazIdxJRZ5
tnB0tl3t97c/gOJJtAuTxqCFXf37NjYkM1oHyJmYtoWzZMvFvotUkXFmzzYTqYs2skOi5NMGPmQn
UfsuvqT8/UiqCd7VJ5iv6ZfAg6mqAOH59c/O4OklBBSoo0VBMaIZtqdLPNyeVgAE88xNRo1wUonX
+SPtS0VIzXUP2LuQFnNWxhTssZb/Utbf1UeDz9LHWeNtnpDteVGeB5lIS2qc23qk/E0Hm96Ew3qs
2fiUvVIs7vJjl00myyrcZiqAoqFlaEinzHN06pyaCdoY90eOk9hsP8qo34LpImK38VHtuneab2hs
JoWWqtiYCmyVuH85/EWXbNH+XNSxQ1r1omBxxhuzYYcHLCEtE06TQj7dDwusIzbiaDUxCx4neuQQ
hKvCnBNzoEUp+9jE2ij7H+9UskJIXfiP9PH0Z5p/XJmoOb2XfnLJcc1/v778oCtNH8epHPsAS40m
XUm35abqwfYC66b9ZZsAfz5ZKgPpmtNX0Muv731ENez9rkJ8rdmr+h9fWVxv4V2OEr8oz0+ZCtMC
5spA33WGwAAQsMsClB1SHGiiWlfDAs6x0upjKuRYBhHZJI8VJq4TfTzReEKoOWzikmrjWxDD66lO
q3EO4UxgCfNczezd3rHntm16TbP9K8ClNQeDtpsV+Uqi3zagnDAD1rsrNSkO5MKlmBnpIBmNDAex
nzDo2SbShGgOYwZsxKvBz2ZI+VKrOFM42Cyc2yEN7aiRzPB2w3e4P5Hy19dv4zpKc1Vu5b1QOwqp
xkl/ERu8Xq6qmqjsuLrlIZmQFGC2PrxWPdXg/M2pU1hSXhnwEtniA1pXTVKxs7ioC05eXc1t0iZ8
Ashd69ZeZZYNpLnuaD8WV5XZ+WNZWOWrHOzl5Z6crD6XH17oFxgcgAFI8Mj/1eB/i6nahIMpgxcG
7M85btz5FfM/zyvZQUR7nWiAEUpK3zdPDBY1NVBlcLsnidIiLJW1Mu7f+UiNIGK4H49JExayxE3q
p36fLAw5xjIkV/5HLPvumgSXm2ztCBNLhizPy0kSXfFb4b1d9l5LkeYsZWMz5uLR7J17Hw2EF9C/
yM9m6+J7Dl1zw1GYvudxwF9f1xp34WZp8P7hiMWMQWXTdYRs1u/ro2q1u2m0FxBNjSx0rVYS7q2X
t7bLqwbuiSCs0bVrMgM/Ni9u/KeyArcYSjeC4AWjbt4P0lB7GG/TDDZZWHgxQtL7+iNFyS1e1BRP
w76mA2ktu3Wptu7lYEAAlYPPGsxvYyJI+ay/+JJ54+OObKVgg5Tvb/RWvyJ/ADz/UPcI3/IZXX9s
26kQ/DmJbW7MahQZQF5luv9a9HJZdh1uF4ONozHTSGPb9EeOuYy2vJSxrKrFHJXFLfgzurtucPqM
s80CVT1eXRelTYI7TgwqlgwxMFVNmUQbJhbEPnCH/lqpAdyaEg6IXlwQJmhtU0zZisTEHcJaCd+1
b8iJBXy8++cc0HHDbJFvcaKT5r6a2B8NbCAiWy4ZQfHrAjupxiu37s7prZsugMhzX/eWpdkbQLUK
BruaGua/F5sgcKYGFQbuvSHQ3JPFvlG1vqfhHSp2CA97Fvk0GcVRjq5kyoaO/eSVjnawem7z7+pu
bXwKqgXDGfPQw17NewKhcLatXiTWJEkFa8D8GEp+/n6okH95WPwGc1eudCitmPmOQwvkyLirHwmH
ps9fVxFq63PreaIFEQDoAtuRI8FUJWc71c6sjVc3DZi+z3Y1B3uYXWp1DQiSXSRCzPRlvZ6YwBGp
HtrkqUsAiFYQjMxZR2v20FGQWU+kQHH1jv3jXQw07v7X/YAZoSJqzzHICgNW0PxzuCqDcVuvfD5K
XpSw/8hBL671FT/I9NAfgdWpirAvakSMjNbIt0SrERfZVGPHn9dDzyoeFDpJ2sXt2rFZxZXCnGXN
3caEyCC/Bl6Pzf0wx3RM5dWU9WVBXkbEaGefk1l+BK4Vase/7l1AQCb3M+/baw95aPcrMmQnK8Sj
cSMBlsy7xTXLtD/bkttimBnG2EtzcBLiVrl239ZhJPVlSYuFt1icbq/7GRFLH00k5WqpV46Tf3es
gVNbbqdJq0GdWzXRZmdUd5W4vM7ETt0K8lV1aEdWsVnOootuykx8YU+1GIEbvTehZjeHrYkLbuZM
gP3dQM6fBBtCAWYEIIKpHLSK+FoLe+vQywbKnMgal+zFSz92DY1cP/Rw8RhYNE6w6TdMrAtHrNfo
+CdpOFFq9iVa8EOCeVG1mL3y0QeCGF3x641ZFkhYt05rKnlHXnA7jEY8RMZqrMv71XJHRw3b/q/E
MLvEEmUfYFITX3oD061nFilSayuv55UmXGUlzycXnYIkL0E7qIhsyYx7oYGLHNzTd3HfsGF/qbH3
QZiNYvs5vWAW9G4/+KovZXVY+8rjD107m1c/wZtR1DwLte11WupPwirlW6NrnOv77P0zHymcaG3j
HLl9r5aeqSr5Fa+iauuBlNqmCNSq9kxIlfzzzIlJ4NFairYBkA4YfdBNWXjXMQ+ULaBRtPe/xgoj
2zBsrPdP49Eh6V/vCBLH8CRkRdr3AZlpIi+aypCyqsrGOObGFpOzi1+GvpMtqf18tw2DQ+wXbiff
Mf0vNogkfZCFmvVO9N7nY4b6fYHaodzgpctml7lJEd0jL6/08JE7JNOeiAbQdrWW016xtIlWqziX
9UP2V1B/HKRdUAJh6zkMCw69tpA/o+Y4FO4Xp/F6uytXQNBahKcCGri2M1k1eojQdF3vJxGjCqvk
J/fceyfKqJgKx+dk6U1oVPR0JZXa8QsSwLPIOurGLIEI4XSJTxvhjQJ7NjG9fY02IxjOWVNp8WSr
xCGZodqdaWE+ogpvt+cx/NTvFTPjufH0MlHHM0tXeth429fjpEOlsL+RPLPpG5QqaNDxPTjXNuaQ
biPLrF2Iy+efQUiHPYlgJLyiHjUD6xpCubWsM/Mg7L+OH+m8/1el8JftW39BzuQZiHF9o+MAXT0c
8suFANvDmdCMhgPoNLo3azHTEbxjYBC9L7/7eY3g23jBf0bYtmLxId/lYhXS8tL+wsVSEmEXzQz9
ioB491RAPAUYfGfgKYAFVivUSuGXjQ4O0uEMiQ1dOOTf/vy3x+0USdqE9UFV4jb+OFpWq6arX/5i
Bnv5rvIMVSNfyJJybVTO3OU8cOn1XSzOq+IcfUWDYPC+lwM5Nd1WbluQ/EsmKxbuzzpdgq1TIk2R
nobEQHHOG5DlvDmeLLQKQNK+vtSY0PrA/D4mag5CT6Twy+fbDlGpiYRenbw4KlPJNRBtpK+bOQ9D
FATV6ikjZUtvKkEBWOvGWqt0uQ3vpXMU0r8QdRtAjmgdRZzcyac0N1JpnIbwvXYO9oaQykTkVryK
uG1osveY80srTxeqS6HysZv0GQDkTzuB2PMO3oYbEmqvQ9TQ9zDCFU8SemwCa0tcQ/r0u7+aNyBP
DNmKRnQv5pEUjzMYw+dQu3LwsrEh+iUnIjHVio3RngnbOcb6jJNwKatABUvOgpwrKLH+1+BxY2my
lsGtnN1uoufcwMUvl6buJy0DM9DFHQ2l5g5TSIsK7AqeeDbgIGpDtYlj57gz979L5wNjx7vhI28y
zaf66E3U7Yt1ToMi4Ph2mNOdJVKpiKlFZFxcVS61k5p4RNpZGJST8fHhGnrLjl4Zd8mqKf3x4t+c
ojvGvfMnX9ziTs7X7NSR2Jg5dbuVAHbxP9Alx31LZOkoxvAINFdMqFmaaMPxgijzLutEtRcxCN/T
5CG4mDDGUO/sTQJ3X05JlmaPYAko1mYLsAJ5lKKBXYQ86Xhc5Dj9T2++YZVorJ2CwpFbc44mxAFz
hhObCxfDEsL4GTYYH31W5c7q1pLxLHk1kxEKp1bUP9uUdTRvjBLeoVtDMrD6Dg+eNuORFaGIkh6I
68W39s6P9mUN7vwJUBgBZeUhLoxqV8PNQGEuHb8E7b/vWgv8e5XFsIk+Slq8FnhyUK3tisrvS0Nj
qtDm2JRNLmHC7GOriGB5w8i4Qk2aqhUMIkGzW3vT6+cDSDcYSNc6qpnDa+jzjuxeaDrtKT3nmHEY
O+9eUn0MMCY+NVHbzS5PAa7dOCPsaUnMj45fVfhaQd0o9knOw2Dpp5HJ3nPHLTUra5X8VNzSlUbY
2QzjxagiYvsPkmboEvpowM1UvyqhOqnPHv+BW7qgNSAfuQU46EOg/ttmRbT1QEIChHs0EJHM+aiH
FnA7IjxO7nZyr4l1UOW1LuHh3UPwcokwfY48uSpCsbYOqP+x60vNBVddea0JPLFMRRUL5xX7VVvn
y8lARHcg0yi32f+pljDcMCn4lYxE8E5V2brrrjuSHdRvMH8bdT3fYU6gBIm7s5aEjUvTqf9n23tv
4gb6Kfmtn0hUCyEPt5ZonMROJIwK8Kyc2YiNW2XCEn1vQaDCWh+k+xHwCiGicXTTEWNB1H5HLhaD
9592SuxQpsuHtlpCvl0xk3hCqhorQXfXktSVF8ZaIscX39sfMGUEHBjcwgoIxN19hVVUeK1zmMzQ
RABJNh6V/w7DA7YDGUTGlz6Y7gktdVrlAhHfhR4XwW51YmIOoprBoQxVH9cQHrjpXGj8JHYpAkP7
F2UOBed5amcI+eA8jDqIwdWiJECX0QGJoy9f2tOjF149pZTQTyAMFhmU7NFIdxTgLlMCf5MoW/0K
85I8bAgcUb3aio5w5i70bGMvOWrc8zWP84AaFSSNe8M+tX1B4mHLccZ11Lp3wfhdmPAkkZCyJygg
pppAfWYHbssHCvJKAOiSNbkcFhIW8FFMMkTF1k59yBeOAiOAqDcoptHU5Dcq9d91o8n9SEu1amjV
mNFOMLnGAWsNipwjomxHtFgSj+MP2V8F2r6hdJwMjuNe+0of1VyRZlHBtwNpQ6FJZdgUeSuVDJTZ
g4Q02EEOUuBs0YGyNBwUwOvFOlxfilD+gnKtsceEy687OZ/tE0NbvG/pJ3Dgp/zEwlOR1Pw6ktu4
wQUp86wlk7bOcPcX80koPe121K+Xc6jqmmfU08MYlSBvaHMzEqcH7GwhEcszEITY9/+zmXqXlzYr
IosUEgdlpg3uuyXlTutjh15ll+j2VmdetkkFN1GrD3e6S4OgNKr6/ayhrctMwsQLbSHbc4DqQmA5
Kx6TgPiJuu7xL2j8Gcm7qlarbr5/15+F2/70WuAkmbsj6U9fEKNOH36fJoDq2ZgBJVTC9r+QueWS
a1SAnDcFZsG7c2oTJECiEwo2tMy6jAHCYyxX6brd6IoceXe7kdjzIe3BOZNQUx56IbQvH23EqbMF
NFEsskErH3DxneUb60RwHsJ6TFf+gX0Cz+T1laQNSrrAzkINL6EJgKMQE/c/wFradFfzpp+P0Hhx
cE+Q45q0lxeJcEx0k6JIYkv8ES+LV5ZG0zNxPD/M7I0aJzMAbTuW4BSJ7fIoF5JFEZI4WpK/6lHU
IRpRlyZXsEH4Xh2HwSD0K3L15xmyzMq/hC5vH/bYhVPVZarJ6PJONbCkTALoleNWrB+X1yMGFnpE
2h4oyQAsbR/ptdKvPpTFTT0fdKbndseP+2r1QgCMjGqtYMPUTSfyiWO8kut9LQMyhmuRoPIj42oB
RxYu9R/mlxPJR/Z0oU2fEvojMHvKr4lfLWw8Yh2fTelnj8xl+WMZMw7aOcdCM79kFsVCxW+eEuMy
y1zIeubxfv7sP4f0St9c9PqjbC0mCNF4IW90F6cbCVKsWSa8gSakBSqWJeivhbuPTOoe6o9QYdl3
z6XBKEcKQQpaSFnjyhqrBasadnc2l5jok+Z5V6KWAZv69uZb9Hz+g3J+euBlxMpxtdilwk+LRUUm
ApHTUk5N+kkGhEfvM3BAk/clLc4Te9K+23hpJw+xKmuA7lPg/joUy3woMAWOCDxessE/+OGkJoON
EDfFUx8mN8ARzm/BRMqV+PUYvEr+8wcPf+B2azZhAZhXFvZym2vhaTeN32gL5N8gOBj6+JMieQFX
BUYohAXN+4ld2IOIE7tKFTpir/L/AL2itvKnDLLBhHUzcdjKU2QtYPuv0+0uYUFnh31N8cmQyGlS
v4vnbfxu1kU1vQsk4j75DGtmZIEMgjqfRTIXL5i3Pp0xGJWMTrbxcUYBfoNH5xAvuphcQy8fu5v4
eo7r0uBBgUFCh5GYaa2PoxZ8XuHHlH//Z7e6fMDDgPKYsGT589atUeihgLWW/5ngGY6kPqnA1oU4
oXN7Pnx0DFHlYCRIrN99I8JAQ6I8VdhjnYTVBR/6fihdldnR6arvKF2UkpnT4QWLS3oid4T031ex
xJepczFuEVkWgR+OevzjSS/mEIg4daeYoA5iDc48y8GOi4OINLd5yxiz49zj0Hs3lfEcpr25WEZO
uE4p8q96/DfH/3kJeYFsve9TsXoI6sEFXrJIhj3ZfT9pvxR2SZ0+yBS6bp4W+fknsTZxh0Dg4rLz
JdL60twC2upl+TvpqV857w/4udOt1366YQnFQxtLS1yD5D/23CswOKDpOf4CtlkxRE2QQWH71oZy
5ZfYiG2MdvTxCyjRDIjWxYgsLDy1R5x6+PxxH3pXcB9fR/bx2olbmTrzYJBsJ0RNa5749IMfHnJU
y4/U4ee4CA+0gXkwmFkJwaNqd5K3vw3UqQET3OwwBmOfNsPhMjGKUh3ZBckLRtC53Lh+24M3VVO2
ucplEpZK35QEZpeU6Djp0vjMHFAk6bCQxia8HPSOKjJotgsNZoYFokuC1gt9HxUr9GTLHptzUmhm
Kj4DcHljMnCTA+fIUMsmAEhi3FGVa7xmuc7uPIcgVUMoE0IguV/jNmGpeiRynB/15NylwjK2ATpI
f39gUAStFd8QgcuN6u1fW2y7amdlaqS73+Wby/MYVeHmws4Ztk1SLRiOCZr2q3wHOHzlMCo3haH8
GxLStemFFFf+DZWR7uydy/mO8Y3Gb7Ti/iRp5EpndYh/IICkqrDILhETdGX/HP9Jyg7Ksl1/Biet
0E7/aqwXBlX1qDFkfxMPkSdPrkbhrPiSei9+ICkt9dLsTSOqfs+O28yLZEMaDGHfLHRI2WOtIAat
keWFQZiOt+Y29IE7PTs/Bsw68zPIqAGW2qhrdHYkIoDIExGRYPcDH6ZKfg7S6n7QM37Ckti5zb3S
p8ciGkipetvBajgVzKAJf4crSVrwGH+b3XLPXYU6MvE0QglrDwE7sZOnvS/pxYwy8fHLS+MD2t+t
YeWFxkBuwaD4wGY363lm7ALYXLtfiwaJD3ldxEF+IuenA/f8k/hjIP04yED8gEEQyu+AsLl56gn6
ijkj8E8WxptbxZG7Ub60EheO9kSrCMxkkDQyti2E8nUNHvYApdL2aTsHhKTeNF0OLJSf5m7IcC8s
+qcwn6bSoEag1UnJNVGme1DZwvfSzj2waO0TIZd0EAmgSLEg8X6vyoFtSmeWb3STWIzybWrzqN6F
YR8gOgI4glXGkeOYGES+YLzDWVN3AnJ1i2j5Q58Zr6WJGHIariAag3qY7odp/Vow7S38tCW1yVdy
ErlDO1gAg2J/ge/pdHSirCftKJoxy5N1YeJHT1u5EsKO0VB60HUkreJYB3CQS3eVkSXqzrtRA4gM
pQaJG/2yzq/pOv2WpRJJa9Al+qek1D+1UsZzDm60KyJDOBPSOQqRBtLGowM7BrrvcGGwr5qoKoZa
7HFWWofW9HmhyEEU9s3XN96FNi8xmfH7h3g5FrdZAmCpMWcvWEC5XM6Yy5lBmHy/WxoqJHWlyfld
4dOOwCIfgvUKgmgQ9qw2d831Ln2cJSnAnG7QNLfv9qwtWwOEm6+rF5om3Q7eYlpltwMNdTZLTGUS
8E41x6wChjLlRnZOYd5vTZhlh3OuPlwj1Wu+/7CJy+CKcNyPxcTQINrjgxw6OPLANstc0W3Lm/KI
ZdKPCxOeltIxrRxrKXpww1WvEDhZwhAEmd47yZy5yQplPjj7epvHiv5sxOKOBl3dHWnO+AdyWNIt
9NsDykeuSNB70lLbfPRYD87g4odDy+G3o15dxmShPOg/dnZccW+lSUGUIDRCoSm6SNNTZogRXS9p
wpEu/o27CpdqFkJqhv3N6yqKcnHs1Jl+G0tvnU2Sb4/R0UR5xBj6y7054LD3EGzcEtO8vuy1cfKp
TnSDSuPDb3XD3WLWFZX6jKeyw5b6NycJGrCKEm5WP4bnr4neg+/Fz90KXlGK9LS40NGJ40NP2kBc
3OtSpNRySNUTx2R0PV3h+bsxFSwD2Hyc/9omXHzajcP17/fOkHTxplbTL+LkJO4+AdBLUdCsLcxy
53xg+z7DnH3SBQwvvWdBPU9HprniieJI4P9LURhGNHbVOx6hTYkppursYTK3oxJbZbtLqLjm4TYw
Z0XrlM0nALtvHaRFMKvn8MLaUjqmitwrs43obywtRsdNM5FMmTsERf8fMZHbm+hlzgw5gWJtAUiy
PdciB5opC2vx6/nFluDnDtgBPmZQuT+UAmDkRcW+4r70GDgPhcnf/Il7mgkS5Dvcy51k3+vNNFq7
FPu8XV+krqE86O83ZGo06it7JCxBxvcZm8U3peUZnqGR9/JrKRSHUIDc+s5AjMAnoSCZ6w68NwCz
JlQsEsjjUsbLfrgB/M22UxXN1EKLW9qO0RCFRiVCk+6gK41W4VJlDsielbpplNm58slurf6FzGe/
UTJhoacjM7t+Y1p6no7QgFXZWBKX4fw8MdxwrHPFL7EngAwW4PxN3W+zBgc328+j+Xb9G0ZD/ZxO
5f56schmI63gjd4RsKU+8wAYQUXAafp+CFYT5QDNkY9k7HWHrpnUhfgUe8VeC+BdlW1QYxdA0Grg
b51+uV5zo1BrT14ZHi/eNZKN6yyUuoqDDRRiMALmHrz8xphR2hOgJtg49mjzKcLJA2J0XRMYPryg
jZb+EJ75qFMl+phWxR7LFghbkE2kHCOiR9ll482q+fOkzu3dH9QkTLP4Uwxhz+eoOlaU0kgsImkd
V2xCa8UXaO5AaHckDbxQ1IWq13Ab8bEu9znG+50YaoILKWv+CKFcS8KVsmNPjDiyj3X+zUx1KOi0
88B8yRDF3hO41Op9ZxCQ+8kt4v5xHaNpra4/Du4JKVV34bM+ThAdk+y/t3gHOQxh/FiYp5JlTlPR
G9+iOCWZc3Y3HR4NSdXkW9EdKUldI2Vcq5FRMcJcVXrSB54akq1dqTn5jHUEdbzNGNpQY3Abbg2T
r6tkPK0SPM2MPVLNAGak0ZCv4om4aRibiiuU24YzTUZieHx5bsM26XgNA1gBOQcitPrz+i6+cgKD
UUmr9vVyRk0NyaCoqVqnKnf9pmcJZBSIAHtJHS99bGlFIPgQ+vEzT/7q26SxhX9mPX7PGgehu+LN
xL4d3AyplgpwxG06Cv/e91pmjtcFMJQu/5iZyvaW1jRgTqVn1lc4T4o35JbW322YSCKPOtDRVqcc
XW8A/kqkvz33KSNIh1xju/fNn3D6j0ACamxvoadaF6D7zuJgXbAEl3BaQyWmZeS8ILGTJdlljBuR
osAypwdqJ7DW9A+ZbHqKVL40b//ld/GiwqWVPxZ5G/rBZozQlkC9ZxhORK8C0GQsR5yxaFvppB54
DFbH+oRxHSeW8Hse9kzW/5nJKrBOmAxcZqh/bYUknqHq0sFqDth4J6Yf9fylKvyUqeuPtSfa8w72
Fj27ngfsmE/oanSk8RFa1KTGlSXxdsoOX9WYwERAjGUpGWQhWlBqNEpubgWxeXETtUwu6jshIuZZ
kuiJ8LaQxfoB7eMe8QmOVLB4vbiO64WG9Rdm2vQGUajvEzp6atn8rl5cv04Ov4smYmDyfnM1v8mb
7+9d4lZngcUGKvzOid1vN3zoBO+GgvFQTxpgpPzB2wF+oB9xHSec9cxIfYpIBrxyadRQETE18+xq
MCNTPboOA87sZkmnuGfLQzi7PnkDnBeweyST2iQDNFV02FVIbZjOjN2N1SqJibvnPSzWhfmsB1Oz
9wZVxSnU4kmIuwr7uj00JIHt+YT5P9kRwrPwgcnIFeCNoUMiopKARdZ5hAa3DHexaeHFWSyHp/mH
vqm6WOsvQyd4v/MaTvqyz5m9hamYusrUshL4cH7anJf2ICtQhISe+M90GWcB4FgaSy1L5lj4q/gB
zkm6YTjd/nBJziRB41W+OKNqtNzJnk58Ivz8znSlqsswwYyIDXSneHsg+cL8K2s4o+Pl72Q3shaz
pE1diSU5lMiCoy8eMQizCpbV/EUKRijGhvwaBdjst6PVCjSB4TL12RzifAKO7aNVw2NBWlRuQet5
DkfzEH2fEPtH4zWghecJ/8rwc/JCS1mMk5M39JzijJ37FgksAGM6QQXaj5oDSw/ITVOt9iW/nl2H
il/7W3X12cGkyCGT+BogC4gg9byxk0BnnsjRLajjYSUf3+DpPIGnJjdPKxx1TmHg6HhcZxrD3rFU
RGdUpmM9auUqfCQ45U3PJhg3bPamPG7tSj7YiXp9KYUyBlNmu52KSrWAYq6jkI2PLZvzJNSqeyi7
vdWv+08saIFFgW5XvFZIr1pLDB0rrIzLkB3FJ6WeiOCVIOoCIRJ6UzwC2RL15wllIXyBF5UoUdUH
+9r7AsQrjilpWN2jWlE7Rob73+n0f3NZWGms3EzHcp8GaY6nqm32PTlnmesD87EI2h312G9bolSe
htFgEc1WV1R7UmKcSXgNFd5DQo7hFDCAJVFvelB991QBTVzM1EE4kTs9BAyLA+zK2cnZ66zIvUiw
zX5E6JHRDyIkHeXuqoAsntihpgazXymF7dme1qi23ezNI2Xw+s7tFtAuXFUV4crUDxbyXBnHJbF8
DLeWG0jXD8Gd+sVgNrmuBBmevhcmPYp4mHiPBKDg1cmKzkfpAKITJE3YKJ9LmWhHksuvug7x+Z7W
KhVR0O5QXPN7IH02oek8bGql/NXndxFlMJZjfB8BH90HkLRBVZd4+fYm5csU6kmGaxOV6HYk9tfG
UsAshTNqz+fqXglQzKtzc0Kv76kiznlxq/PyQuadkoIqlPmHwQmRIP4X6uVYQq7k3lnOh7o5FQ63
WwcEtjCIV7H5v0BBpJs1vkXgTVuWWsjx5CI9YOg/ZK3p0tfILTRnDYovUymf3XG1JehB44mWAlKM
VrJQdseMV6jrDKESHCg72LSW9cJpGZDUdr6dBYNwuwukT39KGZgMSqF0jj1yl/L1UurtjMAmSAZS
xuuEXP5fcfWfOSkKVL3ggEQcBpkVxuG7OvGNdjG/mWi00xYH6kaDnIGGY5q+dqw+hFRJ3weVTAsO
JcU1bTR+njNsV3Qc8MndcQmIjN9WDbI6rTpK9pAAN7erHFT6Mh5i1HMxj0ax9RsUOagpBRL/21AW
iQUAfxZne/Klv1rEgqZ5hyCxh2h9L1PnZr8q17D2aRF3tGlNn1mWfnpE2aPV5Ymepacg5/t2kQXA
hBs+uPzqDHtKjJ59/S1lIx2SlXxCk4xMpHkYeOPDiktyxlhkiJr1sTEIudx474SRy+4MqWURD3Y2
ZF4ufrVipc9VJds7kYNKpP/2u3IlUNNz/GwXBQPVjqWfFcYqqdotMxgwWfgq5D9EslwO5jcTvLqy
VUTpO/xr3ivBWSj8jBwfpPtHqlCH5skuyFnYRwNtTdpZHIaFG9kPGA4faC7hHRjhlEmj+2FhnCZ+
YVnvo9i7Ya5XrMc2ElaRfmMK7rlEVzxKXlBE9/vrrQCK3YtW3raXv26bIDdkIIZHBcQeUMwvxG72
pP/5Pd0yds3+Quqo5faNcM1R3Ezu0eI+DMc2PF3RFW16LRwpVezr4yqOfYrwjh5pxFQJ9uljUZBP
F6OhV6Kxj9+dKe01/c9VbHor7pZ3uHOybjgfOBtpBCVMdyZpMhCp9BDXObezJwMD2IoDR67jAOYS
6a+o7ASFwygHPzkJJPmqIxqpvReA9aRXVO+XqPmckM9HZu6vlidLcyeiaVhm016akrKvo8pXVwjw
qnKEgyApZn9hHc6iG95lGDBzOo7fuwiDHgfzjcaxXIyGRYkzeiCDY1DDqd+6eXFgkS4oRS6aLd3p
Wmi745uMbB+xOntDJxgHy+k0UzsZ9tbzXJrhaUpz+iIB75T08X6w/3Qo1RtvNhwO/ryQ0M1WRNxa
zmhq+PrUv5bmYl2sSgmhP+JIjO6+rO+Smj+jr/r40sq+N+dXCJ+LbkpIcHJKc/OS28gmBrZIkuvT
RewaQ7wPBzbvf4oySxgUI0LzGJaXKytXg09n2xYHO2vLUPZ41l/BI2esuosjZN4/63CwIfzgkASF
DCKamRFkdEfWcl732Q7nvxFiwYuhieOYMBE8hiKmmVRQJvPB1kqRwdh7yOjkKgRU963oiR2M009Z
qNsV8JROeiQBsJvdVs6jsgVuawS6ca/uEyteUjMhRcetwipZXsjsOPXHNt3S/qeg0ZoXAkMN7WEr
RRdLN67HRnpI3uiapyzAuZ1hkKyqOjHwKCygR498CLmbcd8wFfGm+mXmLFyt5JxBKy0Y2F9Jf9+l
smbWb/0OZnp1yR+41TfP9x/PV5V0B1FN2kS2FSBm9q3WBtRMB3K55yH9ybNN9bzKcuFtUcCi/cZn
9JNVBfHTnXVR196JFOSWxL/H2Hd8iE238aHvs6YlD1Q2jgpaVLPTGKagt+9WMzdB6Et9E/5eLAwj
aLs6EqKNzuyPP95Jr4SDhNL8wlzdhxWhWPP2jrU2cVTyTSGTdDt+7hGlZes+JQthZoXykszHOat5
uDi0gKiZP6hU0nfbGyxg1Mp3Wek8GZXNBMoz+f0/RWSwTAZEyqFA/Ub5J+Eg21LqEK2iwBL/rRKH
vEIoxysgKGVAzmC9KWehN6DKBLT3Z/tCGrgHegm6C+l0sgr583HRv2Ks4RxCNssz9yvnkA0/+4jQ
p9SQxWJe6bHIXQ3QfCWQHlyIURZbCSwuQWmXIPygTXdeB9FsdjBiM8fk4OaUKMGtYvyT1g7qb0eb
sk1Za1L96sEfFF28ceCnZlkzB6R5PY0T1J0Nh3/PjCFFzDCoBhtgqtm56z2gMbz82WsH4blJdH1P
nJavke4YNUh5Ps6vccsjQYMrdfl8g1WaRW8H6sWWCeLrqd7tvdUq0uKV4zNEHpO/rQz8uOsD2pSO
LFTnZYwikaqAt0T+9mpTN4Zmi9ZPtk6D3NVM6csVDjcQSMSMM/Y2xmHVugg47TcLRSPQroMgbnfV
mzuVkg6pB/l/Y9+kX+xanHK2fjkRgDdie4d1EWFsOF50rK2Ve6BYFUsM+qpO5QxOsnjG8iREjoKc
w66YbYDpxIv3tSF7n+nvOVYuUQEKYjuOyqGZwWdAXOOp05rnGJFikEgv7oBC2Zzn+FQy1zQexBio
/UKU8rnYgtKHQBTofcFjK/Xy5YfuUecwlmoWYpUWj29dbGZLAkD7z/QXs0W9DXxsGa8VR5d8FdcV
iGmZLmQsehCgONr4MTNtpEs6DDcjfwnlvqzFPmTsh9TN7MIvhQvA02IEJdCJw6ATJUZ0weBBUuAj
/qEwrpxWMkw81vR5KNdfI6jLSbPU6BGE3YgXp+LmjTuT9Nh97fUGu0hzZ7tNDLtsitA1m6xzOqsb
w6UI+UC433D2xX4+P2moeG47A5H9sdC8cYZq5PyDRy8N2a4cC+NfeLYGd3u585ct7Lyp+/DV2tmt
YBE9acEVE9sRnd03z4mujyc78MqFlWdf6icg6mbDUgehhnlhyfABnqXbu9+0cKGtyuHa1k0s0v3o
A3zBjZNntTEP6hl1lhmzV3BJEI9RH4Gp+q9CwqONN0zOPFdXEXXE6zLq/V7q55k1ECGgUkjGqMKS
pvluc/gSU7bzezaVEWN6hiSRN/lfYENyKLtWno4ilqTcMd2MvUfEt7SDsvTsrxfeO377UU8nBIDd
ES8hYEByNcGOwCJDfrRTGCqMeiW0Blavk4AFMaJCuLjdCRwIWvdpoYdKAuzt+lkEmbglmsppRDG3
fwe8jyS7ycNzGkHLP0vAH2rWnbp4lHKOGGRpy1lGVhE6uTdW6RfGTz+m9xaisyQ2fXuDGq35euRS
XpKp77V94EFzNdEUulODF/Oa8PTHeX9NHmnb1uEXwtqH/EVOuK9SpzmxpRXqOfIHT3KxG2GysbZJ
mya0oqhCFDdPLQ5gZu5V7P2DKuJJ9HAcdFS/rwpFFsvRB6TyH92JAdnbqrJMAij8dsVARoozTgbN
Fy/MijY1Eme6YPNYjD9kY1P6E5+har9bQaI8eHqnRYAH/I0q3b2nsJ+9f7uM1tkcM31JQweIyvwB
DYmR2SMeZNAxGvwqV8DKqlL62jg+6/VxOAYBmdfKMdTj7ugwABsYy9a/1Xgp9UC3bFUeh7Nf8cms
DlrZJGb0m1lJ5wXvN2/qqhNA7irGwFzR5aq6wV0a8Et3k9CjpncRvyv2Z6yohYnxWj0DQt68QQb2
74FgUvyPlBr2N95CkTphrvnoWPEAsvCRvn/YlPro0rYbIVfAgcGRZcfnQfUS0S6hNJJnUVd5MDMA
3kQqIWFs13XqV7WvMULSQZnpiq7xQYn+ILMnxF+htBq/WgXfzM+fj9sApI7r9NDcVfxEv/+bRC57
WgWdrULgb4kFEohsRtoT4mfb1/SWlFIZXyxoASyOfluC64ag2EYktmRP0Ufldh+g6Up5stSjq/hp
f1celEMYndzudoLURlMJttENaSLkZr9Ut+XI9JBhjxYPhCeafnCIYkDMooy3RvT1eSUJTK4rpGvC
EMgnZZPM4FF6LPjfXn77OGV+pXSlV7YRz+wx8b5PRiFqTFWFyx/IBEVhOkbPI/0yvTk6l4G592ve
AVtTot5ZRFiUm2wvaXnvAzd1yGny+GjNMAq78ITHsB/Ba8OkaHXw6p1Avo8qg/teWDiRFmt9AYYw
cFxKsFRoSmsKmhWMHh1vpZcfhFrSW6jZ+OkRRYa/0rkg3TxIYVC4R4ZgsML5mD+wRaNSscBUBeSQ
TAoTk9SMF9mnjuos9Cz1KgSouKAui7DSZbLJkbNYYhiaBqt/UqTVUllGLQw5niIOKGZQkqS3Sr1S
CKLFS5J0yNF0aifSaTXnmjDfhoynLXPCLw7olZQB86k34bzt0SmiJCj1GpXHwMNMSWpTHdhWxgwO
4cE66VN+bBpU42+w0hApQJR7lodCdAmzKxpn5uz/TR/Iyq0vOaiEZXjjv3b1IF03E1gb5oWummLZ
N+gM56nxaec8me6eOy88AN9AKhJg2+gF93iN6cxVrr/r7u7H+HVOtMa8tkxswX6eWxHEBmS4EjwN
ijnX7WHBA6Q/GJXOTz+cmJ4ZdRPEmwV04b6f3wW2+AnmNS0XsGjxjFuVBdInbl3xe5VTdHIMxxPP
ZVLsUDIDe+ZctP3EKngw4hCqse4ZWVJSHuLsz+h0MPbEjLUydIxq8xNkACSaALmQokF93PnpY+JI
9YpXatfoNk6McMzujhGaI6tugJ6DoQT6Z5xWd2K7Xr+dRF5a4OVYh93TfcPbm/7zVcXSj3MlZMhg
CphWKRlSlJ5MfEhQzv+2j+vEpsjtPeAQkVBa0Dlc4obBwgC1hH3GJqZfnaiy/KPMvPfifwPiDJ/D
a5b4aPKoqWqE/4s012R29UFAno8zillZY0HywxKOeZOpe/tZU/nLcBujIFHc0cEgE/Vs13MhHJpq
B3shlMZn/al7OWvr5YQcTsZyx7qHCCVUQK1j7vo59/rdYhxPA/Y7yktD1EI4E2Vs+2R0373SskPZ
c8E/rs2Vb+kys+wmQcF1pIqpY2sPqonzS6M7GyE4dv1IlBhHrlJtdsYmNBoDV58cFh455OKS4LCL
KwucvA/wgcBH7w7ba2IpKLeU4ME9d0qfCTZcLlKVNpoq69z2oqNjMme7rWvKu0YmBYCQN2rrg07S
pXuLTeK3jzY76lp4P/cLi1LCh2RKNXbIgSCs2MIFx35IgUkoSdR7sg9t1mPkafPQ6Y5wBrOY0OnC
o9jod2yO0e05TpQkJalGXIcIif3mvI4QyJTmEchfT0JDl/7cSVNcS5S5ADx52ULMN0gUOBiihGhx
HIDwQ3xO1xCxFPrE5luaEn2RHVNoXPXoUGlyqxig43UsNkZnA8i1KFAsSp/4hJLg05dejIQhrmaJ
rMqHEvcCEZud4xNGH5oVPZWjmUgbWA8kWAYfolb+qIUp547qL7Tf1Wyb8md15H5u4liggB17/KOL
UkEMN5zovN+H+O0DG7jw1+JKjqDORUrO8s2rqYx7uYa4+GBJj8xFxB3E8qvwSRAeUNP8ZvPJPvwi
4Io00TDh+LulQISJSxcjRVTm2cETJ2f8y37KUKkKv+vGbxaSSHd1x4fmdv6wEiFOLiIWD5qgARun
UCJcpkiioQe/dKWRHEKyScdDxtsr5uPEQ3amiWHJCiIQOVmhxgjXfsbxqVJWm+VSaS8lz+8dKzCn
Cn0QjUaYazBI03Jqx7ZQxnqdW8ySfcrsvmyOrDty42SrEPAYg+26OsGvxpQrxHdsFhMYWhoByIaZ
Ls7vInX1rziDH3DQbNzzQcJ1XV1I6AnMRxvMheSfKwMFoWJMiogEcDV1kWv8t58uBW/QkT2obPRF
I3/riQZouAJ8VvqqnzJ7FkrvsTWyIvWbpyt52ze92/XiGDri7YuohlhF0MlqCjbbX2zOyKnq98hh
WyXlGvuKUZI72q/4Azy+IBj9OMAJqmKKnY+g5pPsDuMrTKRTecT4BZ3vmSDmC3Nx3QLTLehxZyEc
vxmXQnLYMWzDH7Q45U0gjNEhDdrnrEIwkLIwvUkPF2t8++NQyh5khlr9508zI8k8e0yHBAAm5gHm
uBHuIVbvtdu2GKk0KKbP5WAmq6RLjMrz0KSjwZtjUBN1DaCxgqcimCHlnrBRgWZKMa01VU04/ub3
oQj4hCHemsOxLiv9o2X9+SE2DiLxytXGptIQckwSk+V2oAJTU65RBa0zNoE4DQB6A2kj9OANva7V
Z1H9skBevR4cDKDKiyQ9nCpLvF2k9QIdk2ejQSRWLhVqM5JngKx906Nejq6A/opH96LgBcaCnsYN
S4veDumspMgeuuKM8l8bsyapDTe8Th9mETbwpT1Vw4HVRYim6WAgewetMsBNWWnKzl5vF5fh1j23
aVUHDrvTPyIKZx3HuUPvAJDNS6vmwQsvRyskZTHLq6A2vd0cGogoSVpW4hs9OSCslDktSVTEMoQa
IGf0fE6CdAGWX16VOrdgw/LoexwPkG3KPo9cyIQuLim9TMOflZomsXPsuz+UhD4hyjiIAeSMv7k6
98pthvPXs0aVdkBX9qyv+w1yzkszwmhq4EOrxzgQe4H+/NKZTAthp4m2qECdwBwOZFY/W42BvJsZ
cToGEDSFltzQeSUpTyxOrjMqQ6vCbcHr2FBkUGMCicQQGgYvfbPS2VWLeFXoeDWXsAuo8c2uWBy/
lqI0eev4lhnLaniRYjQxryc9yuKoIyLKxamrSAXeqNiZbT601hHcIA+RW1n47ogPnaDLs0PhiaPi
lH+iQiEP7CJqF0nssfjptLmdgMAIH+/LeNyQY4okxOUYTwBKJvtpDbCo1yvGwUxdj3Jar4LdnjOu
pCYWWxCmQBagbWGo+BEqfH2eE8qUDZ4rtGhDIuY3qbpgpeL5tLknBeSK5sTpbwf2hXMoh9wIjVRJ
rbTbqA8lMfyr1mzuEAJ1KghEY7V6+Kw8v5BuktgcSKKBUg7sDZ8agN9nuQVqVZYob+tSr6aX2A2T
HYmFwGtDDdbXxbrjclc+gxeJto81GKbsDqltX8kr+1B+vsp6VjqwUdHT5B/qmOTt/tMyC8N8SIzw
cwNx6adS7jy5B4yLagugDFE1vAfN5n8OkJbDLxTqUj3F98an2qBU6AZaG9vqAqS5qv0YJBG3yJnn
EL2G24GCg7JTquB66xmoG05b0UuGPNY6u7VeF+pPzsTOi2UXF/YBfIBrbkbjXZRTDHbU1tHpKmuw
h3emRIMO+kpOtuXcVx8+lqUD/GwfgkTJ0srgw8XcIKm5qam6X2pQnQP127cVAQXZzitvNUqnz5vO
Bq87wFaZ2ZP3G2U8hoRWxKWK/2vdvtgLnnhE+sGnuwbjCQxZZ6+rHxu/aeLaiHShedu73t0/rysg
x8vIetSvjbMBASd+5h0laAJrjIBD/cslVJ8GjTMBZ9ClVGT6QF/F0jKFVAplfBA6ZdQcPkTcjKlu
ysyJuFFABx4jJjiSFp0RF7+YzKCuiivVGp7IudPB0fQkYqXC0dd8cBP87K+KqBwPMnGvcOpEeJBG
jMPe2maaamEfgV1IYs+WbIhE7jKwibghsMZ6Oh3iwGEDy43qGnPnvfuVQHTqEPTSXm8jv++gQBQH
zUrOL7LN66K2pYpNww07QX9GkPPUiBRcfv9x0dM7rxLHxkA98aPCE3UAVc8SvHcj74W54YDsXpS3
JtPxzYHEj7ZWt31T+mScmhZiWiC+QclVUtNUCeCK9w4ykcBdvNkthJIYryIk/cbqNGDNDIOZLvp6
CRyfOPbe2mCUW3pqpmL20cSQkL8LMbG6vqIucN03h0UD7Q92D2MG24mftRbdEr7ond/WKWxFYCRz
1531pzZkw/UOap2NuOwRZkKM5YT3XWIKJU5jn41hhsmx2h9tHlhsdJshNfS5gSzcWHlDuplbtiSq
WodL75o7HepLR1lRj2zVl6pPmF4Nb+g2qaiFFn7nF9aKEp5URrn5YU+cnyRSXhOUVXal0KH/sqnw
G4VQRFPv+8JJ74UyRyLFFzPWJnIaXiWYk/ttTeb8K3oGShLAKOSPNqLaW/Xo6P7uyrhd7J/ceeZ3
3NTLaFK7ynAlSYnYWoejEIZMyeZo+IJxkD6xB/GWIfeNl2t2QmEhKTZmbQDZTVkFnhRcQBeO9ZnD
YirAyr5Rt1QmG61pg4aPANa9OFuRfE78eJ5uQCddGVZodrWGXy5rGtZYymImUYUL+jhkdp19h/fd
ONPg4zCjcspwj4jpM9bvy+mcfP6dYh3fKTk3AVgii1XLw/4vHYLkQdsgEoEjlIn39sSpPSL0Z/kS
u+1CC5QaT41XRX+PypS/Kr31bfeRBqaDRUEQu8kkVqmMitl219uBt7YvtDMQCeR7teCQcz495DAf
G+/yARUMVwj3FbwqCIY2Mkh70TZBlImQ+lXvh2iAH6jNrsRA13zLgA0t8/FnwTkMzzj157/AnUw4
XPonCp8kCpyKD8x5AhzvBcB7jWWC8m8H6ugA1FEvJCSrfqvFcfUCYbF5zxZi0yGW9l913LnDiJVH
iBHpFckxptSVC5N2qKJn6/R/cJGwTZ1lwKEBmjKmf/XYCmaZb5rBanNl5ENn3iguLPa8ZMYnArYH
PTp+9nIHeZ9YY9Sze61gyBlSgvSTKu7kgknDC5xFAWxfpETNqUlPXqr6DSpzW1ucihUwiYfUUkIL
CGeT7yaB1DbiG/p00ANUjfJOjTzadTHbtZODpkiO3ntYwy43o5OYRNy/rfxRbBL43b0b/jhjlHmm
NY5SPeMHguvKngvjiKIgCvThTug08p5JP//z5f1qL0bt22CD5u4FAuVffS08ns3/SvaQ6HO8NtTh
DEPrd2r6XGoSWyZv6Oor003WKfYorJf4XCX8ZzLsFLBHkkVLGq6d+CHh52R/JLY3uK3qPUrOpvwU
S1pUqSob0L/Pl9m1GnyrrDPHMQk05n0UU4R9bY975n+/pzGfIpuMFAv+LqRC6OFxTjp3yM9LjKqN
o7Lwfwl1y++g63kGNYqNpn/TYwQL8Jitu5p0t2yt5jLcqUa6150VyC7mrzBpRBHiv27QOlanPbMA
nva+3fP+U88eRYs7ktTnPcz8Sp+7wN3fJQ6wXt+HW/3k+kMO4dRZcnt22RMnnB/lKqo2K4izHRKl
PcseHStl5TgFQZnG/RBkw2FW7D7a+Fl55dGIty7Q26fH5WDUFJLwQ/H7nGk0bfjUycj8i42QpTZ/
6g3cV2sxUZtHSVJEz6BYr9c5T8VfJFtyGl01cz5netBetgeuwkTCecMjg4Q7tc1otfFq1Uj5ZH9L
QykCXVevRy+Vp5ztnCrkVHavVxe2UI2X6iOMcnFKTXGtpnKupa91YKFWFRkRBLOP4px+m/8aeUQP
WmllNgcoJ4W2CLX9lYUiSuL3SpWBW81Lot+wiq6fTgTCcxPVB3v7flROMejTcg1lgqumuo6neN8i
yL/xxyXvGsrnNabM55SqwvWfcyVe1YrQUbU1GcBjKBjBph2GAPuGK/3yckICjVzc6UBPXWA2GZro
933XkZGmooyf9Tp3/GFIlIQ8MZiqHF5pcNoj3WcgP2Hy/6rP4D7WcoXcOS3SKSbyi3lm/+faJUpR
7DVeG/KlG14podQ94Is2n6X0XDLN3SyjuoOepDXY5hmHsd0S+mPsqjnXoJKpHQFxa11vPrllLFtu
NikLd7qr9O2gdi3WIty/jj/Hm2Ds0ZSqbPiloiOCezDEtg7nyRovarhaW3+xoy2fpkBvpn/wfVht
SqtCkzhHsQl/Gtiq/khPRmJxb0KuwcodvGZEHl4Iblsfl4jhxUGc0qVAk3QfAoieYCrZKltk+Zka
YGZYaRlQ4/mALbmBdpkzED5eAukjmkso2ai1RwgZEXbLevXQ57kJjR5qtv1Jhfk7vV0iposE8gSA
6Iwb/Rqa2BUL77gJRyRuQMI1jTSrC8oo0ACUsyeEzfUGL8tndoKcdixcxGZscddQUyXAfS+TYpwS
eUMf9gedvm3MkaGDvUpoVVqUmFt39Rx+dVepD5Sj7Q0qlAg+1QqlqeH3ZtRWbsq5TxCAWALNam/E
kr7EMokADqEEYkH12vO5TdYgChZXh1C3qYqBU93cjkEmEf2tY5jDb1ooboN/a7O5cN7t2E61LvKz
PjxehhA6OClE4U1proWqPq5i8TJRuTYIu6a4qkBDDUJ7hoqjxJSZzZvmv8sAMhYyhSLlToKHgUeo
/6XQe6iop6YC2TOMsXU3WbnHuRHV2ivXuSJsWTozi1Xuo7ZTRJHhUW8wJ8qNyJZtn2nItJ7ARCbj
Z11UmtvzdNK5a5n69x3pLAXhlwcUcsFwkn3Bh7bbAaKJayHRhA95Eva4WiTkDggH1DcjnpP18Yn4
xm6AwLUV7GEHZpBWWgWFbswzTrJ/GshZKU2lAdgAIMOapDKRmHxNOByw6/AgzPvUb3tvcrk6Gs2b
BZ+5kKsi2GboCEXtyo0C+MQgQ4ILVxmrz8apEf+TBHjQn38swJIMG+CaxjnULjexd8KQpUu01Cjv
6xtGWa72m2sC/9Kn0khdqQm/d+7mRdYOxRiQCLiGkHCOVAYaQ/spJGVnTLCpaUrEnDJvvxrK4mkQ
ODPoFhUHbp75ATJH8V1sdQj5yCbma6jMJ/9FCaFdGivPeY46gzJIMtCK5dZj1FeNGEUOWVQwkfzd
/JfzGpiuO1J/M/hlkpxqRS8r75vSk5TzsZotJdKVeEa4j3HGb7ShrtmU3L5YepWW/tx9zPBzyfBo
S157dHYPU3Zr3x/850a4aGxzQGFflLgGW3uVLwB1AgT9sUNT/EZI46iBMY/xgUDvTT+kABMATZcN
lgNAp7CJLQPqxoQ9hn+KWAkE2aC9JTdS6yw/TD2OoFgPezbDdtRqMP2LH9QYYbHYXv62rwc7urR3
SXc0fJmJilsi7YHQeZY50IBzBhXxHXSQmJL5NuUXZD+13UdhmmBCGkKZ0+ycAU50vP0gdVbYjRTo
1SbZi/07lIyTNWLgPaEiNaxgCGna7GMmeAeeNQoRzPpl9wVfpG4cDlVoYt/e/EFTTwVTRjQNgddA
cS16b4che38eu5DYPvuk1HCZp6PLrwVElbLij9eIQU+PK3ZlaANvHnO5raOGif3BWAwZsccfmxm4
9U5F8nhXSqoaL4feGIKIbnANzUJyjhLP1Ft11JAOawNzU67V8Sw5DxBdUsPJodFdXjSoYRWh8iz7
NQp/Gp5O8vI3HTZUhQjgU7EcEFHdaur+acp4AwwYWZqRCpDbWPnWNsksk230YLoGGeFTwQHEXCia
ma7T3rpUCh4O116T3Ftc/75lY2o+m3DRntvaIW35iVoVy2rpu9+3kkJgPg0ONhxDTgNwYBZzaqej
9xID1ozgHgRunppZvWksH10lCQDGKTlO+GVsOnQqh5jxqPWj2G71WGbHiJF17Jn7Ruau9FOWam8u
Q9ulGW+9ZSdXGERMk0b1m6hNzbc7pK93nzfQ+CEZVJylSIfZt1J2ZudL2ThykY3YxZA7aDNur90s
3Vcega6EZHGoCegc8yhEoQarHid+4bp0Tgq71NxhfE6hDJYM8hwopSaWUJ25VEDo9OWCBFa8KOLS
QOZbSQ6ZUBgpa6Lnrl97vZLLx9BSXIHFUfy/Wey7I5W5FqPCkzXdz4gt6Sr64zH7Cz0lPAykGWCB
cF8qBUa1kR+3um99V+bSo1x9v8+Ggjhli7F62cib4uJYggZqeCyN1qZ07e1GRAQMZRDMCoTU7+53
du0wymGTAC/l4E5zlXihSodm9Em5upRx4MlOqeIvGPJS/7QrRoAwqTTUbhvpxR5uaytur8gBgY4A
rMo7DpDz1nO+8YnLhAlf5pnGi9+CWXCbhNc7tARz5xV18LuB21/UCXIRodOOEvSpXkLGf//5qiC4
/hWfCUx8VTKIv2nva4sP3KksgL6sHdgz3E7qFbYzqil9cEdkXOqjkHvVWYnkPud+jfPZVkG2MNZx
1NqdkgfIsooUdziCbMDxvTxE89uSO+LFVlOm5sPRtDSl0l2nFqTu/sqBv5uMa3soQFOzIL5QGFih
OBL+qRm9aJDKSE/gdZi7Sie/oWJKOecPDdbzPxbPrHyKzaYrG65OcHiJl8FPsiaPQydeegQt0t5L
VpLuai3AbWqlPUROXgmipPuvEE4+Gq/ACGBUw/Q6aE3sZOYi/yni95lGb92lnDKHr1l38LPr+B7y
eYoQdSv5jcVRilgzSHvXAgDs8gjq2eUzQUwcAdNFNKU2WuPTbNNKJF/BMT126EV7x7mcjQCQEjQ5
vosYJQrR9iWOPkmaP3diEMFo7Q6nZlDw8YccqJuoSa2XrQiDUklFixQFZeiUOgiTQq+qGMtEP3GR
Ps35aBycIcES45bDXfRC2eS945F85fWXdeFkQPjy+SDwiGyPgJHLYmBppV97kILAtNAhDSFtObxy
hpWqRh1Jy76R27sBq7/F3QbwkT/vWJ7iiXi5UKggGHyf0RkQqEDPP7ql0khVDaaz2A3K0nqAV+pi
JCaQwrULhEynMX69dj3FP6QEbBUTPxi18lJl7HNwvUn70sPzJWfuZV0VuGe6FrSPa8NvnwdZsti4
nW7dByXk8YuXVAprUx/iRsfqcqsvto088JgLPORthNnCoNpQ35YFgSDdldaoW6OdKoWdRr+kOGIk
dcbx9K+AUuvQXU+eTPJ0DLM21MCKlBPT7/582zSqXOWqKGu2zgZ8lVRXQzQ19n/se1zRE+kRwVt4
n3gB+PYtMZPE3j2zMO+FYjUt3HM75xecQKaoZw3cOcH8GQq+Rq04ythPO2nw0ozIYgzX62qwlhQn
T24kmQ/pjDqR0tx41InDGE2MtOfrF2i3Vjy0oKkKuEN1W1wPc6Ua9diJ4AUf8Qy+c9gMWYgq5FhD
ysOi20UhOo7ZU9lxRfyEVqEUykma072uRKuPnp6Ix7I4ZFfaZPtRAWDZcOF7Uuyf/Pqvrn/vx20h
9xGgpbzp+zUVt/90Uv39F/qNXSVxipuBlGSLB6qgSigN8D95wdSwVvd0IVr2D5lzjoicYVDJHUWK
Gqc7ijsk5E1P7S/40nk9Rp1VXw27mWZVMfoD03SOGS1sQiobm7hRzTi4xqUtJQKmGDZxuIxjx4FY
/7JaxOC+AiVWysFXLNRTd3D89adWPsR8ddGKLJMegmCqnYkiiYdOTB2LzhrRoL1JdBA8pFRhi6tt
vJudiHLmyOEz4HUezvOdPR1Lw9l2ywJY19aJ/S8LAfJP3rTlZol2a9q0mAfeJugY7dEDNTdxAXhd
Y70qrwiQmEqUFUtsqMAwvPnfJlORVdYVP5S1bwL6xx6vquUDJREoY6+wTM3/j1sT/UV622Drzqjo
mAPJMg68m6lykOSF/dYfYP2wJRp9V9P68671pjk5vPTtDprovvrTwNuqWCKkpRlxkuc+LMf8ucYB
6ANWXzx5ojb9UyypEoRpR1UBHwE7DGZ51ADrFKiDWCBGm/Q1bS4aAnN/XRBP+WfQjqmSQAnMtnnj
tIoGvcEXNHv5L3wAmv6cvox4LlahBSqH8jqSR5Ye0ikGwzZdbWJbw1XmxEYGUisA9e9gYY+0SVSl
i67O0uKRkvoO+TgWG2H6jVTqaRebnmYnxNq+GizBfAZImeZbBzsmUtFWoxlyk8bGc4XCAvulKEeR
YoKFhM+Eia9oEmlDLOAI+awv9msRanzN0U+8q3dJpQPj4conQ2ugS/yWD4vFrFR0/MGQB0/dCj7g
bIBRH+yVG6bnjZL63MjUm4rgqVgtayPYfDVENA8HoM4Vr25XNhjWO1nok7GAAHYX5K53ZaS+s8kH
oKwo0hwTEnUuNwIhul4hctVOF7t/YcaRpsqRDuGHAvhGwokIRT4y4srY/70MXEXR05XUh7jqjg3/
c10Pj2jcgAmp08n/RGvRDkdwmAcM1COSCx64F+ZOjUlCB4l8CPv+YnGhcwNSgTbCesnx9A4sbkSn
0IcSGzfNZLXf9Wya7mFVyKL8yZh5AeTlhag6Be/Tq1N6HcZYvEOY7mj9p8WyAqWMUxcEKULLL1vu
CqXI0thkCkGa9n5Cqo9WdiuZAfnmIXSyKeA0FN/9xWgkxL9CtOrB7fMc26/hsST1VHqvyD3uaB6w
/E4fdjS0MTIR08fuobwf1nlVQ3F/UeGtDsAku7qLD8RspKn/JIA2KoNkmp2lVh1M9tj505W1BYho
qLQJ5vPToGJG7dQZCKSNSEh5k9ReKx7dw16RUMO4DAMuGEmYirbbBZQqllheGV895GBkmwMATgSF
MlJrECdwAew0iHQQAPxw2duHwyKpq1GK59WR5QlqrFKQSTMSXsWzRUwigiJ830uLPiOV68X01VPl
UreWDji4lNDdqLrNmibjWhjQ3NBt/kyotAPYonlDQc27p1qpoej4jmxNyL9Df055ewRd9TB8VXao
1FTCyKr5Fx0/2tHha9mqrqcLVGseTde8/UBvZgHUjJv0/5C1kC2EIbVvV3NX7nSc/1KPMrhGiKrw
5JaJq+zWurnKaUF6h8cNrzmOVDlv4CmpV+moLS2VJ6Ndw/vv7Trez/jxJ79oWTi8sn4gHJRuybjn
peXvol+GRVCLX/t43uFg+jEK7P8C2qiZGkdvwCOJQ5/z+1FPmd4mtkOVhdJmQHAlvUCej/JIb1jV
cOxZ2KpDBBfKXCTfGsMGOcmgD4T15f2TYbJixaI0s9Z0HzJuFime4+XU/gfeVFYRtfzjvlTL7fEL
ugpbMWBF0QYu9FxZY1VKLZ30JAQPQHN4gkppc+ohpS+G79UohzhmxlswgCidgCZnYosd5GOzkWwX
xqEu2IZkGSToq5CyuuFZ6O/PGQfYlvdFpE/LTak4aYBfKtvaIHAI7kscml436FDduibUQuzD6Aij
Lyl7TnDcsnv3qmnxYlmZ9f1AMVAbfjugnI46lboU0/K1KP9jFj/J0LLBpIzV2me5GUIlYUihZn5p
qSsjHEw2RdUbef2VFOMbQXUyQDURJ4loPiouBpeATmPGy44jaOA0F3zEbKfMUkQE5h2Q4xEPvxPX
BKrEq9nrmau6RHUow0rriFq/lleP6++Dvk1kHAAbUlFgwixCEEWyuD64jtUHpzNTgAADv906bja8
Zenq6ZJ8mSNwBUMAANhKpkrlkpVnX/RHXVdlNV/LLVgAdVrwKO23NAHYSiKQllEV+N+KyKbh8XBs
8kzorzdkxCJ+V9Rs3EEMCfMc/wNvm023VICTrJj5Fo0QTRwnkEwic8mc23gRBkBFxKCf/T2YCpTA
6QM3/NbZmG7eLeJs9b01UAlfxsu3E/fKvAeI9sUWHbJ7OpB67lvXI0D0Bt9KQjk/aBfkWtEFfrP8
WZ8kXO59B4DOPoa1E+PvNX6cMUS0KrQ4XPR4N8dGKW0aLkNsL7MmpvjheDmn92LEnyt7yWMIV59J
PXj81D0BnfL6WN6nfzl9jua56lpa4HvuXqcO22+LhQ/+k7GEBRyHhwyzPQaevd226lYpOjXclyfi
+8H9D9hEV8uNQXexM34JYXdAzDtomO0WhC4QHN43CWu5n9qc30IYbRs6VTYDlQbsnajUhVSqMoJA
U9X2SZs1fSnx4KlTJni6sha7EQ/IYAaVJwuon3U929n1F2w2wXrG9OzqmY7IqoyHZNw/SFbthPX3
e35KJB8uFY2i4LFhCUL6RppTztKX6L66Xjja7xcAwEZi+RI/pxJ90d9L5BklrCqXBekoZZQwCgR/
yXLHynqCzCfiISp55HFthSrp4NIIWmamH74QDeXipgx4flPXTrXuQU8WoiHNOBpgXkZqQK5//6Bw
NgO2xeAnnjWJ/qYg8J5YFVMdl3R8t2kklDHWHjfcdiqEDafQdkDf9uiC5SeZ3Eky/rkGW5DahlF+
OWWNo1gxYTZ8bbCXkB3f+xCyY1dyFuXgGixKif9PMU9MWswL52bNkdqMTtrgbDamxrxa+iVUDBML
k59cRrIl3iUNLqMctYV5/CG5CG0HvKC5kZuvBtneTlkkSjcC7f/rj02MLgLguPCgb/xJvpDZQY8D
puAAZoLS0OQJhm7LY7nWDIIpQpJ/cl9mWoxh0VPH15q8TIDB7+C0/FoA5tYDFGh0s1eXeYyvOPrX
I6PJ31jVZlm+Xes34bibwDmTXku6uejgtEWnWBwu979GmJp6v0OdAvK8yAC2+pNpGMo18Ndbbis9
uUeg5Y1C382vxRwnRxBVkQyEP56FV6mW3iRKIkc9XcXAEZXnEnayXIoLCoYSs9FUbpGzXd1J2O3Y
Ch0A3QlLUe2gvZg3zx2PVSyagt2eeJg9Elm9cpGMc+yFQU3Zbu784snEDue1h3d7TV9JNNBvYMDc
QsO51da4lXprCWJsurMkuWWX498LQfZ/tU4T89nyCDdHy5iDBYRL/Vxqwi9TIJubAOD90mBEzZA5
r3lM+wcs9VSYY+E5TYNijsv19raHa75yDiQU8AV4S6uatHdBFpugZxFe/1mnNbe2k4pdOogIjT2r
cOpp7LU1Wbnv39i4IW/MeXJlW8fcH0wap7Ys+qaDHmYnOdasmaqPUCgPbXaWTiGMw8XmMb7KFtCV
8jaaxBM/gRWXPC4oE7rqXlmhLKOuxbf5HeLyHtcSshfSElzSaIXsummsUKPWzR01Z4CI7y1Ta7hG
DCN2FXQtaziQA0AIJHmjsAaYYnNPZHl6Hwc/zveD3ORem9QdmLE8gRU6nAyFa+ad6XcJPhdG9J4C
fk3cxJnZk5u9QNpbElYe8thklxEQ67VQBZh5kWNGMH7C65pNnPCM6gRqoHkVFcJHzU6HLPochTEm
1Z0uNS9qj8G8SaEtruJRaFww03Up0A6kjfUtcd8QWtYxGC097pZoaxcz6PGuxEnP/jfQhVO2lR12
QUlayb+Cubm4Q+INUTRDPs+IDqqAWki+ADLp0Ex7YlXIMmwJ371/hv5N0u05yShTuoQHYyqXd/Sd
rnsvH9G4Y9dvcGNxwd0SFl3sOk7V1KEr57c1mDXKgTXIs4Cm10YJRto4I0pbc/IgpHZeDXsRhX6O
FX4UpKtLoRE3eQX7WYrs2ugMMoCy2Q2qLgwecMoiYVY1JESPP+rLcOSwPkT1rvB8ZaTqhTL58ghr
MZDPQJkCbHRR8cXbu008pDcYByuOi0AZS1ukx9sB6vbDxF1LRdNw6+RbiYLaH966rqtmCh8DKJqX
Ds5PxVYJUSOKvGG/Byc3SVG1dMhD8XnYNcav8uR4MKwdPPy1aovIBrJ6uFjfTph9wl5GSHYM+FAz
Qp1nu40ALTEOt/4xzKhzhIDhW1MBQHLjwHxvEutu4C1hdBtKKhKSXx2s+mJmYxe7px7IegWxon72
vZ/dEL1W7PVsLY6A1MiHVZU97lvwbEE1VrCJ9i7lhY6eIDy0AWr9WoVtLp1UR8WB8yT2Lz20a5pA
xhhOimLzVyYXCFKUcHG2DKZ3JydgBOX52AVJpnYgD1dj8DqZqekF2JdT7eXHxU38zsV61rsL4prf
i67FjO3k5fK8w6vKXH8HX2D+6m4GYTPeg7FULXJe8yDCtfdRxjQBvF1ML8XOolOtTl79DVB6jn50
QyZFuM74ZmqXOgZn0NVtaE4VmRxuxAA3AK1k4OLrcyS9uJm/LY79O3NfGuXCoxsFR/dAc3E8RN8e
K2LHIph4oNv0hNyM5a+fX1ObdB/lkv9T3xknWhcJ/VkD+X8msQ+D53JlaH6umhsni9aTpltYVBLD
U8MSVkakegsjcQMtspjd09258zglFF0I0rQA9nFw74ZeTq8BPf6dHHJa0kfwgj0dNtMjAxexn59h
e0PILUew420qmKJXe2/b/knL6caMqCV3ji8soWEJXkEecMSikOAkr8yLQTKCRnTXdrptpOzz1ZwV
hsDxFHvqbHldf4hG6Allzk+imjbgxlTnLx8ZqYmP/SqfGB5w08XZFI7ljXq1RD7CYLvyDb8Iwaof
IQW/L13HvRjUqMLG+JQ74my09+xN3/a+lkkw7wpRvNEu+Bkgi1cb4TZB7i2FnTQCByhffakwDI4w
LBfOfL1o3J36BqjLUj53BagDxjD2KxOyp6JHiVNMKf65mQUHkyLPIqqmq6MV9WmCmiA/eJfyalbF
PfabAuFnrqYlqphKDGRupuzmNdShd7Eea2v5u8vhFB3AQnReuoUdA/3AqyySwR7+imoxdnsNbnjJ
r0hWi08ZyBQfkP42SHoWfnhy/uzSJxeI5vJa0sfE9xwc4fvBykRvu7S9fwmPR40seBzLSamOq5Xy
uLR0Gog3C8zfHffi+4JSK3e4txV2F3KpLiKxuY3dcg3Xytk6G4xa7d4YVNfIxguufmegu8Q7B+GW
nPKXNEwJ+a6JMRvlmIx2h/04GoyrTKjmZDw5SH48cRrAcNv4fZUU+cB6nQzY1RZdgS8DQwis4+MU
zxgz1pi+/+Lu0c+Q1/FZMh+ehStdGu+O+DRJAGiG0bI4hyh8hqT7WeAdAhckQayI8Qmh3OapiodT
5UGegTfA6MmLOEjPULRH/Z8jm5+xSCkbgbV5aLfIKUlXIpA/1D5v2zoWKyYKJiGT+EoVKYr7QYGl
qdHHCvVVStEHEQz154V9Z7d5yeqn88Bdsyi5NNtlha1vfDZk6TZHk2w4/sfOi6Up7zldX+1RZJpI
LP83wrWPlE3W47gWEL1Fa9zfS7adoSFUW/6JLOaObhrFfGq6rHiJ5RHQXFY/UnIjvD5+2tncTkGZ
gT/r3DfN8jxOfw5gx39jHitg3HlvDd4GkcoLvq1MJFHKVheHQTBuKEgKQEgrwRSmr2xR7Qznqmrm
C+9Iv7a53DvLh1Q5IupJ9FP+bOwC84dIQQQgj6J2gA649PeXGzOIHEqE2DWqcLYydYvOPYVlCRVM
nBEzqm30yWS3XTeP04OYmRyAFRf/G8MAh8/31auS0GEySGLSte3Zsgxfntj5xvu25840cfYsasbo
2XzozTsL4CvzfN156Q9Vhc9yoUzkI5hWr+ACCReN4r7aHdPl/5DD4VTjeHja3IrRLQyHFRGL05n/
+JOPqOhq+l3PHn4MO1uZDiP7rMhkO7te6HulTPq8fXkn1IndGIBAtXplXMXck+/1u4wwc9XOmLxW
WeoK4avSIvYfhJuC5/WAxLrhlAWWNKJUwvwuCtbBL7yJQ8eqP1awrvLcbWtD7bpIAN1P179flR5o
57lmvWCW6cvi4+H0v2y0uAvYLEOE4iqD4oIVryyUD8jvQ/xoJKu1POAbh3wV+sd0wHMg37bqcEX7
3CR0Yxe0XQNG/lohu5Lcslf59ZPU0yfAm/uAlsHNxjb2pZCD3Uvojf5JkvHEkJT7GCRL7KsKclxL
je1piPF5fH/R4lfOcX4PqlOPl48ksLd9ETxHMhh5juU1BLFO7GLjNLLthXN9mwmuPR3m0SsO52PR
U+5B9+Kkgps8XwWFbfwXeI3CZA4djLsaD6kBkDBzbU5R4GiPoOwNVkbji6Oefi/TWxRwEKIGLDkg
FayFaiR7rip1zSnWCS0J/YxOMzErJAZSkQTqL0PHot8cOay7Zq5KPsDeXKcvTmllncbqlxyjDqfT
SlHpWTY4H9AlGR2DufXN7ZdD5B5H39S9IIfLxABMVQFfkz7brJdnZcMnuSLAIVF9iBhta/lPdR5c
8W5hRMQtwV9gaWGycuerEYTuSVLnyFLxeA/rG3TgT09FiJWOJu9hGzDg/ZFcPcueNh4h/tPhsnTK
gN1LwsTCK4w49cnscv/srMviBQxeDDebT0DbFfJ3D+atX1HAr9SUO+NcnFxko/07pE26wLAukoa/
+liGo1X82BQKhQogazdt+D2/FdeGCMhTk3uR6xuPl4azuoamuvZemvECj4TwFVSoGsVEoxGR06Fo
w1InSVejmFzxk/1RHuBT/AmQfFk0qa3NHaV88fv2TQEND7sZikSA+BUo8oPWA3FDtbBysFg0C4bZ
wDFOHT5jxx3McFHVvCeKvTUbHn6+GVyjnIPhIn8DGgCJXDeA96+MeoMwO5DKt8+6tdMsUy6gB10b
5bl75TdaeEqjq/dmsNGCwiFqDY8RTf2jRPpEQBpZHg4R1lCpQrrO9UA65C7+xSbP5nRIbh4pqQ7S
9rVJrHy7YstpHOPIltielHrAnw8IsGygkJ5JI/XdmY+Kwd64+4AtvubVHtCQIwcBRAgw3BVJxq6Q
tadmilM50sLTokXliun+T+FQAv+TNDdowNphsTpBssguzsKyL5WqV31cQmuEuXvEcI6lJS6xn5/a
7SHyTv6LnqCKiQ54ZzxjeNyqD27P8Bpcpcmb4LG9N0uPmsuml/NnY0HYx2S3uEqyx8tTW48Lm2af
E83xxp+dLCgCs5OFw6Ae7eGUZ1SXAsge5lYYaGf/ObjQOP6fPymCR2FoUrCxXNHTjJe8ZHWp61FL
ZqEqiNSuItuNrlOrTw51s1Fah3WBETc93Eq+YnOh7cb2DaMQLO/ACqzjHWqd2t3Bsvv6H/qIGGso
ruwzjmBYnkfJc90zOMTGNhA6SkSHVpouOsU6hPdJ4mqB5LNdvvZq/e7N+R7h8Ml0DyO9NWkkzQDX
q/p5BWBUlcL9/NRIA+Sv5xjo70H7u4BLspfCOBKkxtaLSgkg6OuFb0QVRApJFbwcIfecoAMfCwNH
5CV1Ntx0IQbAOqhSv9IOekGlC9Hkn0Hl2jgXoOe+4oHVpkd+jIXJCdDLjHysjkrbK4ExXCos4nk1
W+6hKF5T/zDhNClfqN00cJ2x47147weGpsj+8n5fziiJJ/fEjiZ1bhn8NyKRQV3CVYj82Zq29XTI
UNjAyBPtya6wY7ph9GoPnQaf8aIXUHe47lRbXFVud2+wfdHaKW6lCT+Ndt12Ba0bAhiO7bKUU7DM
8PnoHCb/BcSOxEHiJdTMpXyr8JytIkI4h1yQjr6aHx/TB+3spYXCDGbRn+LKtC7vWpIY7tmQHvPT
zIBgwRjjW3vSkYqvKWuiHqOj/H8B2mNe8notL8vohG2UwFpGYtcXI+qWF5kUEBWOUoERhq9Tg+nF
BWHRyq3+BX+wItqWZh1l5PKanNkksN2IDGMdsvT27tLb43gRazfNoKkPXTdz31PiKhQv7dM85LW0
yfzmS8OJWa2L/0PmPG4akLpQ9pprSRqDlA1HlE/U88r4psGLPdiJeQhYplmMgeZesfc24dSZPSSb
JZEpjs3/uIfv7bAxkgph+u4NCD+jd4aWLsjcQiMU5wb9CSiXrR3ccLoUl9/SZ4Z5LtDtgIMpADb7
WsEJ+IC+OWU/xyS9fxYfiG0D9LOsfKyIQNwrDk9wRMTowLHjiPB602R4bkLCJ0LABWt/m9iIDomH
vniLASDcXwqBjHnXelOWhBU1lDuEDtdFMczGU+XYklFQMHFnifQTh4UQ2GUTEI/KRj2Sdz9kjATG
gtBZJgTFH7cEgHtXy7Mf7r8q8AV3aNCocP999XZa3HmQ1n3oCB6PS6x/brYDSXr/tL/vedVtOUe7
mwH8A3AJ6mdxk/Z+DM/H9Q/TDcxt0Kxvr3BU+QESSoEDY8h9aVdOk2vjiLllSLYrEdz6a3eEsy/9
gTvExf2H+SffpHvKI/34YEr/I912gRVayW1nfPHxWKvGSqXp2j1fqw1L1sF+NIPBMlK8pYzgHRsN
9PTgC1WYagEXS7RA4Wzt8l/DI9zW3SmW5E+K9GDJYmAJmtm/tKW49kQNrsY3XnZ7E40tG3sjXX72
DvRRxJ7EyY0ly4HfrsUVqcvBSSBIPk2LQWVUXyOcoigEEQXOzBottVlfig7iB0cViOZ8tBGCz1CM
M+t61a7OaXMbI9kODWxc+SSyGaqp/WpgYFlszm78oT17iEdRyY4YXfuovrKxWsvad6rvmWQhfag3
8zOSrnBeJjlSQChzGDlPvK2TZArM/Fr8gsKN3DBeD68o/v0Ps1PwNP3mDiov4I6cWnTcCvCL5lQ2
3wLURza735bZa66lx60S2nnNoXi+2b2zU1+3Nmzk0GTPkPuz2D2cQP72uV7yID+mmw1d1egasCfn
5DV3FRx40pINbt3vVSlShYNJyGxdecnCvqZ39cc3lzJrfGmwgsZzQGmUg4IZJrOXgeHFrfGWZmtn
wdT+D9fPBD9bh+EQuT3rZDArU4WifRxoJnqI99Xv/zTm1kHpD4NXmjKMfWUdbLdZl7YRG0WKA4u8
j0Z+mHhcChgTN8aP34LOMNRJ7LxKNNq+S7res4cKK1YD1HYBBFogE/Tg6515QGHtMbhSdhkzWyue
TjhOdnuVDDeu51+xNi/pg5ae6iuUd8cj/Hbknfb0Vbu/Gksdq6nsvrr8Bv+8HnKkcN5dh7JRH2Nc
l8jSAF5sx8n7mRjwouZ+3arOTPoxRx1lltfS+BOV8Oc/WnpnMKugLt7lI1q6Qc0th5c3C6oZXsFr
tcxWbDpz0BFq5il2sc4iTZq6tP7kWQMyF46s6zak0qP+mxK5v3xpICwPd4bRleDls+Uz/16IsM9x
6tWaqn2Mkz99vbxhnSSwM7e2cWUE+vyO9xHCbBZwA6C5UjQvUbrQrj1aO4Jdyzl7vhUTTYX8rVcZ
37JUdsxKSySfRF1Be5yJTg5gfkVeYR7xF39e1IL1Taus0NNBq5HPFNtpYP+zawkA2l+bJoeRCsrP
a2inCKxuBZb4JQrTwv1Fn02F9/z8y0ck9otyCUUJGN6a9qkOv/Nt2KbLwJtQ5KLHf0I8Pkxp/E1Q
0Y2ljhnpvbzTqL1Xv8IG1n8VVC9OIUAOOFdDqQHxHYR8z5VL4C0wg0YhZb2wlT6+QMw9sfum56xU
DgRXXuBKl90M4OXZXCN68/mHrdOFwcD8DpgDn7XZncp44l7CKZDhmOEeyHA3yGkqO2SWYNDvvhtj
cT/AVQUk8+0IAIujfpc6qg+rNP0WHb9HK4pK1nUVTPc6Hp9R5JPzgunYwe0SyK3HCbdIWSVG0QdD
JaIjwySgjZWU+CgjWdRoqOl/OaXCB9rIaw0OmUxU6/QII/K4JHRFrL7Xbw9PPTIdbQ6lNgfIc10G
meCz42FZFmGMzwAtSmpXtYN2tKH9X00kc8cbb7mYqdgLwUMh1uVV2JUBYj3j3FJ4w6jDWwtIv8wJ
LzbUnccZzUWwfe7oLTY0q8lMswn32GDmZxFKSlBx5ZaWgkfTSIrR1V4nCnxzvlT4N4dEaa4wOBn2
lW7WOL59gcO+s0o/uBuEGtBD9npGJDeLZvQZCsa1Wtcfm1/Xq0deh/ErODLFilwlpjX9hKYIRVAG
f2WzyjNCt1aC5wfEwPh/KNRglnECEuJidSweDIJz+3we1XjZzJJQuSVTrsfJWbN8sve56xSZc18Y
aUPRbjpPCyB9is3ZN2AF26eMRScCEcTIHkOmPGGd+rkn4RoFbZQT7tzr8B0trjVCexflMBzup07O
lZr5iiz6cQv4ZMoPlJRvqDsw5n9srJuBLuM/SE8Kgo9ub6ZT6t0jqpLQqMVykrYnAyeZ4Nc/1CLt
tHe5fvp2s1YzLfXFCLJmHnvhHGAfK0U01i6J7PAwheulMza+UNwYN2SjP+eVXIslBt7sCce+5BvP
hoXrDYW62QdyOYWu4XRk9c8toUTHoX2rxNmsBPVsyDKj17rFHRyHJ/mYn7UBZldnAy5DCTnzhJUB
SyJO66K7pjfFA1osOh1U7sy+hOqZ8Cj4TudICyxUd6sNlzAA7QMNzEVx1HcpKP5mO1V+mA44Eidc
snQ5UmueVgBdQ3TT/iOwZv6a3xWeLklgC7NwVy8/h+QGpFx/0/ENxCvBc5k5TXZxQ5eklhb+ubhp
We2Y7g04zr5E1lPOqzGIAnUmoDyTnNQ/I1Pj3VOSwxpRPQmXeIpRzsGMsGGMdkeRnGql0MCnBUYu
zxoQDiQDv8nlozz+cC3vhB2AIzISmdH6h631uTNLP+Y2ZJsgoPiiYc89ZBLD8zIM8M3XTMc/O6sX
WzUZwzMpL76lzyZ0JbMxFTkoYy2xQQGwd/RE/ydDVYsLUvGpXDK1oD39gpRx3aqYLYfNC/VYl8Ul
2bLkyo+lfHrrkqQ4TsC1kYuDk/WO2UHQ2O5JD4O0nNIJyOTf2amk/J3pfU4KNKIx6CaIsF7Pk0OP
0TBE7pmQpfVsgIrfWLp/hWQy5aATHoQQBcDSlsoaxSs6kx815WW8fwKUf5pVZMPDJw3I9ZL2rlKg
1vsXk15LNerXtRo7YNZ1/O4DuHfmWU+lY91/zojfwO0kpb0K+WpM4hsVqSXgcBO39IsVxVo8bi/B
qCotQd4DaiBKPy9fzSg/QX1p1TsG3CsyZDtcqyA6Luq0gTEzcgMd++vu4UiF7/Dg3fubV8d1d6zR
/a+rHTjg7gxQ1AIBQGYPFiKPK5KfoF89m5XoynB8tP0YrzQM93SNZxQhi5R8Tj9mYI5f5ybaSJV+
hnqfDI/VLSnjc/dvC/YLrH6woYS4P38v7W+n8cLyantpT1DWPLb4TOod9gvrlS4DvSpaMvAT8W7y
OEORB/ukKWMjlsSh2Sf2pY2iHcMoSQ+YmPO5TSNq9HX/t7tPXWU+D0f07pgmnlCRkmllDRwly3ZL
7VLKGTZ2Lc4GlTohoCEoRBy1SyerIAgjd1osRDlxZnivI25X5RY25CyUSQP7JtKW67fOVADQt/0D
Wo2FIvVG7IdSkH0Tj0bNqucV8USThYUPMWTJXKeq5/LFQNI4GddbT/vmdKPXreD5UPso/rPVVQ4L
lh3KEYseqf/4g57k+WLdQYA6b2PIiHv79qBhcn90ugNM2ol9ZnmB9FGTufCwqbktYqB8ncOEqsyR
HQz6DMtdxCLe+zJ/q+35dkedAFIpllHFxoj9+EVAMDBhq81rnxll5uJBmlNd/Este/eYZ5sDbLey
NUiDGimg6JW4hldLexAIx6uGQFinLNNcJOpGGc9G81Zaj7ZaTghjGv3TV1NxBSLvbilxzujIiriD
GHGHxKtCcaezPPQtfI+jKuy1d0oIJgF53u/ZCSSOM9jaWnq0soIpdCy6Kew9R11SbUwLcetWjzH4
U2LRBIqo+UoYiO7khNa8sZSvSUbx90yVTxZW/mr6gGMBD+he/YwERwN7FXH8s0H71SK8F7BGFOxS
pNLi0lpEOKRW8wnSE1+rM4MB2Z4HyHFAaUGbcrKPkcenOYNO8xINdcGwRts+opd9z2WaMevwIjM+
P2IwGEoEKYchJxhuL2xEdANAFexM4zOgmXZLPyIkEB3GYb7mqsGWyo+14FucBFJe1PI15VzETisf
84wN+qTzMnldcTX/ch6LMpqSPTfxfAc0HyIntExBPq7JiFTTfDKmkXeMKjAnqOK7/Zu13a3wZFL6
QBNCbHSi2UJONksbjOXcgkP7VcFmxS9ETm3ORm3V8XpsfEjyL252cCdb4hb7xn8Mlf/vWCxXNdND
m9epKRKFxXhBm9RYVVYQ+9enSFTHdMl6X1wf3iOQwIx2qmB+7dzY6sqegw6xF0vqNkOM36rpYdcz
PrycsJKsNUEODXPI99Of0Be6b6GSPwWhQkV0KENaBCDUVdRCy6rIxnLg5dFEVsdsQcOZ/mG/FVC/
Cm+/2IMnb1yWwbRHBlNoK2+rR7e86m/y1HFx+yzB4puorPeDRyO4MpnfnEpkc7m17En5/6F4IFAy
vxwpl8wpKEHotgG4MGXSwvbraEYYGdvjqY+TCHMbHgpMsoEm1KJcle42O1GGlWvtfwr/RyhPJAw1
aUfrWrFzkOgIKgxpsI+MNFJpPUBvnpdxoA417QYiInZCCLXLjEme0rdtyB85YzfFMRkg+7EDAwin
qb0EV9DMeCE9KD/e8pOt47JpBpoJ6fM9XX8H1szvOB5ByMg3HwVxO/Z+L6Cbb9qVd5f8GSfYLjqk
2LgA6lWxhCuOi4J1BlXCFbvxvNWT03pGU6fkDS1fxUppZiF23S3QBdt9zwMC2kGaQQlb5KDG+QBU
/rMhjpc3GjrljZksZKuP1svEm+hVhBnHNAONeygm1vni9qHVH/GUFedI19/zTQ4U7pyBTLFV9CIJ
XWCoh12ag+hsXLfBAxDa//4xQD6/JK1A7dRkVNRxuHcZPTuj1VkhMBOpwCiKtyfIqRPxhinF1rH3
d6f1PTqNej/IIqmpmx2n2KyU7OJ5x+f7qEEmbYSHD02YbtXj0Iwfj75gcwXpqx0UQE88qZB56UfW
NGZKhLJjGaE127bh9d6mU54FUca+v2a7yZTl89RSTnT6hYKSC/wvohER2sRbQ+fiS5C5FX8FwGwI
Ut3Cggzaq97ytPQjNcVHcXgykQ/VuGkB62XwFFFxQNBxnyTW+hkDl/wvdB1khsO1xWcZvYB5ZPsT
Uun9c5cpE5R+9xOQiWiWgrvMg0JODXWbMKlaFgu5GDMeUZUvOzhwYsunkG2L8LJ4Tcl9Eq2t9tHA
j6IsF3mruG6+BnwxDvIuZKtehAlz0cnqV/zu8MT/PUeih7FoZSsiENSV2JIuQVCvTWZIilxD2eNb
v+UcxeM9LZ61NKOHyiwaGeicdevC6x9mnEnEnFmI70D1kEuZUijxMYsKKeu2oEdpfN9CRh8qEzAj
KRlRSPPz9adqjWPKIE1neECCJ9hrUHZcrxIzcAsY0lz3FMnreFQLKBuykUYDs3iqLGNi3mq+xi1h
w8/uLJGvWYaj1oProaGwCB4kpjscnX9IMOHePcKzzJUGhHBIZN/JHhRDV3j0ocddjgszZD2KCE3T
Bx0MDjQSdOp91kM4kFcmg7C0+31z8yDS4xNYV+sb+OtIjUoHKIVQ4U6lAOCfJqjuMp5UaknRM3SG
VC+ZhVCYdJSKDuhsje5tfFHgKKvQ3e3IJkNGHCry4yUcfb7KRME6q4PTOUxU5ZVHLCX1Eh7v1pxi
GsaVZTIOExtU08kAJtoBLBb4YKuy4SD3fwRXw+6NUs98gjwNkXBx1R29NehtWvwBNc0AxgxtqVCM
vz0FrMGdSx8+XdETgr45kIwzqNhYZu5wGFSHKepF5a/WEgyC82A7y5Ucn7mNPbkOOVbPraxylMna
Yy/hAaY/1UTKvMDLddGjwB1naKSlWEhVWvJt+ZFOVblZgsPvAfy8NG8f4nx1s5L8O+s8tWMD5qMj
kNpK/VrWv+1FBPxSSTuShD1ab+xEBcF+VbSOi2p6GqJQqWKZWrRnUV1qeo4MJOuZJE5ABLRYXTYF
zpDyVDLrk14Ynhvd5Pey0k59COzBYXYvfp7CgKpeBL175AfVpNfJzaqbdPINeyvQ0KDbvAvOQR1R
hFjkpMQAGjV6EYzwGVcLWCVFh6mIKPiEwaLZ2EYcBD3QSXWRNFBDzgwgbEPLS86k/ZISaIOZ0th8
SPtSK/I8Jv83/ispMFx34VR4cYCGJXWfElgG4n2AkWNUc+CJS3aTw2ux774UYcDLsodSsEihJjU9
6MCBZ1cXtPFts6jjl43xwEJ9woxT5/YbzuMb/IZ62cnocZs165atIR0mG588sK1lg5cz0RaJYkdV
btsF7pqAw9aPOx+HtEnBjqgKR47F8nrYVHI5Ch9PEsrMZWotpYl2O0ITHD7QTN+NAqZsgKDRlc40
ckRdAz6sypEOXzYA9nYV5d9WaViQy+Tt9Qd+hglFA85UcWOzStGSap2fFrV0F0L5SK222n+gEkHD
eMWV+m+6ophhBX1eFIQ52xGB6N2HCyV1blHm71JOx8KIyUTLGc81BLFbSJqzWMdx1JtPFCDL4zIJ
iFc2TPKWtFTlptpQDV6ndBQ5s56RPlE72Nya9XGMHVGgErsdojfeapBBzn79jGsEVJ7SKjR3DG4/
FBMYYdZ1vFm13tkf7rEHbSpoxmaxezwIY18JClwVgYmQsDjgILYXL9N8ejX2ArSojEy6fQl/VMPg
W3Q89i6eLa1xKPCNZ4bi4cNvHEKALiKynUQTa+HaihdYvEFRyawBLrPcsMv9pZTldq3sRFQTw3KZ
4crVXjZaPnBv4DbWcucGr1SKfGovwkWsAQdJzp4L41qaOv2AhFrAA7CngedoQ57kpgok8LM5ZrYP
kW4rcu+bG1d5OGL3fMQ1FWMN8kgBCjarQCEr1h/Hi38gYspYewzv2tZyHlwm/YUivwS2+I7uY+wE
7vOMsFKxZS/TKc0QLXKhpYn4ZDIgh3Aqhb3R4SHClzNgJ207xen+nX6LcrIkmWVtOFxMK0zERfUM
OuPB7u3wn0AlIIG5OjTfTlZviORSuye1OLNTvxCgLv6LYYc+LPHSeYyMYnweNj2jzGLhaE4butzE
z4u59xHpH0BQ9aQQh2a5OBXqUWrxFNc4WHh4kTIN+FMNR/IWmbzNYrCLbF1EqJ6pSr++CZ3PipFc
DAhRmz2kloiTkhjKfDRsCaGN6hH2JsKXctYLFq02XQ/fe7Aja7MuyyD5e3p5C98JAhjZVSh/mLbH
LuSX493fBH8I2PcTNMkDNWqQF8ZDLu8gsnThDyiq/R/g1ZpqMKEVyYz7ofVQG0A13cHn7+tuEvTv
E3xyrBi1d14oSGGNbbTf/96Z0ZMs0DQhLrvop4faVoeWzxc1Fs0HLEc9K7L0CIQjWvhZSbY6/41L
JBKY83Md2vIvUKMWByDB6K6F4NVU2AqRMzrve2iR8g8JPdJBlRMPETRxCJoxt3+5fdUzZv69zviY
OROrUvrC66WqBUbKGifUEj811MbXupInBQ+XyiQXGXUSmd4BiFBsZAwF/rZcLO7GMAiP/CO38u5k
dSrOcxxU9XYi5XDrAH1p0cALGD2qVKETpmH9BYzCLwcv4rRjA173g1rOHYgPZnD/FBIXhszpIotF
yEC14LiQUMQLeoDBRqwYnBOZETUl9wNaq7b9dERrqyZyjAswHLbYeNxbxdy2rBqqtgfJmQtXozJH
vqaD8o8e5IrUt72yyex60FbeKvaqfioX+ex5XE66Det2u7eo3jdoSfJ5ixhpttA+DRTzHakpZPUs
Dp7WEXG/5AfQ5eEajjtR3ZMrru8N2wdbG54UV9MxbJe4Bu/WaoMSaqJ5o0PiXKBcbO+CR8cKte9V
dZT4DMq4MnH3ShySPHFiMLI26jcJ0tdCXuhx1ixok6XdBFBskepfUVxVC37CifGv23stbRNBSdVi
rzQuF++38agTvmeogvJPGX0t7bGH1LUg+4j2sardoL5Qoq+CVqg7Z55vvmd3eyJUrdfZ30AGkvbU
SHdhGDbDkc5vw3Xve+KiKKF6RogmpLafmoJvCg5qLpCfi1zgeVP/83Jb7cjbb2eCVlFpZ5EHPnzx
NuqbWbfJcuwkgWxzTIu/iwDvQxLEDQl7MWK0PVdcXohl0xk9ieBTL154dtB2oNDaascBELPh/bsi
kbpWr09F4AvLEGalY1Tj25gbNfq7ZvQ0wqj/u4ZMF5ZIuout4cJKdOCjiOr8Celax4SJyWEtdx3V
Vp76r56mG9Ub9MBAOQzeCUyD8KGh+Dirron/YNgye3DjOzATlpD7YROdU9ftoXZccpXp4sU7QvAj
hWRGvo+BIZkwWUKIXuSf2g55EygekCokjVx8WAcFjezL1rNgJkQ+ikuYNrxJLlizCnJAyFFQ3UlL
cAIDPPB2YULKLkI8M5nV7L/VawRyRykxqft7YajmZsIrt7/5Ib3HzsH0Bqr8TXigFAtmfz+wiNY2
1B/piXUw+Vof0XPjnC1ylWN1pGxTVIFjfa5LvwRxtjiLCl3Q4+8CSszgoRjilKaJC/NeToKi7GmV
r1vapXoKH5ZOb7u0bs4I8k65Z7W4qWdm5lCakLf8oz3Lov/h/qegS9Zxzc6Q26UTNTgpx84/xEmi
eODxcbvzKiINs+QNF+Nz+I3vI1QDSMxjXQKkX42/Qd4D/rHZafI1dDyI70wJyXhsf8qG1vrKNmUw
MrrBO5ruRkkaln6t2XOMpmQ0fU7sAMLEj3b+FxXyUiteQkrtNe/c9nfQiOtnhyEHflhUsgHPqwpU
hjjQNsEVkTQuUfCwiRRKUR4k/dVMf16/HpFT72zgXep6AF3xPlqCWXb8fJtO3tYh8NiQmc6Dh3J/
A2uqhq310d36EIW6DXOVjcI029LhozdDBneqH3RQl7JaXb+YUvzAwSf+kET33Of0lNbO1xq9kBwt
PxkNlH135aXGWrPrb4HDTIgfzaeXmQ3i6OQ0K4nsdBxsSllhipyG/5u9Zr1W307PEDnX9Gt+vVg/
kzMoTzFv1ajux4qy6k/b6vJ1faE7hEFa6s1gLJdBMVyO3/NhQAE6qR5adk27vRYCkdNFvyPln4Mw
htM2Em4TX4Axj6elvdY56Q54AXBDXw//e7Ob5PShtgbAGpKSvG3bM6Qbtep1CnY42dEgofv45OcZ
7PSn5tQ0T4Ox5VA2E/Z07NW2uvG4LIg3YUrcd0xmO8TyfecRn0QE+elPTcWcl+RLkic/v8js7d2c
K5p3X8D+Srih5+4wvXrauI+S8IiZvzUnvinBeWLSTKh93dzcBB4fCwZTCsbc6szZ9dhy0B9idorn
8wjHNpfcJ0j9b2otXk/pbixTAUOLIobYUU1lqlZoVE9Bj44mbfxkEfA2FeWR2gNobHKeox2NsapS
e6Ba8GwqjQHCjqcvNhY1LJ6sM1qRUJx5uIpKIulIwBTaKVy3ZKNGfS8M8OD2ifPxMlx10qMbbWGb
NiVw2d+TBx0ylF+nDT1GvCiTjVi6qJjG50T6icboQYv3LuefY99mocJxF7HY9jOPllhuNa7OTiQa
ivCMG3w/yMoGEyXPBWcFWas7mTENoyKDra3oj8tKuvmWD1IA0zuFKG5CDXP2Z/CCjNum2kFfcFNd
e/WqK3STQmrhMIIwomMQFxsuEdRlvj05VJoy4v9hDwzDPSs9EO4n+CAXa6g7Vl83AD/xAINLwbdx
g4t5QrYNArFFmEp641DK8jlDKLH17IEh/Sv+N9hundEuVKm7eVFvJGCQNYequGdJlZ5n+i6w1sNw
JMR2gdNYiOTtfjV1+/zJRmXHIFzmhfCdGaWqxm8DXrCNBu4MKMGe3tAR/CFUWN0Cy4/gmZul+KSl
hp9aGpsx9/xfF4f7ySVfvfMFoC3SF93J4a0biGFCt2h8bRPgQOr2y+S7Es/6iOELpbyQQ8hphUCp
6jOW/9B4pJ1f32KUSxewu/v1AOKpT48lgmggTYw8bnHGobCW2/rbf7liEL2fQA+MgwHJub4yvDB2
MOJJFFiirZaoio0+//huy4EKZbmuAEw+ggLSm2BtlXVLiQQO/lGPFli77xZWiC6AqvB3qnSZmraK
uPeDfikluEDIMrCdi4UE5IXXVo3dtWZlccMbMcILnQlGy1+aM6Lk2Emir6KBYqeZMIy47c9S6yYe
OTsYbIW6oVC+AFfh9TjkBbmyltpaJp/xEqwCOw/+GD2WVFPX0YzAgHqxSlx3ZMOnoCymMrixz1PR
tBINXKC/j6j+F5BVWqIetUkRqqx9K1JqsuKiWnLJiV/Xkn3DdbSOecsBHZq4Sox0vxslPPIxL314
hBj4qA6+RtNlc9d3gSDhaKO538YV39UZfnWQHQ3O9os/gHuoSBOUq9MLFi3/Rh1z/ho1a+CqbyOU
nm1kfyAccsMf/2egCCm3W7zPj+ra5F9vfWXBsAE/2u0jYpWssKx/p69awJL96gSWZE9pOtnD8Dcz
fo0x4epSrAa0G86IQp4Rj04Gr8yBk6ChFjs7eoIYpY+HQkp4vKWjxe/95XlawXwRPr+6ds3xiDQy
Roi8OwqHxJIiCEUs2j4Fd2alAe12AR3Va+zEwfcQC/iFq2k6/LvLSHg7zuPMNZsXhshnsfqv+2Mw
pHZq7kZ0krRaoqBengROhDRZ7AAmW+oiGDbW+1UDx5WtKlU9cUAmTzKet6oPgoZUrMrtLjIcbrd0
pQTT2HJJ+37ulEeQ+bG1LtZySYO4mn/HxjbU666q7xJOThQockkQufI68jgX4V6xHBwyOnnPxBK6
UGm3z1JHmRI4GjyhPniRkZ2gshUKl7lHuYVJaCiOY2Lv2nkZI5LoXH5Adw9UkUakBn7fREXpGMvg
W7rmzGyCPu9mThSgsA2FXkyUw+xK3I3E5n3/0lNjcqkYComYCa2ZfxSovLprlj3N7FBADQGR4Xod
z7Bu+WRLCWjfTyRBVeXKjNrXk2FTOlVnCq69JvNg6ZYNsPwODXZkpwf21YKtq0x3u7Cz2ylGmE1+
gZanQ2GjBRE39/WSpGHv4O6JUpEikWTMPcdk1lJyWF5XSaeywq7sul+OHmYK/7iCq4oGmbzvHp6F
foe2KkGm9Ft5Dpvzxv17TZqNlpPwE3YMMg1j2JAVGHM4Ia7tylFcUg+3bbR7P0XnN8lJ7LWGgmzk
xe9ZawhCbjE6i+THLbTDCmRlTkoNacC339dwnNpvdHjOjpM8gYx10oKdpwHMSeO8k38SfzlYRuK7
Iwy2tT0hkvs4fhuuuTHk96L6gpJy3YMnMVWiPg3kNT1EuDdUHw6Ylo4LKEacTLCbdywhRMxwts+Q
+9V0XhVe+1w1sqR0iNDm7wJf77tTnBbBQ6kmtVrDEggAqj3p9kfFR0hVhHGNh0h35pFqGifjaRgi
sGehkFOTqhoN9OLo19qnN/vzgaDnm63VFSLu7oJpr7zojZo0yU8CIHfxeYE1CN0u7qL60/pZLTa3
l2DG3MM0Wtf7wcdQ0YnhtzldT/YlyFLdQ02Yz4n1Uk0UsMKcSPXhw7/Ui4lmz+VhxuKnrRDeDRy3
5pK2COlfa0qDvvCxreD9oU/QRxJOoVu2s/q8nlBG1+NUPUAVTFUTHQAICaF3dgp8DeDE5GBIPnVZ
AuDqEJyl/FHjj/bXukUW+hW56alEzBqByEJhr1RpARLQvQiMuoaK7aCsUpHti9mHYJPh7ZCoD4HO
/uzPwPTUue5iMLPnlCCMPbRqZtF5PyW8XPmkpJVaD35TDTvxRddEKF4rnKcnYMfbBcUYFMQd/2t+
1p0sMAPYbgWRvhAAKe2Rn13AIaJITE8ZF6fWabFJy3j77CfFRhq8Z5J8nxI5Gq6l821sxzOx6/og
Tr0ZuZ9woIYMsNCClcNOjxuNGnAHr/N3XRGauZ5VaCUMR/VaDZG4MrM9Czyup0aIfj7HgstCfHQB
VZgdDF/K/KGNBRbudFUbez0dvDNvj9HUPCWG8hICL5Och6YOS7Eg6CFZg4mVllohzj+c+vnss8pf
ziBbkOkct9h5HkB7Xi3Bqqaz2LsKJKNo2CR823wQ34mCgV7lpeqghEP3r/Pk9xeZRdZ61RxPqxvf
2JtlFRfMBVUHGNnhRkDBvVlL22BjC+PBoxjLuGd8hsbTBM0qMaZlFZKdp4QLSFrSxTGCSF1LyVfm
8RsV4tSws30iIuT6NOhqm4bYXby+iwTLjY+YbuZzlF2It3Z33bafGinBYyf1wt5erIu9SAArO9X2
AenDfGWimR2fnzlVel6SzOo6iUGQTwjUk4I9ay2WifeItfhh55/KDFtkmG3p5q631ZF/w1OHRVWr
xmnpEDNk9e/9RoFgE7tRDt24o+kqh0G0RJ2hrGa49AWAlzl1QK6LFCDY2RA3bZ0tvbKW2xAZf4Gw
Rld9p2zSTEf19rDOjnbO+HrW25xggYnBYosZl4nm5+ba6V3CL1QF0/kI212T3h7+Ic/AS00LeXcd
Aox+DS6ZJWwEnKfmDXSsA4G0DuyOY79sRRZr3zysx/K4BmN+Mt3kiKAiXcHVO00oaQPj4xNYHNfH
5uhTbri5HFFIIp1k30OIaHAl1Hs+lbf4hXsP33llL1DqryF5gHxUMLKXo0l2CCXJwFU7qBgvIfB5
XHYHbfiR/dlOBRzc6eU2gakTzuImrfyqTfim8gSX7ysIjUvkmYYvDjiwXU2HYjsIQg0NMB2lRleX
zUzmdd2do11WHFzrTCTugEbvRbijAMNSSWxkW3ENYSrSjjh9hgqJ7W7LmkaeC7Dzhn9oiinkJLwT
fEjST94iXiL4ttxn8Cq8qYrAFoM2xzfxqdbxEXjvhE9r+J7m6ME9Lb5hRCPm8ZJvKDojqEnV/wg/
Oe1c29Mr0WJBCf7VMDbHUt0BAalhEdKY1AJlu3yWqjqorW5kB82Negg9UOqivBtCkrJPrNXyqe99
BFX2MvGn6JNH1voN35FNvbB0jHNaFLv24fkm9Jh7x6gbfwYnWBPeQgJUEAjYkaJL862OUK5m4yhq
qt+zH6/2LJ70rQ8DV7oEiz6YrnzJOz4wUmbIb/Py/NvhfH1LBDp9rqWnYLN05SFmpfX4cG2MU6n8
IEf4imxMiQtYuDzvZW/5Pwb/tlDRdzuxBUklKFtkumGAEGgVchbUthp8fbKp/MAOSTQdwigVOkm+
KHeg4Y0S5K7pEMuOpHeBKnLGrCyL6lCAdRvaqWrgySIolmCgt8nbq38KsLrqogjC5K60ii/fIhXR
Ct+nSH+Ks4tNGQgnFeGu/AaBLbuzwaBw6A6FX6zC37m+jd68SFcurrU75mtG6Y0AFoDdan19ycsT
rMvY3THuPaBRMYqfwDY3H/KYo9a+8+e1wEw+V6oWKIp45o7N7RBSLUIWQZp8bDI6f5IlEufBO3un
M1r2J8CHH8nufimOdOzbmhH/C7UXLrhNZ7Oc3VXYKkfY7bdLEcSh+UOUGmZIL0BFVg+779kMy9rp
BMimPlY5fl1nYbyM+ew8+Tr+YSCr4WcPc+eUB4kQsMay2d/k5KcTPcZMbtoKCxX6LBPEsmqo3mWK
gWkqXBd1GmaAWPQRxoY7dgCt8qdVsQmvbj/v1e0EiiMopDpmpaXtbS7Rh4D7rxdLeLrtFlLZLVHv
Bf6MUbKs7hMW4IjBouzLKFON+32qPDVOpJ5wCNMSo6wK0qA1Vk7G8fB7Om5l+HvmPFvzSXD7EfRv
zl5d0u7N6XZMHmj3DrpPomfaVQhLb7NVHupMoaLxur4fy50mYEUmtKH4vKLoWHSMoJyDcUTP/WKm
exHWGykddim5v6NMdeRYqEaEIRtnfV1KhYFaUUv8b3edHOZaz4+ZqU6jo8/lUOiEnkT+LArnq8fG
+UIIDtYTj0SiUdPpNWHoZ/Deuf70eZgt7RH082nPSEJaLh06dA8pn4c1nYweJzikqhKWVzPZSv5s
fxCxN1Uc34Gds9vfs66ZVgK5Rv8YHHo40fs3DrHWj1OSsfFjghqAccAi6s74Q/uuWTp8llLDyE2k
D5A5CFMqDbsJmr9TqON9FCzz/YRRy+rYkPgpQyi7O6aftE2iwCICU59i1ouhsSDimRO+IsnA2xqs
nN0/f5XQiBRZ31f2fB+cD1eUw0RG0YkdnMx/UD7i4pp+jhcluPpzE4uw6XujHCknsunc8WgBoSyD
yHMPNzZBx6wfcVTpNw9ric53814raW/o6nlvvAuQLMHdoXwBdG6PDqo+RRd1b+0JxIbZ3qh9PAcL
rzzF89J5qIy4ZlI9y6D8/8rI84sin0qbm+MaNM1dsPv+rq1iegsPDn/U5bBCFCtbwoydoy4i50jK
CLztVPj4qe8Eqfz9d73UVLI5BLnaYoEwyM9Ukhhq7ECEnPA9YNTznArrqYArDCtXJOYYxlKDr0J4
AydGFfx8/6folhJjVFY+MvQngMp7r6bYLVMpkX3HiOnCqIWRoTRjMOgqTHYrB1KEITucqljYIAMr
16ImTmxqOJB3nw6l5EJXDwVHOed0T7gBJplxKDbBGZbG85yyVoXs6ZVIKIOzrXmLH8pQFN6Zz/Hq
Yt2GXp8HvX6G4UG4kUumHyk7mPUvgDUaU4cl95Tuwz5etc2QtJok+Elf1p0FvIKkfdsY15lAjDUr
/b9D+cPl2AiX0LwY48U8XRvjj4CCtj1fGKFM2Hiq6dDHqNCu72R0HE+s3SxXxFKXwxNoyG3JU9Xh
nAA7CqBRoQD0Dkmz2e6RS07R1TQ+wGkRhraVH0+61wjGwsHx6gJQBCPz0MEy8juZRPmb1dmTosph
ZxQ1THi3YsULge9ghb9gzNhIg0OP7ohmis35ex9LW7Sf/5/IMmuwBMerjuyGx4k2gGo7yd0ADXXK
eEqM8ubHy7Pzc0ri1VrW5pEAO/WG/heA/WUIy/cC2nPe78HxV4Vz/dg+WyX49jvg5s2IHZfaZmBF
agBnrRWU4397T24eHMFgod56rmpv2IfGsEir1he6ESaGb6Bs8rNMMh0AvNcTsOrc2osOCiapPjTR
RapaP6OvGRpC/AIvRMMRJTn7UKGBNYSIMraFslQ1hrrNElIFQOf/KF6r2JQrsjA7tfaXHBpfVJAA
9nH1708VhbG0xtJixIPPDMgmEpXB9bww2DvpAfFCYkjCqrT9POng9Hfep9ktAPCxEXLtJELNUD98
6rhDoBy1XBLiUkNv+7Hzy5ccUwFOBAgS99RvpPXVp5xs+gs/BovgcErFFcNdtqoxNsJFg7MllNkE
HhdbcHvvaXhc7LUtbBic8SjfA8e/7wLxIitOTMbhdtQuWLfIGZV1d8UU03jYcrtd9EDwPKTvXMqu
D69DpMdC/mhXVepZriB/hW5Pw65N0inUHitdo56jQ2lkW1Sc2yHZo8JAFURzVQ1ugoxewV4fG9KH
JQZRPLK50haFQRZPQ5EW09mZvut5B/CdiydUx1i4CN2VbjqUqmKEvj3g4ieO+h9SpnfPiwgNLLOc
mAICKb0uybS7xTu5t19U3No8wfF1m5eFmeDCquUgudYYtd595RkS526jSyZl9w5Z4wo1QrmW8Q7u
JKM0LvoImS4YA6aT95ud+pKPr8mhvdBzaP0AYoPmDj9X8iRaZCMgl3gpHZjk7IDnXTzyYw6kZN2I
BNqEy9g8YzqG/k2gmbZFcX6XEqRXJGp3YrdjPLi5cfwGDyeAHzXLHzJKlcw0+1Dm0JpAHnRLCLVf
Whq40FwJQBAVD3Pf3abedBQsPcE/o3qq3/DFdHhpp0fDoX4cWIaj3CFMHak6//Qa17EFki0gemLY
R67xKCdUewVgu4LVdZg8VmWd9kQYTCE0+f+llR0FToLvzVL9NQALLmR+5r6ocGebfnYwZn7wTeM9
nrFU1H8nkjClmVWMNiw6op7vSTP4hjPfHQdIwg97RxBAqrRW0NdN7wLdWMY9N4YSFkxpUWgHxaO9
jFPPR8pKGiTCYKM37zFwE0fOTIbn8c8Sa0u3zwvmbB5GImCssOChcCB6/uE0ueodUGyrfU8+6OCL
2bhbOA3SRVUKeEVPUzYIeqomwCay2UcA/KULoIB90b/pUqJZbMXOZd4JdGL/M7lQhhRwmWqHB+ZN
3uocFTjVvQBMojgckef8ti9PmmUGYn5C3lU0mWu6p+bOyoiqlu6yOegvjC//Md8wWfWLiGunkTXr
q/it2Xyga37AUCCyxvk7rJ+TSORd5X5SkvHlUvDAq2DAAzuCb1XmKtYCJ+Z7D5FRV3A2odsYDAEW
ayqGQL60yAsSRyHxDnPzbkWFLKM9dmXHBSIxO/iv05ChUD0EfN/1rmYu5G0Pn443FekHs8qxHnbx
mak0h1cmJ5Px98Xgh9zMg43oTI7+OsBy7PxoOXaQGLimUtz9V7e119JTPHrsd/e2YxEn97CgCHKO
ogW5kzcV2T9t6G4YqJ4ht/jaEsZWxDr0SFYx0Ch90p7jtTxh3wQX2/D824GtgkOCn+n+eB6WuaD8
4AzGcQ2ilavXJIfFp9jcR4rHfOlX1oVm8x2/zcfKFW6a6h8nzmAD3L34u3quU6xtIw1bEKg7JYbW
Uj4s63ZDLyvcVJ8l971IS8vfhnRdWrSwEkOIHFECpPJbkLCBrUcdVRiskpWVV9T1AQoUQNgSpuHw
CboEQmp2oHX5/PEJZu+cQ1oZK7CiAkHHhNh/G57dtqulxStvCZgMb9KfrhRaJSXbu6QqW86FP1Yk
0LtzcVqwYkncHOazS471Zb/HSe4kL6PSrKOKaCJEzlYi7iNQKQZA45rzCX02pduo35ItVAxcWmjc
w76SjgMMJeO8oW9uncYDArLH8mT6E/AyrLw2TaQmRmR01wd4BSg8x/Ur/LxIaqQXpyXgbEB8s2PW
7svVzn9citqIcAuIocYx6HAreeSanwz0ABQVGmnLmDWCPN7SLU5W7GRswYeVlTd8ix68/vIKSZrp
rIjZFZUwqJBZFhGVBDvCq7wRGd7OBoG9Tjqit+M/r4fAxQClR4GXWDeH0tMtK5PFLVKTbafd5aja
pYpvaapucihXXGRo3q/f4AVf3ASXqxHoGJYIoUdLhddBfe6uCskxEVqnO1S15WWfLbVnXaScaHIo
1DKbAwRoMxaJ5lOJu5ZbZLFpU28K8P3KfV4YEFKTi4mf5REBQfq8QaQZceaL6ppfLXbeUrQC1mdr
I/8qHTAMhpdgPflmEQwRZMIax5bwUbanEHt1fgW5AF6sSDb3v7rBZthJCZT/ivPGSvqHLSvDiRiU
BzkVe9CXM8wyZmV0Iod5akHaD7wuUX8mFc2tgRIznBKQHAL7Iow1f8ce9jVNJMmgqyWZ1klUEFkt
B4nTs7kXOIvK8osEP7908RWmLc1D9doxH/Tiq1zGKEjwk17zuZc2JXKxD1CVZzjG+avMlkB3tRzA
lOtFRAouDEgDqq1DxROpD78hygAy1yvMr6oBu9X9IuGmWKSrUxGsstpxCKEuhNVI7sNNO5w/l2PY
PVmu0SUUHLBPbHzlfFSuut9qq1NMGdyC4Sdyq6E25yUJLUOlgEZIXxjJfDbKn26SC9G1G62oOJ/8
enOih7NKr6gSB5VPR7zsJyAUWSBvsxnVUynrQNrLCGNF1VCnf5NeNLcT6tu3H11nmv8ji7fKfygJ
R0hnpyrw1zpHDdUip6L2sjqjo1ggVjiw+prxysT6RmEbpTGcf2LzKcFJEXm0iS0xkim8XLIgBR5T
MVxJBTsIWP8irwybYo6/625SZfLauxebArH0kH4YxP3UL34A2/1Zx9hNdtB6r/vnqdBOI2Z1s38b
BMaa8os8TvX11faglPs+83sq8nprBZD8puwEc7l46XVF6NHzQF/EA1595W0umyPok4XhEItRzA3Z
aIIFOGfQZArLqyU2+T4Q3cmS0G2Kg3s0zz1JX+cMlsM1I/c6dNm+KPbogxqLSP4pfCG/r4ckI59c
2GBXgpxCZPgQk05CbvySORZUJpbQMpeH73YhxM4Hra8n3BD4QTy4Xjz72JeGPkoBrwcfMRrgTh/T
s4dRZPNsNVa1ed8mn+hHS7KcFHxyF95jwHkr/aB6dpyVuJnS6klKylH0xRG01QElivh5NvtvQq8Z
Hzkz3XZip6iV3KMYQkH4Ir1hnkCTQztjqcN3f7BytEHipQqq1m3jmql2bjZ4r4rsOpKn2QIX9x1M
Y6I2y/YikaXCsvwKQbrOdKDEo/V37tN0adcJ7nIFA7uKN5/OTBoz9TiuxVbRTfnm+wnO9vWK7Byr
gBuUD6cRT4JnaUkSoBgRWB0nVkqgSNRxqT3zvcVzhQ08q5N2QNBhzGKvzE/jGJaL8QY6vS+04t/7
/6QqHgL4SIsIsAi6ynOQDEQit/f6kE6OtaGG7tAKDTaqaCA6PGjRUTQzSWCWv4S6hmisgiI4TsPj
agwnak1jkT8l6ZXDT0qRDkGHnPWoeb8F7UJT0Pv3iqTgl4ES5UcEyTCaLvag8r4Rve2qfCcTXAi/
33y2gFBdYTYartXzRsJO5Nwo8peWX+G+iiW56gS0TdZatjoo4mzHGxO1IyRhG5eD8eXtfADvPxCq
vX3IKhRtL2VOepEsTfyjwDJmwCsV0WzhD+5QXcNXRZoLgAKPV6Mxd9uX58vDmhKyxRIuqkJhniNA
Cc5DDFhxtdVQfItOPgiGkYg/tSsuPggjIVOwyiypPzBzDO2fda19Vwd29gXDQwZ55sQgtu2YiJnn
IbeyuaFm7jzd5Yoq570fGQwOAb7roQlgxki26/xSpKjRVRyzVVnwytn1PQWuVS8fqAGTCevadJMA
iudN8Z7aA4/5CX0rj8O+GUQq6582yXgg6lXTMixLor1tlilTrB9mMFdJXMDh6znbFF2GkQSC0tiK
Um0BJcySuRyAN0iAhyjS12fkEKMjq8CQWaRLPZL2GpqOBSk7n2y/ru31Wf9QdTTqjQFE7n9BIMDb
zOy2+4170lQnsDZ4JX5SB8UJrENavvTaymNkIdC6DT8hPTnNqWBatCIZEtSiSGG3dTr3wF/jfSst
tMnVtJukLFJylYut/Mhs4YAkr7+AYb0wZD1/JR23kZuwO67wmse8dcw+QhBMxLaXYd2Cva9L7T1U
d8xh7YM/zkhQIBtgr+hwUS4QuV3Hx2sp3ffgmpFogTbZQIZ5Best7+jvVfCeu1jE/jUIieogSQfF
tFB07z0X9AZ3wu+8BGeNzz2CokRljr+tfBSXKvvjsLQ+dHPhepHEVk4J1F6u2JwDyneJwNLBn/9B
D+dYSAYh7hbVY1vnsIkHYJCha/hdQLquSUh4fO8xSsT3vIN2rWQ6vExD0MFXVuqWzuC3j5qyN2wf
zBhi3GuF5Lof+O4odrhAEh21TndlZJqod+zV/VH1FuGozEQIcE19dJQSRQBy80YfUw2jdqfZ7oT3
4Xkyg+RibnSZ1pf0r4+yVS2lohOjyiz9yZHARSHoxKfuKTuWIL0zjI06t/l7sY3PIfUepNB14EF9
mJ/Bicrl4Vb+3/uI85Ijv2AnA6CRU+VG3RpxIuQ7Rbcr7ysSmUJmfYH9+bkIzlhC1x6uWPL3dKuV
AgMFrCljuDgxW/D5w9zAm7z8MMjRZY+GFXgmV/SIYKp8KfAQbL3ERPQk9WG6e4jYLudgg8U7s+m3
kSMWk4xZmzgHxtMYf0R/e11C3NXoMeX4KaWJHP5QNEf/Qf2CLZb86ciz3nBOD+EkwEpUeR6rxIQ6
28QmctuQrbe5tJeT+zEgaeCcmJ6hKydIjnFTf1gerW3bSvSDzdgxqo024DA37SuDvntFOMAHUU9S
eWpYE/fnBcLtbXBdKdoqVmyl+7qIRSorR4Y2vbw05voYBoeV53gFr3kaA0c2jgCNlrPD6Rf37o7c
DFmaGTbhgcKPoWvI8kGxCx73uJW/hfFJdisBq7ghBI7Zjfz96ZEAtNwPJCuY51csruefGga4G5Is
0xgMkbBIvcyg/hIlWBBqjwEuC2Srq7rDBXQFStF/lnNg5VvwJaoK5DAQ3CM2mrM2BIn2wSWCqZKc
93Kri8OU59LIJTHWK7JM2WLICJgnJagWl5533Eep4NWfZZzfCVL70GzYOX4OwAtoqtTSNIqknoP2
Yt1J7CxE9/Jw0vyjMfaW/Da7NeIy7zQ39lbwnW8xX7v0mL25FiJGOQBjMiZNbWPQsRKPNfZC/eWH
NATDaYKpC+h1oVFG3/3GvBd1uWlYZ0nf/0ZUhIdXJv6tV2p2mEaq4mSILKxCXt8A4tDiPf+q5kBE
A/kxfza2I6yDMD92DfHAewf5/2NDOplvwNjs+f0AX4BWsGnUX+Eiui1Nv7pYPie8Yf4c3EVWUO4y
vWL+pn4YlDZVlfmTYpZ1qmxJQw1d7frwRjkM0xYOKoySDnBYLU2Vyt7HblAf2Ut1UYuuMOoDaCst
r8hEjmuslis1rbyinieA5M2eMp5xejcukL3ooimJ+wwVAUBrZTa1PUdJAO0slBNNBg21f96n1B9P
+gyyBhQJqJmQW8vc1QhycI9TIGpxzyMicBxlB17uHa7eeDgnSt86orH/IrENbf+tA7VqWFZzbR9J
QWilm+5MIFKAtU17uDAyy/pOMaEuWQ+X77kdJboIxLtOaoQ1EqQHFem4qSQ+P+8Fz5Mh92I/C+aD
SOg2GtrWznq/EkGA0Mzr9LppmCz9i8bdGT8fqudxs3CPRo9vIEkm5mrT8HKkACD13w0lEP30jzyY
jNP+VBOVKHxutt1qyCarnjXhJ4S3/ZU+tQUCfNDgyqi2FWwwWdMiO4go/7tToHWP51BSAWgUjflK
Ehj0BT3L3iRqfQT/wFHAcCola7RiShUc6w9RQpul46X6ES2WNwJPMIxkSRG81Yzi+hZ13k2+oRfl
HO49P0DGbrQPEgSH19PI+NDmchpRKfw39odgW0YSdlDC6aNqjX/3dJT5kDIzxuEYB1WpJc5WY3es
t5uza3E0yj4RoWm3oiEox73KXTpIiythHhaReNxTlqCZU7LdP5NYdVPmbpuYAhsUU8uTMJB5z0Lg
6IJTBNDS5k78Soqnblw0bkkkn3D2gpx9LV89pKr8Y99PLvQiJj8JxAjkttSXcHYcjtN6/bC4VqXu
bxd/UWuPAD6mMHRepu1oY3DR3dVbKIfuap2ukmWEjhhERmOLPrxyiRuYVrw7WcbxMdItMfosGacF
1uZwv1cAGhpIMx9KmAtuCUt3oMR5CQudML2Wvjl9Jkwk4/EjgUTEsd9xbl73NDoGMLOuU3t1S0Ce
cvQY3YnoA1EDUoH+YxkrWDHRBf56+xCjFU01SRqzsOVy9jqvQ9M8SAYPP5BRWUz7y+x6lTE2HZxV
7C/VkTlhbxRgbQjS0UhZ0iENctopgfz67jAjCYKtwWEW8DN8kDGyjtJkw5GVNEZdN/6lOfL3+iR2
OR1PxtBNBfaBjjlIKH+udYz3WWZ0KWwmyfnpbgJ+yggx9hxsYJ2e3XhJidJLRhb6drf4j7DsFGYQ
QJ4rqKRWM/h5RA2NSFAqoporjtHAORUSsUp6xUOOF1qbiKvIiXva1h10RYrsbnVJuaGPRPiDr2LK
vBzXRbmskHn4AVsrdU0n0RW80Bwb4H+HsZ5XfQmwsVljlbD5ZD9qkuNTj4lnVM3wxQ/9rOERThFZ
MuDJSuprwzcRl+LQJUxh4PuJvzUX/C2j91FA30bSlOfV5pDX++IanZBatFdwjkDVRt7NSO//FZPL
ak6dfAc6O3RfFxUqezJPTZln8GX2sZ3LQ/utt8LukdzcewTaDNxk7JGZdyyARLh5y1gKHQ/H+gFB
LuITmeFtjEBF1qRf8ewKdmMUVgjlFiqQLPmvMY9tYDuVaUAmKqQHNzEe+tGLJk7WUJLArnfQxA+h
HgC1OBYfsiX4nAoVlIYxQteSqp4YaYSynJUF3jG0cboDPPw3+iiiuRccaez8EbeMWd910JnDTcT6
v9qd2SfJBnCwPLH1cnzX0iOQkqyXatojwlrltB3TlDkeozcONiGD+jnADfxzDIRxYU+au7fuMn6M
eDvfRoGlmSrXzUYdQApfUmsMGOhyzL882LfDoas4ezFIWbQx+l5++s6lHXaV2yvybbjveL2r0qbw
tl9IgKTKtXtYD2FVSv7fZ+JBrlCP6z6+8VayWECBcFVrnj2ne4Vj3/FZLVAMN7IJTOR1i8se1K5z
lq7knnY5xFBEAFqdSXwdBDtjt2K0Ssjz6tpU+lS6SaCoChq5Fh/GdqSB6xNvOVMBLC02MW+KO9CV
jJyyppXV08o0uJ/FQSPmzaKVGJtktddQlj8o/rLoxOoajM06G/o+83pLNbTSFnfa2njUZthDqxJI
1CYrs09bnMMFy+/rS1jicNs9Ul0ZR6b0gvavHJda4cGhmAo55Lw/JUe3iY1SoYeSuB9ckh+3w4LG
vCke08RNL2345KPQyan1ibAyO/K7ZJo4CP0G1gy/7qjl5CWi6Ej3j1OH7WfaUK2fGLJB3D72QGbY
lfPll/eWwGMuSU6AtEgWqdIF75k4UPKhdM44IIbLFJyAaCxRhKIJNm2hKUqYqX6wz2w80uZlpcvd
rphW41T1k1vbvLXEkxZoowadbb0J3XxOzoi/gwquWf+/XpJz6SDqbBpmNkfoh9v1dBvgj8mJP1rq
ZYOrlmLoKuV8ULjwvGGwRYk9rtjHaRIyRJgaEEcECtE9vQ4HFO79WrWG35p8FQ3E05DBzVZZqy6K
Ak2ET53IfcsO587OMqcagrrKmVOlCYk1yls/gejRZSqk0fH6KBuDomWy8b7G+jslSponuTGEcQtX
fVCXqVQeJoL2qI9Kc4BSm22xZmqzYY6ygYJJW1gFjt2xbMP639D4vdQiBpg8ESfKA44yi21dFAAD
olA9miVUU/mZzrponA/aD87qKOrdedLBecP44PN+Q5pHUf6u1XPhWmGNOrK3Cv2y/rXbRNAFRoq7
jGYD5ao5WfG6MagEcyhFRnxR0fg2BI40rZeqJrJybVxKSZHLAlDETrVLpOWRk3KBlPsPUMnssIBY
wnAkhlfTJXsva9BpQLiUWE6LpFCzxD8t2vV0yYVgknWhi6fIx9PgkFQ+zuNMvJYJZlimtghjoYGn
vTKwRPP+PHjtsu5ez792ZjQ0DDJhJ1dRS7Mr1n9DaFXqR5GH7RHlI6acW8FeDB0PabENISn44zWl
YjafaQYa4uwPLiYsuyoB7o+JHaLga4TA3VfmhnRxQEn5ifOWAqyx6xXp+h21zpJ2wSw9c4YN9ZOI
ZwO88mT7zalGTlUt2o2UU7c3V5sYDAz2gm+bRBshdL9BIaP4shiuDKTADD3UkGxNoqCUeVK4AFbP
gNpN1vWSZbXdVjaHx2s0s/4l1t17bTtSILm6efkdIDc9y8vq7sF9rVuAXdjUOxnfBqXxpNi3RXTv
KtyW8N6m3EoRMFsARdA9xfJtt2U7jdvD8k/Rhxlx9jchLai5usVPEeyLKm3UaqfrGxXyPWbDt2wR
peBGmgEW5Z9H3MSxnCnWOg/LH/WggwWw2WbbNoEkKSEFXL1ArUDL8K4H/Kh7nC9udfmM3SING22L
t5vgxEm+9/eumW0Kg3TKTbYAMcuG1Wuzwf0JDJZdlJfqTaethpScbdammBPyVv8zZZOyyXsXZt+N
mdontRdHHkOs8dJ5IxovtvYZMsTTdlPsfCyUVklEUpRkdI0tXmf8ZYuRJHChgjaNCriYy+mg/41x
46B+quiqD/8Dz/nxaSEQSYpwQjCF+YVm3AAI8toNZDqDZTpl8yB2yFmZ3IKv9g5VDSOpYhYVmA/4
rPB4IdjrTsrcNzPPpykfEiGD+Ugzt6QG/o15f3xqsfai+7yuGnvX+jyVI67MTx7mI7gr1kRxf8nT
QKPrC1KdBVkxpcLMWNvC4ljTy7bOLi9vwczBlW5ynQgLxU5GiB/yrEsPFL0pwQOUoc3chgq3Q5js
Sc69o6ycPiKPcTX/VV4HtETsi8sa7NDXNoLGc7+7cJbTDNVfiaUcerHjW2F2heFdwE7UTsc3h8o1
t92i73cYjtr/20EANdk+psbBG/Golr4vLPTBiFn4HsMP8jC9R6prk7l8J6USVLA6pox0N0NGbiVu
L+SzAusBuAS+lzPNcuIbu9tMOWqysfsxDdfNp/54rfGKVDEO2gPwpd9gX/eE8+zUNo6n6aGXT5fJ
IVNXo7HfGQwNYtKS59uU0Lzu/gztu2HmrL40bbWs/Q/FhGJsm3yMwo60lqLvU6dyMPa7gaLdRtKG
fTIlftIy0PIULH6jPBDP8GyUxuo2BHbXTOg5oZ1HKlXCn/MyVahYnk/qhhvYNnPr/atVy2dOyfyQ
1c8xKtFqW4LwvwXDYMq0WSz2kNTuUQHZ59V726OeIsg7okl5e3lpz1AJ0vMsnd8q4wDBR35rZcct
/7keyfobhuCftZYe27SqsauLLOEtZKnzgPvjPx/nQhN0Zi3kgZJKlcQ28s95uayhUBpgd0Ns2gsq
KWlSk5oUY8Yy5W9pR9s+1J3wFr53ywuIXJDs+zsPHHxogYKDFmotTfvfnZP4T4XLfJ4SrKZ6O2Rs
yWO6HxoTRkYUXMDHACtmq/3Ar/ZDtNAWlKrPAE9E2giGvhd/6rSbxWFGjNwLvMZCnyH/6cAoLqrp
Ovo6f3GnZZwSfZD+Gtk8KB0q5a+daQ4DKp27SkaEQdC7s/URmWS8aHaX6rHHTUTrK6bOv0k53MSP
URpamGxOL9Kgy8UJk9hhMMQxfxH3L5Q4T3BQF+a+1lqB/cWw/lyP+OqbpCdHTfIT1+FMcZXHQXho
Ly04s6LwjqDq5S2i8QVg8iKBPY2QhtT3+Ck+jv70ao9l8gKPcsqjSn20jPdJgbZBntolcl3GJJlo
q8nULlnN5DonPRAygS6nviX9Tsgkd3b4jRK30qXtu4MJIS2daDQfUyLh7GWQ1iZ8VKINhs1Y/rbM
ocOqACd1YBzV2pA13ymSrUHivPYmJWsggA+H5DnBGZFuTRs/k2cXK186kdeenhoCfAU6hv8qbQBt
20TTwEHcCYxleZ+ZQcsFp03i2zLoopD7NwjyLE2Tjm3+B+qjGkZQzGfV5CyXDA5dbgheiF/SHspz
WZEM7IegBjOpaCoMrtpQkMRXKEsU4ksZIEuqOKv4NnQePXjlcZxnVwZ4N6UM2pLt4CBQfIbPe7OK
fc1MXMPBLJl+vuTIk+ai0XQcQe9qnjLiYVLYVbcwp/RQDGKiWeCZy/A01ztKEYKhpqL4Bc1pS2Kx
Rxe1S7KQGzzTQAyhI2Hzqu/xToKa4jyZI4KsfOWFzRWbrL+zFGkJGauspSfoTll27ZkB0d3ZJvHl
VgNLa8pOhkzWuD0vhJgvyETZxlg4CIf2ufp6Vmk782RiEVvhTXQuNJRkdfbLqgsy4tplR+BUB5qK
2tu6/UsgXF7IailYVtBRW5k+jlOMMpVd9a2Snjl0OXMJEG56hfPIzKXkAL4ckz9MykB6cA5CohzU
j3ZeqNziKAVufRBbtJ3utfOlWahrJtSpv+ghqm5VVZYFvjHtZjYH/9rHDYeJnsCpOXDnBfuCrMFw
qHgpKzCXcnfjW9tzqZcGDqRRP+CARQAJKRyQPebmifNlLub0m/2GPqINJ4nRRURiL6FHQfQJbwuM
8nuK43mRi+/lygS2r6YMg2+Y6X5c+UpEa6kNEg0J8ZMrm+czPE5x3X/INu3bI/GW4XtV+AOwk0Ke
hXvQ372Xg44HhlTECSQx2GhCSbrtf2ulllykqTAuHEud6JE/9runbBcqoefAkPLw2spi+Fkk4rVA
XMbFxS4j17P5B6JkZH4r4Fxwf9cLl9CB2jJfHmPyPkG/dDwibE9LJX33GrOaCoB/V2hthlYHm9UU
RqcrbASzR7bpJEMt/vsbQ8HGh5ou0xvGLGc4oJnyafPhVHUFbEx4fdaYlyhh66Y+OlBEfTAwhPi2
/9elSLUyyJLApcRfiToMA+orZTrw2iS9R5nL8t1S3OCqxhls8YwM5dKvjnk6+OUOwWqbmmKuzgZS
8KaXMt9Yj/nMD5jJ+aPm7rzJw+Vf7H8PnusL2fdTb3pRCND6VWB8x0w/D2Xhyfc2jvpM7rHZk/Ft
dyZB6JLIgRABUsJMFZBq8vZ3pwI+3aMymEOfAJQI4ibFyN5cYyoo8EOwNguuBHGcHV14dSzTrWFA
HfjM+fxfuk/vhlldfj4nZzyj8Ej55YuukvP9eaSQWm8uxlOjV387aiEIv86uOdbL8ktiVsTGTihj
n0KkedQ+7cKAebxHOmDprnyouXWzU/f6IvORU7HK16u8udNAcy8nuAwjmd/fwi4CI7Nh5oGSFEn9
DAs30LfI1tZkaqxgITxIoK2k6Tfme/zp6vKxO6e/bi0pFbGqeinippsyGFfUglnO8JlnYn/Tnlk1
IL+6mJyOVGMpGrcXiDX7PwrmN/03ySftLnyNvAHyBDvQTnHNkOTUkjrBzEUh7fcrCD61mKJiJ5Zf
o+PrW668Ox3M0/QMG+B0xuzzjOBoFoCwCAX3BxntXNzc4dk0mkaVmbtiDTr96JXSVytasBBCg14d
jhOBmUJe+42z3buZ399MfmuabpZ1pRx8uOlTsTDbnz+APzOK0bYaMD31hLfWHQ1q53cI8DPHMwg8
NmHKBRxVmXLiySM2GkwE1GCrm/0SfLU0sJIqI373oyIgDd0jsAxx8B/U63OxPtqsrAcq8JtRR6pO
qOkocYuu4SHWu0CZebSiSGm3KdxmpG1BA37mVSiWFlI7l4Xv1Q4HXcisnhIfQfNjDfrkPB2ur4Lv
nASEbcofmjaFPFTCiWnInXEFo2hPInHJci8E41hwJjw+O5T/snTjwYq4oIANRG/52omRWDMEA96b
vslNZv6RABHIWQZdttOmzMsLeRLaXFUGi+ntePFxRjdpTivuvrAp8pIfOkzjgs/2BxmPRHxf48Iv
9IOGIOwjv6UQR9Ldj1WMICodV9Ulu2vumJbbFIh3y2v3Zjlh7GRcr3UcCIgLltth+6PJ8jn+8cuZ
+6yGP8qu3uaxyUR1TgXks3bVBPRqBOrNP032H0yKUcG10Kil0VuTGjR6DI2oSG40c4hdU9LCoqq7
a9Lv7+hOu9//xJtLHwnhpsyXEiTq+5+FT0S0Xg4jtaYOgovcTQDHDIgSxbRUlvTheEv1AKUdD5hm
El1Ux8bFtCUOn1iRLt99x3DJ0ha+HBzxSu5l139/4LJQE0aFWIpcLy9c2GFZYI4URqVunHgW3mVx
WwayqsfGENO6xFuQ2zRMo5x0dOkr/sQe1id5w1PebEX2B2U0m9CHuDhAhRkecPUi6IIL9Rd9wBmw
fFBsIrsdIwPr89Q4u5RIpWPdjBVPQwKO2LQbrcFqZT6yYON0gHasoZ/8idHbE+8NeJV6oVe1gW6G
POZuIoWhpbCGyKk/k1wKBhHLAAHFytC5E+SbDqABeo4R63n3eZmRsurVMColdSR0W2+FFkYE/kS7
Wr/vEC3rIaRO/4J1PPNL3kZ49gNudny1Nr6bTaHqA3BERSt2cvxzWuhCooSBLYGqfKcQU4BsNyR6
VJuYn7p+oEc/o/t/NMY85wZ8mt2NEDGpNX6Im7KW69gqFJspSyMr377QFCSbNGZMaCDgisuexQ5K
pLyisX45Ya7nmUq/0zjaEPLlVJq5IVLRQH2nmCN1IvRIJGj+iSZU3WyRCtVkQOLpM4FdfIzx9NQp
+mK+JL7awSUKDa/h/uDdwtxirZQAkYCfJCSpCLSn1FYvMHyTkoF/ZcQUUIseAsDQLCDBhYiXIuum
SZCp9vx/qXCfy6Nm1VPjBQBCYvpJBry7cCHeFVo8j+Z4eteNG56Oqt4tm68gt0xt9ZtnxDN0Ah5x
HU/1LxHa8qfBq764hznftmE3OY04BZqS2AarFIP3FekD0FcdBwlPqVXRKFBYVQcBASm1QnGmpWwi
fhXK2h2ev8MU5TIfAfkPUmIKJAXflez9wBF7OEQqlDYArwkBPTXLH4EUa4oUjuGlXH/GUkTHTi0g
OIXLq8RuYqcYloKZOqJz1XX7eZcg7OQgd/1vjXguLuNkJjpH9iY2UpHe8IcK5hrjpaY7hgQrS/Mv
ur9+Wqch9WKYD6jmZvUYVfVtnZ3KhVio44IPTKO1yluvbz0ZgH6ch3gkIeAE20j6Qk+M/E1MIJMq
vwCCJVLGAYwsSmUrl+1/ywQpmptqoroOVVmKdvq0hP3iQtJzuvHLY6oyA7tv1yNWb3HXoNuwdTmY
lIzlVbgaQ0Sh4MaWWU5plTZL2ks+nIzjZwyCVT+gnNFuOnIqI73uSJzMCZjcytB/hahs4ePlA3qm
YXKEI27B1GgcdHMx+fufq8luOvnRRZf7OAHSEkluXVfFoRi24VyqWV5ywU1S2XmNYIARMxDTm2dU
dEXYNXJ0Vitzpdnd2j+OjbWq8VCs3NbAE8oVE6WLhlgVavwrZPa2FJXtS9SwsYcl10oKKkplMhN1
SEaUoTTZ2AxSRzo6lVkmnN1zH3F/qg832aR0u9seS1ZhGmgjYIDc3cbpFLuj30acKoSvqNgBkjyN
Pftd0lq89dsyNJCDdnUDPelMvIPG4FUZSuTM0xvwMqtOrfuRqrZAZp9XPDAIA6gidGrdNiEQgK5i
SEFyx742uqQT4d50H2qxVc2ApA0U8g/1wh5wXRmLt84Cejqf2/qN6Y0J4wGwAyAiXutMC6fUWVBq
F3BVCLalq4V512sTViJbGc1nS37wrShV0y5S1rU846HC8k69Pc9jdgQgcWuEPAQyc3hFDNVl8edv
hYocOLllkivtUx6l/x2IIUXi5M1UY9EgoPPoGWS4I0aZ7+MjWSgFz/SUw2Lo7/fkQqgx8fBCwt+u
HZI26jXN4spcyHHmplorflEZEnPIBdzLXf5iTPIIFpjRcOE7ie6n4Hr5FsJ9wg/PrSwOFoVru7a5
jnxtQ4El0FE1Q0Py4+HvF7kYU02V84U+wbQR/sZvZFjPFx8YjkuGayT0Mt5mLjCQlWZ5L14AyM7O
5ZrIYBnhcntRMaqOsMPLqt6HUl/zN/UbDmhCTSlFbHEpZNNp/kqinCXrhvIFhV9bjPLdmHJGCCDf
1YGrmwJmmpJQxaTnF7BVskDD6tgx4Q5ftFZLuhrfKaKABFTYNqA3/uy7zaKZbPI99JN+9XiwltL7
YbShbNS11YJMUfPkodcDMCyNlJfvZXQyP0HVGESTdT8/2jvQZCNxxzWIWL++OSwPLloZcAqzgajp
IpRvZUJOk4foB9Zhb+T5zsMGQ8HUFPkbrZt2YsMBogv4bXpQ9w00dmoio7HxmgoXBLaMD0fv1QIF
FpD0t0pLq/Ul53nLLEz0Iyzzn1Shs9j8r38+jHKf3+3FXPUVGSKRl/xz+EQy+F/dDubFbxV/xp64
pF+2rPnteOgeqgxISu447FDDUpG+7NPaV3wQa6PLN8IEunnSdGnAwy5ZY11eFmdYq0Ncnvj7hD/f
hfnUww6Ey60bxNtCI3fEKDg8fB0wmFyfM3pW30BVWhq9b+bo6Yo0fre6YOhsNDGX85MlibQGJgJM
kA1KEHPrTNtjeKfDp9rykaAPYNRv/XTayTJNrQU8Tuh/2vAWt7DX9eLuhgqS+07TX0LYdtUbGr/k
4qc6YjZugMsGFb/nO2niUSXW8tN7kQRpWcROeFCM7NSKtb8MfTVgBe1XXajekdGG+1U2OPwmuscv
MZ7c6TvjMBQqqz2+niIlyONi09B9D+YlODKokKoHf1VRT/CfIUrUZCiGWMtA5YdvLccHCGjojzTt
liUZG84g+HFBw/G0PQ93O1dNoq8H5trWh1hCWHUS2uYoekU2N8QXUDHIAsglBhulrnzcX9VcRLc0
sYyQnq7D63YEmm3vQAeG9VVSoxmv3hz+6FzKD6iEVxJG8T+zW2KWfqBAfSw+/tiR8VGDKqZHa2bQ
vcKvlal+FBNknZ3VOOX4kxJJVBRl2kGflG33DtmPNy+Yvr/38eWWwh9bqJAZ9D/vVFvYbJsVY6mv
NXBz5AUkFVts5BbtPqKY1K/B7ThWpl9FPlLHkJAZsNuR/CfDpGaS2lcLM7VUTwIbq8fFqD6TujRd
zcsWu4fb+8l4wl8NzBXYZJqu49nQg0j9PTiDruiCnGqbUqcPjEkzd/Xjw6HyKalbCe/NdqCNYwcm
guJmU0FDnccx/u09yJfzZYQHsPX2foWtjde+XtjET/0Gw/TpjXo8nkcpl9Y25mDjOpdR+3LUKOMm
McSW/Oyp3WyCQFX30TeCK2UD/E/OjMXBguYBHuUrp9HsF9XI7szIgh9vB6QoAcvy6hvOdg8hh77e
oSOHSxjQi2IFvwCaM5DPJaqdZNfN1R/oaALgiLVcKYoI/lI/cDeXTvo/GAC5zla3LFrwA1fvLNBD
GnEMwzLdU84ZJ5bupx6I8GaFNUSn6xxmL8qJVNmeToqAJjVmZ83uRrMYQ3qgGMa8KFjulvQgemDp
q14eVEvX+miJ/KGjr2qhg5dlEzLugVIlNZ8uIz2JAR5N0vQwL4vbiXMMaNtsMsOjBI2G7GcZR5qu
426WQVTbi8O5YVxWgx06zey+eE/A1gdkq/au8HrkbYqYeHPFmk1+FxdUZNkuJF1paN57jYH7C5Qw
GISg6otaEhsPEA5nc7qz8VWorPE/6ujcN8XIB1MsrXCKEZYQ9aYCozgZMMtyNNXDj27Qos5bD1sj
fQEqXV01sP6XGnLNSs7mPqbjGHsWutFooz120u0hpOtBb0tbbVAo6+fQs3UCaXlNDJYrQZicxXmY
KDcndH3yFsDETU3oIZmeh1q8M5eOzYu1GLk/cSjzwTbanZ63U6tMtBDANrrPUWyjv0To5Y7TS51C
xxkCARiTBihzVUPlteW+0YLMcqEEmZBlcaDME9X4/9mP/ydTZ6LQpzOyg7GVkiUrA17R27xKt0s8
SWtepTnuhYk/8xEHWUHVzO5aIke4erGNu/5TAASDcVqJ04FKw/waV97xa8hRl+IaN5LAuVxl9JvZ
VgdECIzVZREnLkAz8u0W3Gr7Mnl3MKSsUTQUCBoEs+DcujFGW0YILvO1QIDeXi3XxbCmwPaoKEap
ScUBIkoqsj+H4rCzphlyanqLXBq/Was8qxE+ys3EbldFCtD6iKGM011nsiaNlmECiDzxiY+5Gvaw
KZKxbafr90i8RI4F8JV3nBnS29bb9L7blYXSkb7CXwS49hR8drtkM8ZPJutHKi9e6kBQplAX+xbk
cTCJsFzT0LMo/YScAoZIwFEEo+tR59Yo0pZjtlWLStdRmTFn3GJmDs1jwG3cZHCZjB24nTk+w9Xp
Q2EiPwH8PjiYgcwV9UOLf5334OSf4fQs3YbsmxvmuGMCr1BghTPCxYO3SBWPwIgW8qoBCYRr0Q5E
nSZJzit/ArkAHlZxFb1MqSQHQYjM3/bhV8GL3nW/LP4KCEDJeBK0+v+KL47RC/tDWSRxz6FIMeO8
mA+yLZBmJrz4ryeOzqz3Jowu4vMhewgxmBV3Y+gmA91ttI4NLfYVcmNoLBTAwwuim7o06nU12hqd
0OSZgWBZ+XcZ4Q8r6JLYHkII3GzHtgMtwgi0kZotDTMqQm0Yca44AkgNdDoCYtHwk8BBF3a2/QZH
a6O/p/5/0uT/lyT3OAndv6NgRHzLN8rVcXo5psuyUbcSFZFxJoRERkf3bNK8268rVsl9PNGYg/gs
lOyAnHkm0U+4cc53SAuAqQ04jiZHeG6xokXcbg3axUKcZ0OaRF9G+scqYex9wR0qD/oZ96TxfgH4
V1jPzNprqCpi1yZqyuG/yrFJxwgRB3jlmaZ34sxOf9IbUSF+nFUzAq5ROsZfUUFBXY3rs4GKYc8U
wS/BdNWTRxsa9AvWrUY7i5wCBKveXdk9KBH91sPcbHsiNYIcHuvGKJ3vX+jiXY31FWdRHmmwqyKZ
aWkLj3dXUfg/hYYWBwkiEESp31iAwmVOiOSPUu+H2MnzLNJg8iWSRmoE0/x5IgBW+vo28rZw7diN
W4BqSCB77mxC1IK6ADjZcR59dOti131Kpu/NJIfIXmNMFdxg2IuDhbsodJWfyt21cek9BJB+Tk92
7FbSLSOHyJuWBw4h4L2UUvrU2bTcFOLxFnZNJZ6ekqHsIKHCVaoYmODlxO7p4K7f532xJpMlYiKn
ga3lkocUy69YxxpaDVsOac5HXn56quFgasjejTgIa0JLI5G23hSlAfQUI4IVDQUw6j19yM2dpowx
w8ugXiwg8MhQnpNIimni1L0uMiywCKV9e/lNnulADKSHsiLum046PastVV9ITf0Tb+AJJAE10Isj
ImRQKyf+0i+nciOnIrdSquFeXwAG3dhJOtR6i6H8aP+EL86bbOdy6AV/0+s9FxW36gxXISPYKjU5
wdiFOYuVG9ZvmWK8hhyjAob1IvMQBm0HLnbbaLFW/mCIv2urXj6Yy4kjcULd8/LF+zO+3ua3OsJh
N5kAQwvXK5HieVAhCCrZdGsmNJG93vF3czwdX4iDb+BSmLRUL4iTO8FIqHpq5RmAK29ZgfXE50ms
iVDjIF6LHKUOjHKRxlq/4h+ixxCkopxzUt7hrk0ZOC68mXY06KhZluK7jKzNbqMRGZjoEMtzV80z
VnGqrxxcZQ6uvoOsfULfzKzR9iSNFXzUGg1f+Id7t5PtpI6EaQ9ZvLoFWFwUTu/Siu66iL9EuriQ
TsdbwAMmZcu3YW8163Smr2vnjJAMe4ewV1zqSECz1bkS8Hcznmk8UbLMqDNsckrk/fR2lnzz78ee
/gg87jiYVl03uyVZ0Z9R7mxsK2S1HDT3G7SbtTxDMxlMHUJRDINALsE7KoLnZ7pgDAwfjYEPMNjP
6p1ywVtz+oRcYn311HQNq5Qayp4oCVXtfShtg32IbikrfVqXOrDDtzs6Vf19aadcYPZjwbY/OikV
7MIXjGTTJ24GV6I9HZZLdRhK6H+gsySfWqU98DYTxY8zC4Xw1V9lqGeBUyzRERPRbEXX9k1woyXW
GhlDofj0+YrcumdMOi8TK/1ILe7MBh6sjMsVlhUIj5fKdvTEZOK79yMJ/CaGLQUXK8lGISGooCxr
g19fFVArcgnxp1a7MWOy6CY7tVY3KDStkrUomubgCPdotfQq2hHFxTTef9nXhUpejydkdzRBgEoD
jQvX32STVx3YupxjiZekk/Ic7FKfayNFQeDloL+H2bv8e71+4sTH6hS3UUapUQFgvIplJUdRY4lS
2medNQv4VwbdocdL3iK9BQIP+MqipY+FHb9icXHsn/Gj5BhrOexp44bj9Al5h1mDuHrZo2lbODk9
2rBeXU48z2X/ZExtshhO8PFNFiUwGltCTKig9rjHG7Apc6RW6x7tV9mP+HNU36i9YBxpVHuI5yfj
24rW6+x5TKoF29hnxILjMRbMTrJGVern696c4pgmWXU000zpqTiUfO27CJfOpLb59aoebWlJg5Ay
OuDygjpkOHYgUeUib6SxObDEHOrwUEWx39gREJOhmsnR1vqdhqBCfuGQM8azfpND070rucX/HVCh
cM4R9gzRssC/rgcKFCqNEYOU2gIcOCAaiqORn19TXbUKNOQTyq6Q1hO67f4fLxF24sI8xADrNnsz
DPGjNn5O+o0tfOsSClH7sIbD1Ufx2l4Z5czKuS/x4E0lPg0esoV69rzofn0K3yJzb+G+84DpmIxT
lUNXKryuxAUcKARCJLfHNFj2DbHQsVCmhhm2ufZTmmFbqIr4lJtfT5gf+0/PqGJ76szEJh8HGPVs
uCje0oNcI/r3dlQQ3Lrst6yKJjwmVPke/3P3XwjN2/0sJ8gtaiS1DrrSGInw2+I+De5AYg56ipQl
0IP4hHzk9AHxkS5KFAJ80/W77kdmy15tjUhXUeKf483zLeqHQbhsunHW3/SK5jL7nV8+3Dvf86Vw
bwz7xufR8yoHekSimrm/XFBt3sNsu4b+Qa63rGcADe3JcUbf8jc5XhSmPOo7D0mDRsljvM38s7vr
ukxpRi0y6Ulsztds5A55c/wgXRTbXFCRxY0DfO6LMqu/HGz+9IW94pxE4RImFCGy6Lm6QaJkIwUV
WXuK7FklQNAVIOFke/QEHYYlM16Zs1ThmCzb9TfoVe/wSgI+pfWzkIaUotX1lVjVAvVsUtWKDnxE
IdiDNjaUwiX0Yo7EH29XLO8Zyt2D5dT3gk8KWOW299K+867FX6JRQx8mo42d8gRwDzc5kQOEQFPX
HkxXyLvzjyT8UHmQrGQnNBggKtNRQoczWYQTc/n2/t2b83WN+DOYK+E6FD6Ou5b8VYTpUHlXWRcF
tYGhYK1VyIQ0ynmrEcCFQZb/T3oGvu9eljNQ8x7KVwH+WuQrVIeBF8oiuneXeIsKy0SYkRyrKr8u
GuJZfWV0FsK/c0ChEH4QsbgDLiD/amcF8CtLBm84Tntfe3z2iIB3NfIghsOk43Mv+u8cXJzu89o6
muXzkl58elndd7e+oA8q5DXRp5fKczguX0tbSRokXgpVwhKCw9QJnt5/2jtjMX2CFauAE4jSvnpT
zOykdXMerhx7SSQggNDe0PIM9RgQbmjJpiR+mlUiecZSfzcpwho3TD/OjDFbmVyx00LNOU13MCLJ
ltMenSiqxZgeUS5qTXtR5sC7YsLphIIU0NwjaY+d4r/FOGxFP+ghtJUGuGUD9EL6YZLomeenpZx3
S/aq+2rtGfm9+j7NBoeunaneSlIi28HsHUcavD1hTk5KupzfluFik+TcV183MGFvcnYMpQE+uq/q
Y5LjdUil+cMDH05FxEkjd0t46hsrGXVPSonLlkQTltG/7caZ0Tuj1raPpAbsOjb2Hisyz2InADRu
cNzjyPSyd7sDAOusWNnYkgUfvsJsZJAE0bT+N+O8nohNmn8XMIhqbfX6HFL7TmNnfrjCsaBKBMja
TelLOiD0GwgkxGsMi/VRChhTp4AhpL+PMUX9phYQn8PPB82qJ5yghPK76LTS50gFAtPYI5dSzYAO
X+yny1azhTA59Mcw6ht5yWmAhO3LoovQ97gKMwOpmPzgK9Vn0FFUTGca+4atmtVdcT9BRM8qXHNf
zulgVA/Yd5PzkBNr+478QbZCpAvwGjGCb1j3+Cvi0t571CzvvJZkMKHwYcVH99JT4Kl4v02ouNxD
u9+ckzy5uayHpmF55j7Jui630HnaastGdn3QhjE18OYQmOj2GIDNm7YtEQYcHEXd6o6hrp5JpPgu
TVkm8GsgDHrNvzW89/BNf9PFnNXB8HRWr9os0k2zmYkh2xOXtp/B1UphKDZPfj7TJh2AFnspnNMy
gwZeh1eYEoWZu4Z9DSAi6IwDL0eosDa+jji62HETjBhgRKBQJs26rRBKnrVj8WCCU+JylDfZFGyC
e4KjRy13XyHspiRYI3IcH2gH4ubrGZZ4nhnMUBoR2KyzVmjJo4KEOolfoDjy4XJMr4mHV6Xgee1K
Gez0woGhWQkGJh4VksIKtvJHOdzVBeP+3UAFeFapBK2aLtnqscPmzo8mgNa5rzObsecH8U1CSjT3
xsuwAZ+YLgRfLJA09u3MEWAL8Tgmr2RoSYmHrxAyQLepKs7Uyx0wdvplDzacFbjoTnVPAtGMS83q
jnS55Sm8OgW95Ik9VHHiMdZsIVqmTp05BUW0wMt2c7TU0xzMnAbV9k53Nzn5h0ZEpJ33g/XP9hU0
JshHKas8O2PzmmKyij0fzt/HuFFqcIKNsLvzmGUheKX4gg5P8IfpqgUY4YJBNHlFWXwydtzcrRD2
VSlyzgbOI2SJTbyw+B+tOh2URn3VcMLYE/itfp9oIZeAxUMLFlKQuJt00EaxSEMYwykMvuNwVnsb
0MR7ZQapwWfPQb/ll0GJ+x0iREKfZkVfVqlme5CiSCfe8zVyerQtjo47qYY0iy2uFrIngHbwbjqj
3CIsuBG18X5iWJnu92Hequ7Jsw/2Ie9vqVER0lY7/nn9/uv6hm/PzYrkZXOm5Y9C0uTvFEIQuPmg
qLnc4XiZrVWGFt1C2fFXCUTTQr/plYIYZSwun0mYkPu+D/cVgGJ6vEDaLFzJsiJDHKI/VX+9TxiO
bJu5+h6qB9Dlp4TAcL71NIXNRnDfG1DNP0MZIiJ0q4ES6YuGBD3Y87MJUsUHfI5WEOvPOXZaC//w
to+cQmiQ/mDxtMGKKpKVi8DMqY5+kdroSaKPN6bfQPB1nmdR50rr1rvYz+uZz5gsA3ULLvFoI9RL
Dp2oOGfP97Xx94cCSu5xQOhf2Hyc85iKmc9XTwRiVvhCsNbGowD3xXruUWF1LFoBDdp4lDa+QaJ0
HQnSstXbg8YwPcnv1h/ky70sW6cTM+h+/JgxEndpDw4hn+/TLXSaWEL5TMkWLMriZiZ4qGBYNXoh
rBt11jk0RbSF/rUcQ53IxYZDAsGRjYhm9l43mJUHT6aN7NXBxUuEdkIE+wE84He8fHfw04NoyB7c
zVzn+Q9/+FH4fRNlcoOAvaycBadI3dEFlds7YyckVmQ+Io3lsv78EbZIFCxfgHoY8V/NAglXTCOl
/Edy4OhrJQyA7M45NnHGdKnKBQMeb7T0N4BvjWGmMHddWf53fs6r8QrqnYlJ0xEblh56VGEJRa4L
AR4io6u+0LJn/MSZy0AM5ogFO6JqPzTK2Css5a+FwjkB6HcttspYuxeO8dE45jH2kC5lDIx4N88c
IvK2y+J6fGyA9qEqDepucnu6Qo+wctUpDwZt62IBCvO2wzahgdhBFFMDRPau69cBl/SEzW8w91yq
sKfimILJousEgIs6MiK07r28aTHdJBJXaqVwaAIN36WMLdLDpTmFjNF1cjRd0BwbsFUeWTWr+4aX
9F3WLB3nI3LzCCWXtJGszeKou4UCqPxoSqfN6/K5aFnRiK9+tgu+7EbLWNtzmZ6qB1IgEughL5Tm
mmyXSlui1uRzGQOVJXJRDJfoKRu6gx+26agWeO8lei3m50p1ERVk/wGO8zoTh1GSNH8XuArhfM19
mTPxxBhdrx8Y3gNPf3htSxZ3gPlRW36wxAXLiY7TyqO4VyqFQmSMCmUIo9CSQ+TZbOPqfL0ZT+vj
P1AX24yQFGxnVBfUJ5pK33C9zQ7fabGo/O3+YJDsAh6eqOPZOAy58kLCnu9wdPEwV6xxEfCePENz
w6lc4Yawv4oO0xo+8dlPH7/aDvhidIwA/OXxeC2XmMkrZ/IHr+o8sDDj+KCYONmKSIJHF3Jxghg6
1WbE7lK9YX1PSn0+Vw7tpUOSiO53PbuSETYso63q7W8Wj7jzL5P8yf2yRcFyqBWRA3wrSQsw+y7J
Un9z+jSDfH45BBtPypBV+HQgIGi2z95tSDjG0Kj17CeuA3Bns1klQm44gsXKg1zEaoPjL5jQX4CI
jHLdjLzSLIc0chUKbgARXrP7/Odg2gCokYxukJb1XQmzJ7bpm4YD2kpSuDOjQzYzOFzwX6I7tccA
5lthnLDsgU3YZ82dEhHyLAKfeSf+LPmWAIUenUkVlxse3w4qb5du7Je0s1mCMO2F+hKn81ByUNU2
9lgsTkUKgCQS5T3hlgkRNZmQToFc1qnNrLoMNgsRmMWvW6rZ8uikZ/qhu/Fgnce7FZzAWWQobuuM
8xs6BPu4ebu1LqMBsDX1Awf/ggCtK0ndcscrgZYX2GWKOOJw+LKrXroqzXfJaiCfnZ2eCHxkpbG8
npX9FAfyUQeDojjdi3StMUhI8Yh412/fWkKJTd2AEGX/ibyX3EqdMzK6s1u8BQVubpOpW/tgl4R9
edNSOfRwzZ9qbCPPjaCmMu9zrUxvsa2JIc1MRDs1lruh04AXhr8BKuGYDpoMf9SU3sRUH/rILO8/
XWW5MePsFTfIzwjTwUtymN5bvleGZrr22m/ODwD4/lWKoocGAnlRGjc3unQKe9Zup4hBAo4lYMy7
TC+1v91hw9AyJF8NnNIgH9COGAy0aWDG6/ZjNul5gNlogoZkZx+jtNRGDiBoBzSjtOwRMAzEiUqw
FojWtGbHe9i8lkjkeyjdwwSimvPbLvnIcK0UGUSIc6P/52mkm/KTYY7rzdyMh2+parW2EiEXxUmj
KE8CtNPGRYPvZpYF21rd5RWA9bWSBTDVz6AqI/ykxpXNyPaVWreCUm9kpcAu7Euu0b9S432e3woi
TXQ3k6duFmxpB1JW2f3gwb9WEK5UoYCJe8NNDntxCajQAh9VkZYeJoZJVf5fV/Y2KTuQM9NTLhzj
CzyvZwex0Uqmg5v1GiYAdlOHyHfjz6GrdEx1WpGNhXNAqa9J8MjmUw7EAjFO0RhlVLLmZCaHjS4L
294VlQG8QcB1i2uHHA6Oz2XN68det/wHzSO9iWd094gvT4Edqoxk+iZJwlV9R1DLSEntrZwd9FJV
5Brwzo8OFmB4mgU94ezYe14XTSLPryhDszLAGTLAgKCLpU3vftL+ia6Y7yzIxb9ktR6WiaCGKT+w
p4pA3dIk1jlS4L8derFZIQkg0Fzb27dmDF5ERrC4cNIA8b+e4HLX4YpE9G6xtIwzF6M5wfX3QF/u
+g2KNG3eU5LjZHaf2s7vAcka7c5TnfqDxirGRm29GfBviiJGgCMja/yJseVR5IFOQ+rVGOLR4sqC
71f89h56uf3Cncpdfzgt9IkuGQZxKY/4ip9j0kDfdOSasCNPCT+7FD7oafiCZnU6lerBgmR9J84M
rUDPzy48tyho6xZZ7F89d6nLaPeTlidQsO/rS3jLMLK+cODbU4vesGApiFuINMOBIcSC/JhcZKXE
yKFP+JX66ZivxLcNSa4NWaMLXreO5Ui8G2guSjcGBzx6txyiNXpdJ6ggyGdE/7IAM/OboX4NH5Ao
fWh4NY64wHC+gjhC1AyJS1oxP7TKRPYGtDeE9d5M/vW80neO1HEoSTauKTbpQrtxJ6oNWOiySZZy
wbHTvfaoABs5J+wDzKyNQEiskPOAQ0m6Ue/fK451+Ng6BBXZUhFGdSgfk95lodE9fneLJF7XVbl6
yHIMg2Ut59mvQ1PTb0pu4Zq7kF0TX097peLvr/SJxy5uOsNJaEFGVIVO8bWbBzQzxLS52ZRn9slk
iWTtaS+4fFl0ooTWj1wOymLbBjJ3vZK2JBQu+DcNk2JRb7qz0m9fR4Zs0R+Y41vJhon4Zq4MIaHx
lD+uGQ23hK9+W7l5qVshtxAxwx2RPrpFhabnO7IbV3zrFKqxVf3YzpNr6fa8DkQZD/IiCE6HyFDl
Waika982Km4O/e1Ecf21CeapRjXyDazPepgKf4YvbDsrAMeU7UfSGbJxEK5ITWZWqts6qrSZ4iab
/cczjFpwOc+aSS3RmGQmSg6YMREU40Z3w5HcO4Lgjq8EYWDckAoIQPqrp7sXMpaaJiHrsz/BivnS
rl1CExy4LNbXTAfy4j0MHLlKTUVP2uNn7MSD1n1AmC31owJ653FD5QIerA04omnvLg/Pc8w9+vMz
nBeKbrl7sBr10vI6XaESR2GXfDnuyFYFxRN+4k7KKHHYPli7g18AJ+kbmglE52nwJTzEh//9fb/C
PjI/VOf3rhrNYB2U3HwhPMGjjT2+Qau/FASZ4HUwXOhCqxNxjayqqWsXqDQsMy2acrebCQXw/z/D
qBx6nPjSoCjGz/DozeBYLSLM0d/rOdNUtK+3uqOgLiy4thhk3smmlSRg8bPMLD5kshKkXidSbbtt
k6AhCSlP0trwNvUJpqUbR1xIuRm5OYMdtDAQI1dj+uN68r6AVEKFD3h6ikbVgEnxn4alZ4M8yD5a
bdDFMsIVJIQ9Za/LS8RruURmcqP92jhdZErueHbynedL70XC1iGS2Lu3mkaI1O9MfZRoTUbt6a8D
7mJ5ljDOPFrYYQ0ztVluVJHpiEt8XQD08UmStx0YxveWyDB+9ZN24qFbQvsHRbY+kFZK28rKl+Ns
w7IdgHo6ouFQvRJX/3I5J3OlNv/cTp7BkV0sQ7jl8x8Lk8Z4oLbSjEGbxK2Ppz9eWBBLZACFmERM
CrJi2kZiYSRjCQsNqEw8Y9JZgBs6OqDseZRzNJ0a6VvTfZYOrAenqB8BQaq3Hrc0nO8lVwbJHVt+
47X78WvARcYKamfKtbIllPZ1S/2J9l/KoNCnNo9RI0O11/lPGLqu62frc2utSrH4nAdoqVe/oZBI
mmoM/e0Q8ujEww55s+ZoCxQju9c4mhR8gt2LQIOHjHAgrt55myTWv7yhmbRaMHQexfx3YI3iSJ83
OoPnEQtyhcGDB8pzv2zoFETN8XBvvaaKBx4I/kumMhGbGQ+0FW/hgYi8ofEMoodWFzc4LOeNlZ1q
DYnoQV1fjC+nHD78u59tVpX1RFOTSxj/X98+QxJoWJRKUeYrOYkW77QFNfGwF5Dx0i0tjL9tiwZc
kn5tQd9p3sUfp5R83ePTx6dr1k7Iy32WJGc7xwf/OmPU9n9lEmMAag4giNtDRv4Bz1A+NFIiL+lX
4dOaHg4Xl7fzCbowwILITmJyPhLVNinjEmGcnbGqfeo+TUbRFBoyqijoccrMjK/HkFeq+IcPrXUj
XYKcwm29jNxQWGsR+CE5J//RyFAoqV4mdnSxp/T6I5teD3ORSr73/nyxi6ncNml7mDl0f+ruiL1G
GCieaTjZFogwjw/wQN2h7Y5e8j6dbjNaUtJtF9BWYPDbmny20xVPZyBGpyqM8yK4k311IToTsEmV
02C2P5q6kOcBMWdSawUz+NMsAvhj8he2dSowXd8pPeAHnybWhoKhkTBkqobRvWmMOMcWc3zzwY5x
kpKMLd7gZnxMMUKFrrZCr5Xujl/X+QyUPoBAWhoFlxX6zfWuBzziTte/FLMIezLJ8F++AV4+zZlO
rU1BIhjclJtfi4lPZ4F8KdeiHs4aoCyO8H44/cKTq8sZpL46oHCW59HH3FEtbRRgB0AFWkn7aKyB
1BA9qBwd3ZsEEoJ06VPNAPos62YPDupsy7caG5y9JYCWuFrZIrq1ffC8vlycKoOt9HbHmRdZ9DGJ
NWo8yI9moWy5ur5nn3nVOYrld0bxlYfUNKyXl1UMaEY4o5guFJYFSedXkoMM6fEwYL8W57st5xg+
2Sp0QJYZ6oW+fM6SrZUDleezeamAgIuoi7G0CEuDs5QRE715SaJQzXd1OoC6nSbRIUTbaGd80MJs
ZPO7ZfwUbCQl0M83N8FHwKUDywvpjB3D1mbMVUpNSlL1l+6z6Yos6C5b0d+yWvo/sCKxBuXBh/m3
R5gbDpUcvacFFwnp8/qV9hk2vhwhO7UJib90pPaVXqFQqBT9okqFdKoUK0TomlUrGU6+vkUTbO06
1E0X22veqYCFcmZRAubSP93+RLjLLS7ndINDFvCR3xOJPc67leu77AFKfQyHyNwUd9hNUdIWLjqS
GGu/VSzff2rsm5c2a4/i67SvSQzPmQSrXU22U6L+lMT/lfwLftKKfkVXIkEr/lW9K0wgr7McW5hx
qeUw76yhmgmYiD/aPssTXbsF7UxaUJNzavySgs1M6Q67JBFo06D4GMr9KC0jqLxXftE3PAM4TH2n
knRbBQrrQbqRk0yHB5qEooX7WHs0nNsPLn/4sZ41diLrfGKDPeFj37LPSjeAU5x4jZyJ2ImtT/nL
AtwCgwegdvO75bxonIuTlydhof8aLMCvk5UELIgZ3j6DVnU+ce/EiVL+QVryIgeHpVGknUyGg9Ql
Zm3/7O9E+K6boai8YwEiGRDUU4P85RuqBv2RS6D7IYUuwzj5hKd8Tkk5Zyb3Z5LsUMXJ3OOWHJAe
cdBKsdBHPpmwq04XcbC4036I+VKVMts/hrbcirzDaxbJq4O0HCAC3JjJyEKcCIhRIstTDb+YpqKN
WZJMG2j6k549u2BI7mSqVS+BeV+xiGUCg+eSQsPECWcSD/UNemcVb+UtMs28bDW86CFsCQeBjCMz
goD61C17o5upHYhcd68ICsAEeT1kOP7lTdvgX321a98LEQnJk05EUuEIiwvaHpWRIFZ3gwkZRw+0
fbY0Tigg4y3vzC8gWlW9X+eQhl7xtJ+WpAiW030cb2wIPKcRqOMIxsgyRoPPM9enOLTrygWMNOar
Ze1bzLiSvBfkpoCF0t+XgqpHbY1OrCUZBWh3onqjI95Kn/aC0BayCgzMLLjK79GwLFPU/YXwNor7
h791bdWffD9NkuAiDeQBD4PKy7O8TZPylr9YYDbVRhL/Xd2pWjFy5Pl7buEYk0/To0J8YmoDLdXA
ARquyPKMWzQZWKW0OpJNzwKcqv6GMY5LSIBzAdMwMVZuxuB9eXlNd0gpFyhDOycVCkyaVZ3LxzCz
1BIWAFN8cJgpu+6HpxI8eFWdQiXLP+w2zZYrgGfKZ9T9lxO3sBHj72PtetUDYORd3VPj3nDvDklt
etmlJkAKOzT/tdtESzwnFa27FAKUELTC2onLCn/rvlG4uoZPgYO9LDf5ZF+dw7lXNJU8zr6kAnMk
hMYc19XksZ2NVgHXLaARPudyw8elw547/v4rurKlNLMRHdhI0/kt6KrTed0PyBwS/62a9vhqAMwc
DsPNEr1QjRG22ybTABpqk8YJoWRtHZjxkbKaLwy+C3Fj4milH1zMF49l/e+oG9+J7cq/jPzMrDqx
Mm8RzfgCi8LpDxW2CV57msP+5ftCN/t7Jd0ZPu01g+iK0kyBxvc1VgUmqdTJKJ+03q/7dU4h+lJr
VZ0t4obuyS1D5mcQgg+WjmSux3vpYTOOYBeo+q/86mhpP7bGaE3mx24ms0fCK/kvQ9ZNLgIUMV0Q
9aDgZPidE7T9zlMGr8pmyggi8D/QjWuf3UZu/emTvjwc6BclbIKxE7vGJyFwaffQQxGUNf3Exf+C
uUTDscHPWDlo9e7xEoxaRHMnZolTV1nQcsNXnSnKZYvTNXNJEhS+sogKyul/xnEaIGrUgqKM88EJ
2vjrTgtIL1/ty5cnUbv/pUdRyjPAggOEcQ4LKdHIrqcPDn0f0BiFlBWsL7QMsEWiHabP9VG8Z4vk
ZmBU0tk8VcMFrswQmBgXm3oB98TlhkaJLWAyUgHsRtGiizj1QVTqqL63Q5p8NOU8dZV1Q+QLt9CZ
7JftTAauJ3lr1ylUFnCQ6FM/GfSIMyIylPpV4nAs0shwf0mKJ3oM7ENmPX6WhlRZP8myvPOPOSjv
dTGReKDuH18bAW3YKXlD+hYr/3xCeKPSkZtt86jiskFCh7uPN7F13O8zxdCxobgZpXU7HqsDOLAz
tEeFiy/9ClhwiCklbiVudz63b2VJRp2/OpDL2/k+NcJEHktCNgAZQzFB1+fv4XTnGZgndJIN7poP
Y8bUcBEyUxuRQdP6HE1AZy3HIFU2v6cEeFWKDWbEjveTjFDGruBb+lpnwMxoCVl9Hbp3/W21q4MW
U/gJ+PoNYnB3t8BJiZgsXnSpPmfNQa13hT5tD44nA8/CFtc+PuCg/LERaCg4WmV5Bb9XMb/bKdvE
AKNf+LndI8cjJ+Rmy1pC6w4vqKWnxwb2rRYzhbJOtc8o9IwQyVUvYE1Y3yl+s7cIaHpyAlG+rXW6
oAIEJ4vb9XY5YxRvD10/WkwqdrofNK2znrUe7t8vhzqSv0vLapta3zVS0ZayMO4LI2BZboiCMaEN
6s9AAI7bu/zzqEJfuM//xLUYlBakH/2enszLOmp4W4v+b9LyzJ6xg6sbwVnTLGgwK2Snb1kn3g8X
TVf1MI0hJUEZjhKkBrsUkr+C4fO8D6a7CohVDT1Q34+LE0pOgLma93mmtrRjXPhexTAWHHYxGepa
Fb+FGvTyircoewc6APY8jifESMpHHLvoCzHXHGqMR1/Rs/HKW6+a8yqn2kkF1hvFUUB35Myc69Eu
s7C/G3EoweLZea9GSwGv57SWqtBb82OU3skri0j+GmeNFLI6ZPClRqj5qzDQ1wlZ04gI5+2q5qON
LNNMzMyKDLIQ+x2WWOKYwWl7XC8IcO1tffYthHXZaMY30RjlEzEOckSPzhJjd+oimLIQ8TrOrBQW
LLAGrWK9QfzttzxxzepE7iEBDNP2leH40wJt+mPzq4G3CjXsVvk5Eptt4OCck9cdB+qD2i87TyjW
37DXcs+59tJROa58iwk0/g1z1wgwLjhl0W3semZ063RCbigi4twTyoPOhT4Bf2cB6bwfN4/P271i
0xzRcb0PhdkK8BKeNa4k6TC8pHrljy1tSsTLTa81w0WiypDhu7PEIXv/riPoajmvQATWNSrxO2xr
K83dpW0u6BTz3iXy4Ufg4Md+Lx5VR8ONAcPOEXbxoUFTKloLqyhhKpJLc41BkBymcf/gRWpdW18m
d16bQXQFk+slGOyma88NSs/ETcGPit8US9TmL3cbzbR/Q07bn2A9bS8Md7LqY5d/UjuzzqefDxgn
dfysID1dShm1uGKaPTCGfEJyXF3Cte62XYZaQrOH+FpnCQIVzGz3pxY6XSr278/YNHLZMWSZx/GD
wmTBbt/7hGAqC74w3FT6YW8Dpzr0fBDb1errTjQ3P5thEAvG6LYTZj70RSmo7nqKVKVrd/Brouwh
zPiIi0KY3lroEBbCVjV/l+s1Jhqp0VgbYbYc2xc9G2M9DUYUn0O1sPIuvy4oNkw2XqCFtYRzVjFo
z6pWGyPabKe4Hd8NY3YQsFsuchrRzN17jo3wm+9dFNvunH3Vpk+0sSseqlKAVou99tf9H5jXw76z
5lM1nOYv26p0Y8hjW/NINUtxOx0DTusQwjh80bjjFQtgZ+Sakdnh4pphuHnaaxPIjxc84QLZhdPQ
eoHTWGIDW7NnYP0c6imnAB4c8W+z0TZ0iatIY1XBdNN1XkHCWQrycIee/Me0bi2jW17RW6KUGyEC
p7Ql1jPwdEU/mGcmbYPwvcYTvE5PXqW/YGFPZLpswyHPYd287pdGLI8e30u3jWb08J6F3tiKoEqC
8p/mZitflUqaGUr3/djyuTUIlgV1I+WbKFPAjyNicVnKJKNi2RiKud5W+JdFfP06XRfqzzSPJdRD
zLvxYidwnv7TwJ1MGnMVe8nhIbgIq2WRzDz/Q0cNeDZyKCwgSu3fjoPgSOlieQx4T6Z/ZDdp3s+g
wEWaP0QwxYU4FG8wtN2pzGA7kxlCY8nf2kSvF7K2zdJ/M2rsGQeTKnle5OR9XO6bNbYsN+TsHCBI
wzLmYdF/aDmIqGuMFkhOGtjTRjrC5lC7cVRkcKZLTIEqec9/w/MPdTyhAKUAYgf39vZ/1QJaU2bW
4L4j11Emgk3slkWYfSULj1u12NlFvlmy0bDdBd2ukW9YcdiSZ6RN6woLQY3Jskfj/U2u5mXv4LjW
FQx7b0Nx+PBDlAUqEjYOuLwYNEKXXxO4jOC/22QEzmyF/Js+g5N9y2SBDS4QQVqVjzVplt1z1vcB
k7puWRJ+teWaqjD5jNI70ZDo9L2CRMyMSQxcJL1fzb/ltnW3g97q6T0/tmoZc5XfgsRWq1vEwV6v
CFtqALVsHZpDe7FNuIopH8txIw+Bs7/rLwuzKrcOOSQy+blOhw9JmSMjvR1poE/RHX6rFx8rz/r4
D3eEQDBeuOR8pQcNqGF8JCMwyYssFwE4qZgNWsBdJecT8SAvjXrCpisIixDBP1SNDvKl4RmeXbv4
xVl9JiFPATkw0wJpAerJUocALBU5UlukH0zwDGCLRebod/2lOjubJteJUSRKnWdwfKiZbvUIwRNC
/7HLq/uk2qhw+n5Ojh26TA9BycJ4TLyGaO11vUT0mIgyVbAlp7dUo9GGZbNEmNBpwFpX2PVT4khs
DxddzyfmALXtG8FV1GoshxHtsHqWaIR9m4S2siZ3/EpedPMHTY8lpfa0CIjoCGflkzTpLnFaQN5z
WnU8TqwhdvnaNAEbkqzOWMeIXPv1aq07nExyPmd1j342ITgEJBK29D2X1F5ZkKWCwoIvc2Jrn2Ja
hUwj8FBWPN904z2hAI9/6BN2yR9ahji0GcxrWXBDVVWqsAF9neWVP5hLVKvzW1TExw/cn2n7Po7O
1Mzuy6BoKiA0lXBuUFBUuDCi0KGl8oY+OREhpFh2h1lMYz64jyurcei8zTbUWMJ0Y6uqlNFlo8xi
YiaWFdC0EOeH2VwxspU5jAZ8MsxP4LjMNdBRaCQGfTncfZAExVG/1J/bOzSm3YIbqxzLo9lOw9Sp
zDCD49X2aP29LikqJfMyZaoHfLNF3435aQJ+pt6KScvon5wYdVomUAoGz+nBxkQo9pd8qPiBqaWm
6ktG0MIMwpZ/wRN4325r9B2N4yTvSZOZoUvCCAVTMPOseyD8Z0C240F5h1e/DkabQsEghkUgfu9D
Pt6DTcN/HnbZGP5V1Bipr8biWu5NYIfnl16YbO5u0DELN/qod0lKGWW8nNMRLl29h6Z6e1Gmaa09
tUfw7GSZp/ncKZuqM9+LXhxlzrh/Sm6tlwY8+GAwHDrJcUKfoZ0lfnCZpBnoXtYK8dpJI22doGpX
HEVvcx7P/VMXHbRUauIY3H/04vou0As7wbkJi0bTMdhqcZR9lJtAkr3T0utzQL77AazpJA48qM9U
4T6MKtzAr1zmBrXgtYmmfHCG1IxQnhwoOYQhS3eMu2kuzmKBfjeysc2RVQGZ+YU0s37sjf0WNRG4
lZFNp64HXzZ8avvlmsr4r59vzgGkUF7rWESFvm5t2klthG9iL87rk/u+NaFkW6YSANhE/jEnZBIq
zI4U3qTZABLEWHXx5BPKDmZWilTvyybi3p18E9Vn0nlq6UIbwkoPlK1qUHhT5Mzjtzl4FM29HP14
2CuaLIEncVswR3PedKLZfo0+SEo4QRZSpX0CrUpcIYxIuzmqURT5qKwzjZ/YxLgA5us5VkLmRXOE
AtbZ8drlL6CuXR4dbUJQXWUckoIDm6ug6f3+I+8Chpztyv673Qt5+D8ElgZRfaYpPPRN1urDuThZ
/bcbxeSp/dZerUicbBSqSb3q13+M0NDheWsRfmEgdF90zyodO9tlSiJP2BF0Uq8lGGmEpoZuKv7o
a6Fl5WboMNKQe1bH+CSeV1HXetzQU+JY5NGXo6RWFlLyfAPw10aVLArgW1OdNwNLqvdCwQQH3P+f
yxGlo4nLHDxd5Ynx5WlnzpYAdo9jxHbeutz3zjRUZPwrsZwtGK0Ga2B7DKtHj5gZPQH7DVg7go61
XMt5nGEejDGQePP/p7C4WSYRpn2GBS6dRu33MvbFD9HohsyIBLZkhYPa7fDPH/ylyJGZHaWgmWSZ
wqjPFpnwohdPFKtuX9+DB470i+hBuVrGDlPT4eJI4YzaB4ejesa+95WQMiHEzQvnCso9hawChhcW
nQEYtz4MWW/HIk5QLWMtp9CBGp9M/aWjO+IaW7N3JNHBeINdZputL0jiStbSxbGi2+6T2PzbErd6
tQtT6U8Nhz3CZgmWSoJbmlrlJlZ8qUwCZIdxN00JEFP04HlZzmQXFckUzzCC+sfhH2UzF5oMuyQ3
ztZW8LsX2nSqbPApl/RBDuGNSavJnAXLvfaoqUu6lDGTJwkJs19FldtYYn8BIMk0Wu40YWlptHfL
d39GV3rlWQDS43oOfcp+4rCzsrK1lNPTTp4uTTDOPv4bFwYGKWxkR5K2k+DoV2g99kH9U62uc5Qh
4pBygjezYwRHHZenuHj5w2UZC72sU/t4O3Yi75bkKKapbQBubk7rKyH7UEiGHnHT8CKNnLgmUTSu
NUn3/rhjfDvm7V34n4a1WZE+a17O5qIPiX8WmxHqdJCwEey83tofDvPyx8gCJ1cRauhu9l3WeFrs
FptH2EY6jr0kWAh8MkfZL6mv6ZH6M64NZHv/8hqCbtmdLIwW0aifY+OpFY/rl6IYjkX6GcrAKVkx
SLbEjU6EIhlXzz/q1rPIVGMcAHmZegFhiiHZG2RlWcuCeS9yMjJ/qBQrmM1ygGgnJc5RerLsOfsA
CEJdzd3Er8xrhkDHQDo4VO9z8hCfshR4h8uqwffGOA1qmM4bBYY1kbjViQ0LrGp+ZHehUcHondXa
lDyFl3GxbnnvDjCS+VwHJU4/iSDK60UIH3zUB88FUmiL987OYq2sHaMzmStTDQg/7EKlZHEOlwJe
2CFTySA9cQr/HPualfbX05rzWvn/Jai7axZfdrOy5Hpul7DvjEV/fHN4+1txxBUvqLiOdu4XDqkn
vbxG0UHg0N2LEnT8wTy8knrzx8mr6DdltX4MgHjhcXImKw055a0jXNSJg7cD1hghP2MZnhJ/edX9
aHfm9+BD3W1BFlw0tBehS/SRKOAldTowOtzQlvZapaeZ8ORadGhChLDG5nYnvTsEunaqJdp9DSd5
VPXTleoZKGyOJkuGS6utZ518x39dtJOlgM0CdKh/ob6xs9hgwPsVgAJMXCALIFlCzBAmsqY74OoB
Y1CooP8kP6+P0/DhCK3ow8ofJLrIo8IibnEDtnN/yX0mjHM6Z+7CBvbM2Ee618WAG28gK3di1khe
DBjXwwHb0xU3Ahii4M7ZpavNDytUfp2L0Q1mlBdhHtqj5ATnqjvW5guOaWwyk2Ac+tmNeSWsg61O
DDwCdsgvSCvvfeZSRlbhwqnuPTikAIegbeUPFioYSaxSPnNEvxW+2XVNaI/uWuBGroJBdwnfS3pk
MNEkmWPAq8cinDc/TsLxoHZnQUH1R4whLaeEtZRrAdkSPkcbRh3ehSDKCu130YsAeKWr/TdbCf4U
Z512L4H7qvMZEInYmnQuY+aLJXQwrUL5qFRAiOHRWar8K2fIavlVqmdH6a1mFIrm9xDn5PI2+WiG
nLa0l1q5RuUCRugOBWpyrLFRInKXSe/RoJg0jDz7Xlm28PT+jHDBXUda8ga+66Rra/fh9zGejXzm
B1pfbrAHTzm7ITcC+8PcvbsZsDPZtzh2uKSpXKA3bZ7gwhtIhDNxhzubCXjB2LSbx3pdlMc0V1vO
7bMbRdTqlY+fJ0rvBrxoX0lAzCX1o7bWU1YD3jkhM0+7gK8Vz0z8SBAdkWe32jTjZPDbdu52m30Y
XhYdnEo+5OGCaL7yNAZ8Lu5VjKckdNPGUvDniA0AztlGmPjOxVEX6ZQ9wPrZzN+2wA77dTNGNqBk
UU4sR1p4OLO6XKJAPr+hQ7er6613sQj0s5QpmBCikutZZmXKTgG1NxASiiqUiAfu6WpUU/e/CSA/
d9kQJUvEIkSl3PaIfQiviobfdWKl2d/bOnZtfJzcRI3FIx+qxddpT0kx3VjGVJ/xqCGsYwq0Kdbq
RzNwA7mE0FMUgC+u+2wIjLvrp2bo9DegdFoLywvJT1j0VWO8SGIYFurZa6SJQfV6Qi9VjsoI5yrX
LfnPCDudjxIJDdnjjGd6imyooX80CUUJOiBhjjyMbS6xLotOLFApzF0NtYsVdnWJBa/12LDnCKhv
pNe+G0fiTG2i1Wu0i8CcO1uMm+yVbo/QssefBT9sCk7jymhUjiixAq0oea/vO7l4uCKR6vJIlqDb
e/tgZVl7NR8gwgkt/2lBsLUikJmmUHnwkrrnDibTLxy/2zV7f3mXavelWbPzJKNzmos9Y2KKMiXV
LkOMtQyHNIi6VeOZGQ1dC/Wyj+CFvhyMTAxjT1xa4lGBJI7M6Q2iZeXan6XRGBfgc6c71iL9it0S
JBuOgVcGFrAOLolzE5xx/nl52mNZaD0WaJ+7E6fN47IHP4SYfi0UnG7x0g4VHSl/yKUXxuz5WfL0
qj3NvdcXAvLZuMEEGYl58rXkBHatDo05WnB9rjCA6vgHv9zVKWChIKzMFQ/k7tgKqDYU3B4PDnag
xlFIyRRf5d797kuZTMjwSOkQmMtCV/A00yfqFUOt3OZXBgOZE16rGczx9LfK47jRHQBBGt12vKMg
KHP/35S2jRf2eZcHN/bmYq6r64qC6FSadWOjopvc1tVCDxQ4sNUb9fU58/U/tSFM4FuapJJRgIgG
kajas9yVJD1M58xIZfJkIA9EYeYIoV9ZBCk2j7Z4x5gixNYgLkCTAYCsE05nP4Hjsr0TsKES1DEx
8jd3h2HT14nLoEwGnJrw/GDUUIfF02iEIh5NgijCp8SjaPIrdvWoT35sFz9sp87OIM1uv06jjOJv
OuvknEjsRux27SMWqz83zGPyNo12en70YnTZNUachqrjSaQc+Y5eHyJX/c8XJu+x7+/Bs7EHdqNe
58k1o25V6Ag2tDxbhb9f4FXegxhmVtrdjuYkQ0ik5vyUL3KX/KC31liPG2MbZe8/HClJKk7kGnex
Sc6OJVpQ82/Odoh3HayQrT+ogbt1epjbuXZPRKIPhyzpH/1N5wXGYbSgi9NKmlcaL48Big86jqx5
5E/o2DU+WMgyWi8gZofxclZu54JBIxB5fI77b1zuFk4Mx6YgEnQzcbSqWfTtVOGxu39dF4L++icD
mnnDOjTMa/ikF3lUd/YOXtrIfGXmqCkipYHjImdT31Hwc9oMLKu5Lbu8Ey//6dGQmGcC1A26+Z2P
7h5lu7e8BNigXwqW+8LCSig/nIUWWPTHlTHgiYLU+fZVaz3KShCC80smR+Sl04/FAv5zvdQ5nG9p
5jeGxS0Q/BjEgYX+nPqoHx0s77ykrRhCKfkgGXriRHqukzhNs+4s4b4GmEAphsykOX1NAMXUhC9g
vPqHw6Wobv+xN4RQkUUUvx41qv50ydhjlpQCTYVcFEOude22xcwWp9WzGoqzH+c/1rB1LGNGeumm
F/JAyvbhvdaATChcXpG4nNZKuqHWasDzYMaQVOWYDRhfl50kLD8iWdPnhyH10IE7CF4IRzDwpPLl
h9afvpxhyEAT5lxCqdUzGPL1XbQAOe4u2iDQTt0drgjWb+3WAhqb9dMNBZzmvmXiUCTttany7xdh
oemooV1Ppewt6Q6T8nPTgvdRRiOjKiJOIkVaNkyoJsMc9hGZQjLpYpl8D7OthhaARyZWQmMYmcJ3
8uaaPiLe848HC6FOkQZVJyCbfgX28be0EMAZDJfbVOFxJoSjT88Ge8+AnFy0AzAIwoH5LLUUSMlq
0V2MTcQDtThpQRPqMPdpBvW21Uy3sooisuuHUzpktb7OyCtN136GyKK17coOaBUvnNFCpMH2U4UP
hMPk0Bh4lzDkNYT9J2CXedcmvIhBp+ZE2QT7sJDfQ5D8fr5AzCHBbN9mDOPurWyQpRh3NqgWr6PG
k01oYezw18lLUwKCEFOON9OrxyMJFEdKnnayoYZjK9dY6tYOF+M1/ldNRxrqwRETRa4aNmr3eS+U
WCt2xf7yNyOhCuNntA1WuYkjXi+72KkiX9fHVD5rtz4+QABj4rgwgov4ViWlRWR9DUT58nW8iG74
IBFZDQhyTSVDPvGpPkulab1e4+cuYxqxm0wEVGPyVyadMrWJHSyRWTcs0AKnBW9P0mCYPt2QS6+S
ptTe5d4sqz54Lt32N3K8P7V5frYsWNB6UWbDOcjh7fO1wk2xck8CEpgqqMKcFUv5k4iqT0uXLvj9
LgcLttRTU/git37upBYcXyOEy+PFSkYncy51SiZoDi0uJReyB+fIPiCIfnUwW8jqWTKc0ICuYf5z
iWcC9NtCK8f1P9d2chtpcjY0TVAN0Z9HdnNNPtT7vC5o0qXeifoY+i633eLzSL5nU66SSMjzOSv5
G0acVyCamT2Vcpx+wzVJrjNKSqUPtGNmHW4p4bdKaDZQGv7SXM/H1AT6Ug0APdEk/ZTXfjYAo+UW
dot8+cOtuSOwOXQXJwPvSWXeQmuq+iSbPg4BL4kpvsTHSlzJYPJPrtwbgb02Ombs0bc04c79DMCp
KMNiqdMJxNZbD1dokxCkS5LFLdB9ZN/qMy+2HeyUBHXQ3DXxaptFoWn5B+QuSu3NPSJ1dHMhq9iI
z8f5gn+epTkbUz9zWtJrVGgyKJmSmrYax206DSVXBSqq8R0WYaX+GM4Z02e2p9Tf/0iOndO6aHcm
Ks+Lfnpau2+USGWeVhlJxewEilqBcicc+q/2rtTW3KFzbG7fwh5cuE5bwpWScZxXXrUNUj4S0xw4
gJnKgFYeH7LboXm416gMTbxa5+s6OS67JExMEs15Dj5znRXnImqL2GJQ5W/17eV7rCbFaEQgJ2bs
cKmmiNKSDed3lMgTQYqXC4dQltseTM348j7koA+USIBAaljmaKOm7+YlmfZN6rBfwS3IXrKclU2y
LmlVu+IrR9I8+nhEMf/cVpf9yUhVQyqx4U7mZt8kwQhGvcfhYFXSvlPxcZOyCsk0FYWXrG77Be6E
keczMvwg9IVQ8OGALUcCjEUdApvjg3wAndtn9KppWMDSjtDB5H+bWiWn4sMjQZ8urKKxdkhsSb2a
FUVjP2La7oUfVkhaTJ/aVh29diiy7EWR1BgthgN7jdFlFryjCm/+5+VOStmKWEmxPVGAIhyPz+jO
Z1xFHzUY6Hre4g97aQbK9Qou+tsOiLlAqd2i6ru7CkKErKpVdhrhJolaKaXNB6n0x9NQAazX8pk7
MMVD9efOw6WkTg+DlKg228vEpcPI75l8RuUgWmbp7MT/RFTIk4g4eOoHGwoH9kpZjjXSTMCnvYng
ax73ZPxIYHx3NUAMr2J+GrL7JAW+wLtOib/HLzlh+nSVxT1Ihx56kI/LAbt+pW8CeLdUGPms45Mg
pcSigCmlZy7gZkVrZfZrbZNpflxa65RVDLyjey3TjEnEgJOxGM47Aig16K3Fo0us+VzoFv2jl4C+
Z9RQx9gXdoczUFJ/nQpA6IH070FycAx4w0eJslIhrB1i9U6xj0ojtYutpYO7aGFnC/w9Pt1VM2CS
ngCkmP+vQ8m9ALp2qPBPX98QBx3QlXZbulfkUT4hX4dUeSUC2ykT/hFt9u2Eq+pOAxZi+c8uJ3JS
VZ2fK8pCuanIwjogkuVqTD96bxoO9cP6p3CXivuYrE4zEYsgrJXrKWYhuNfAk65NR0jNjmBoPuop
8dZG7W0X7EXUXTqZnnFkGLCrb6lZukAEodOWXrvpeXPUkJx7usQUJaliWptmdK1Tg9q08bMdEV9+
u852O4eRWDuo83iz50Lz6KLh3Fb378yAbL9zznIBbn8fzHNWvOtknrIHKqbfZpYG41NtPbFL4bhW
8k4RPoseta43hIHgxQUiFyLIvxZNbtXZso8BTHS3WZSNggZTK/GL+vleVHLTGMBwXcLvq5oMPr53
+2Ghp69Z1ZvfVLGpqkgVuHUEqN1VWMRwRkba39EAp9OfqoBhzAEvG1bpVtiIFSEdSM/qmfqJh+7a
BnMpoWgoP6zTxQKYMSo4xqd76VImImuG5P9P62tp2ZatFuUwFppD6jHutENOD3zhXgVjuM6lC24/
JUG8Nawdrdi4p+O6hXzUNOfvJFNADfHQ2AICDgvJkBN3GD2ZYJrJBjBNaB1kz7pJMNH+ATg5Fv72
zGXmCVC9B/AwZAs5lRcILzI+nUnl2i+N5SYPGE4n3Oe3TatGcu8Xw0aAObXv/eQfpSRMwkV4zLOj
8Wap+cCkk1sDIa+t1V8yQwBu+ehqGI+xutJN9VsFuVMEhGMyvpE90zKFBcruE4gHGOQepYt74+nu
m1njZuHSe7skhVRJqOSq2M2diWCajxWs5W4FLziX/4mPtKIFOiOKqvwVIIYUEfN3IJkFq2xILV/F
awXtVORy3bGSR2W+HKRYCMCJG6Ctw3UOC1ldQil0Xb3JMK4djtFncPGhYdQqJNTn2S5FQAMlwIyr
3bWWqOjVv8JtrfvvTicpVwggr0NLfLpPloTPPiy513xoSEGzB+o1AG6JXfl9wsYxOSnPk1UD9oly
tz8sbxKAYDm4VD477YeadU30O8cGGAZCDJpV71mrlqH8/R1Uubf71l5a6ORb/5VHI/9XeUQTSIcx
uOKtlieCiHhw8ti28waszcp/YVcUC64kw2s171qVvkWl1fF95PJTpi66PhLen9XarmWizxg0o1GE
Xg358AUrHAQdJF6YQRJ9FbInsp5eY3m4dpo6lkdnUciPHcirPawpzwGLem8hyqAolZUcLEHkZBah
ppjdPjeJlndFh7YloCGm9rp5pPEK0y+SpZ5maCLxElZd0AA5hlf0E117CjuAadmLPkxa8T9Y7YlX
5xBsfxiMziftha+W1LUNpo/avreUMerMAKceYL+7j3THU9yp0shcFpV2mCk+ZjEkIhw3xb1Wg4Ol
e7B7luZ7SLrxkdb9+sCXg7VWc0kwsnBtzmQGWri35Aba1zuh1Gv0cXU0gnwAdcEPNJ80Bksxivrt
pBSwY23GNG1JN2LIjA25rfzKi2fNicSU4ZJLSJa3mHPyCd7SXUWybvnkRKjqemPicswyUytHgm6H
33H4Eyd/Axj26cAKiokeUk/2a5U/KEseLxM0KxMMWm2kNdOzhLT539cKUTgdgyng00ym+hRnlJAj
z0vVQxkbnG2QlhN24hxWdJti71IAzXoIyA5z/Iq7/GH3HMS18HhQOVUgjaQjUEbNuTMS9f40kFHT
FhLpsjleUxLIQ/Umqew6+zCrDa0gGZp1jbMLs3Iv1lPGhp15UB603Vzbr/pluQj+GfvoV5HHv7Gt
WRTgBZAC1VYKGcnUD9845FUnigaSqIFvOT64qrQ1/3OcV3foIVgCB+hquCZXckq+ZTQpROKG37MI
GKddNtZpV4yB8DZ1TbVy19X8OGqa9WHiVq6QuG0k3SQ0dn6GwgZNHeJRtT4zlpxgCNIIzc1dPdSu
tKVSXbo1i6Fad6Xis9KD7QM+Dus+0Jr77Hh6MYA4Dv2jLInmBWYc5eHt7+jjBl3Jhn9kYijqnXey
4xjiDGHUd85CuBqLJgpyKLJum2eJ2PzyuGq21UbHpPYqEPKt/nHcR4P11CB+ov9rB+YtEvZSM2pX
W4kfK2OpTbEo2n/kBbhO5dhkqHDGTklKhXTPw+/throQ2YQTBD0vgtouyGvvfdfT1DnN+2vO/yjw
xBiQCNYyp2qaX/qXzpxWSbzFD2GRPMT3GjMooAwomZqhTRNsCddEdekxYy3yF0SgcG2HEoOkTFNd
4SdKZd54oAdvZzVZTcTqVT8aojQ/Ms/0CPHTSjuJplGnZK7Llx85OPxESKWHUHUrfAkHAfpvYdH4
C1qDJpsUkEBKRRZH1KmxBhTX7qJZsAGMvJq1NsJ6/eq1LfLxB2az3ddDVvzN44M/dYLCQpqUbrjH
2KjOIEjB4ctGGXakDrsADgiGk42HYLL4X/uxTkQdrqTZTd5qr0QZvBm1v8ibIwJU3sTxic5zqi17
Aj6FJmN0i4wvfwaxXte/gv1FV3oSp2xMBWb+mTWgnior9PTCVUM2HJ35e3uH0hUBiEYij4Vd5uaP
iMK9o29PmB90212UI0GL3dOSVrVqW8HD+KYMxIftcM+4ZJ+5Z0nsTou86XFcD7Jeuptkc73bztbM
nB47PbgKI6bcuquiC05V3ibaxzEErPbTok4xL7xQh3QUbeDiQ2fHInYdT0k4RDBsueKLGD3JSK0i
+GaxztozWrBSh24j6WLV5ITX5cvkdtduFFd5Sm389S3RjOcAMtcIc1cwTRcYdu9vZC7LdqBg60KV
dTo5sVtGqWkILQ3LhKfBSioO4aZ9PyCqHn3I72JsUC9OGcbBscU/BehHd0NL4THgkY+JrDKpF4QM
XyK6MJsNzBGJT/MKujHPN9Lh1oijfkSmtDt9pfUEqXB7e/2y07DCcOl62tRlRzOiXOtJAyUDVNCp
h8c3WDYavEK3lVMhXSSknpY49Bikzm+fc6iE6UWdtw3nZgwOb8Zd/AePAZfYpEDw/cf7s2ZqXoDh
2CUpknmUoKPnkmKFBM7bhcdPcmJmnYigElGY1osKjl0LkkxxfR0bjWNY22wWESbm+jcUG1hsL2WW
LPfbKXEqS1Ond0jO+jPn8aVp2Mj8QF1qW9sg/Iln3zRw3+SIv8sQMask/9X4OuBfEcGDXwPCPd48
425f65y2h/37sgFaZNevs0bpoAYXTLorvvttXpsQGQnGL5kY7QTiIpnRneSrc0b00iKvawqXEgQd
0viLDBu8kjo+PxZBICWoIxABIuchhNWP3EzJrEcLIBGlThAVggNlwvhKqDTxVrfhu9y7+Rfa4Za4
RpLfYqFDy1Ox8ZCrTRjMSpY3vfw+w9myEXHDIWKdpsd8U+ouOchoWeKGIPywfngdIFfXAL3gPU51
bSrTE/VKJJ42pa7rHDiVcSu9+FVOPsBr+D6bNsluLxEL7URs/gixn4r2jxnpaecWlX9XQa7JsGCS
EI2TF3Y6v82841TNdciA2Jy7YFIFHu2QWb0F5bDilJQbIaA3zmq1/DY+lEOyG9kYTRy3opEdHecr
bFUnXXSWPdQ7DFO8zmB/ae/rr47ewEsGbreFbr02TKYjuQVyMZ4tz1mngP3ChRSsOSgPgIPJPGaK
OoQeGW/BSLyC3KIa8DKRN/QuFI+cw9qxZGd8clf0bDYLxV7P4qKs2kgYBh91O9kSJOinBoZnu8n2
JmfMf7q5L+LUvmZHXDu9GV+noyPV3pVCFfslGoSK4/mmUVYnilLit2dOV99gtMqr899Qr8mk29Iv
RYhWNuq2suf3kUy92SKbTTUjzpRYKmgk+t578TU2hufvDZvOV5NfkXuF3qahd8x8NQkvfGHV6D8O
C6WWA7AJbIqSpjhQ1XSSkIaCWGBmbBwcZd+Unw8y4UyrTfj+AJqA9DJ8s+ek+8KbPeuNq+FPtpzj
QJLftm8/jGhzXGSYjkn7oHl8EhKoNBQFHKhYkLeVGPkkmoTzDApIeMapqeJQvVG8MBBCf97a2Tlk
T4ZVP42u/xCwxUwnSsZM5E7JvY+7I6amaFU3KLGpPgbeW8jY3r6KXDVo/cquip4D0FWjnGyafJm3
zd9LbghkU65PCCqkNV6pkG+9FrHfJXs/xF2Jj0U+mGc3ev19Q2vrI14pCDyrbnT7P6ylWxZc/t85
dkKj1c/W18X8D+2sfVQ9O1xFxmd95z67suZLR8C+/UyJsIjDx/qjLBTINQT86rlhL/toEkiFMmvD
t+TnX1tpjba7q+4LhMQPUKUnsICdLbtoSk+DJBxuNlNG0il3gsG0zkf6xWlQYnGYvj8Fry2XOETu
MCSoXLHcU4DQxqboSXl8FTPzTsaLwvdFoBd4YmLWdA7WzR7Dey+XQJE503N/i2pgDEDy2jaGbxyE
6Y/SvCvbf1dHsaHIjQ2Szv26WhgWchVKcEcig1Get+b34ilngCiC6UDggSzur6V3o8MtT6SotaNF
CWjLAnU/JY+Ja8j4oKF4kYUbn9SNicGIr0aNgmlhiOtpJ5i7L5OFd+PChPR5fZKFBr/gfZH330EF
tcVMLMz6tuTq4usHQiIpaIRJ/Y2ZV0eOz58Kg6IyRF9eLFPbPBUjjp1RKYtq5EXstRd2lctgEjaZ
efqIQzEaEhXnHdMVf69rLo605DX6ClEtJA+fjQsdzFsQCQaJyThYcGYftEHGd04QjvuOqOZrYTHm
T7CTkC2JNsgbT5jTCgqPOvJPXpZ7JbqfZnbnmLBPTeNOKLnV0UjczLUNJaD+lZZpDPk598vzoqWh
qbRAWxPK7LD/xKKLtVQe5NfQsO5Bv/kPR5Yx89oRkGL25tV+f6cFMadbUgr+gJBcBDDDDwgwUMKU
iNug8nnMt91+G8R/BBaMCwKpXwnQz+aV/UK8HvL/Hct7mWoE820WLR9A4dtvK2ljVdRE0rHL3a1x
RaYXNahHbSWSwyYy70D39obsSxDS3kF8jiYA8O+wYFXuEP6fVMB2z3FUb+j9jmsDrEcrWctnOJGA
gH0h6rJ6mIxrbjM5pH2Ry/aKaCHbBsqxpG7MWNFYriR46PxRifkSJlLR7yt+4UOB9C5lI1uFES8D
+ho92cmDiT0OThveYhiZsIUxtl2Hr28enhVJaENzC+xtl2jQpQuGm/EV/dfrv2N0n9/ocq0LcS6E
+vnAg4K95PzGK/zCi+qZnHVhM92PEtUmfBhBXTb9oU5G6VJJD1suW1eX+U20wNccdlmawxI/l6CM
VwYQbriSEB0F9Lr45vaUJf3c9lpIxn+h9v9sL8+u6nMtDZqihPLZmIT0v6kEK/JpXK1ySTRoCgCp
eooIwMdjX2sQzdynBkk6aaWrMO2da+9ytmkrwdqMbNnUAvppjjci5ccGwwVuU+ZFC1i7zbKoMLU1
6FYkf5VRS6HBMrf00ROYP2tjuesi/bEwO6EoxjBYqsuozvKYizPHu10ubmbzYEO0CYPRE/sCuCKc
hm7QhxWAGvHa+6RTGaBAE72yihN2m+llthocGqKWQF/DkqUoqMyvIrqXLty1FpcF9p4NvXohX/++
zfVw378Fv7b9I2h3Kn1IEbqoyVTBsIc8DzHkkE8RR+8G5yjgUfMamME0lii4L3DNpczgl1xNKZs/
cy5S1wdZPLo/sy0kQyuJitWSbb1vyAipTdumh3e1F+nSYMPva5VFzMaWu7Ic9DBjS3sax3WUBuHn
5zDbtiJwSDuboQqp6FdIpHETreJcYJUUFA7jbr2IKoIPMYpGpzUw2F8N2sKxNAnIVVUlB0Obbjyu
e/xC3Onxz06krkkiPcF8itZvLLmU6R5NDZj1cc9nsMBbfn4d1PdZbU+bozrJY/mGl/a8E4lG4YI3
UGHcpUqwyNXt82zyJsOcpA0vzHOYnFE2hOne7yzWudJcURRXaFFftSRQu7NC7zPRO9sNcf9s00+0
pq/ZbQZ08QBTXcT7M9kesS9mr8drqhASd9eRy8PXGRggKgLGEK1ap4QhD2YBO0uhuVoepvs0ubNW
uCFQ/Q+0v4wcHeIcTDRxx3TmOaHOSJfJi9cwk2+lBhnwHVwR+8nICFUxY8qTYKPDC7FIgfSZUT1s
GzmjHwKsbARr9Mf0Im1YxBD5vDV+DK9nD7Is4AgWbXdqUS+h2s054HPTBI5sdGaujlc6xr7LENvW
+Tcc3ARZLlz8Vu3df2FYTI5XdEIbF+QuNnzRtjil01jIQ4bdTU446zQzajn59Dnmh7veZaMpxlAN
nQrRXZvzBwDn3Clpa7bg5blCpwgNH+zEW9PRH5GRNqIUmU8DsaHoDDRCwPw7SLtVN6/UArUkyieg
DJ3X9qN016XU1z2B1oOvjofRCpCwDvK5H3JuAhVqP7z6vOMpk6aO43OE2UbuErwo+EGLd/kwMLSZ
/3g8Z8+P5+DR1NWHGNLZgWku/yArMa5ETkmXuJ6qpro6GT+hWMSjVGplELdmQsXZoWZN+uJchJjt
vcQMXCQsr8MhFvnHApspSOwtFzeW5RKlFLReSAGnJhrVB4A1+Cq/zlAfyF6lOe6eyENwBtUtnWXA
AydsBFsF+0drwXfSJ5WJM0VM3enkjyEvr5Fs/szV856T0SojuR79OiUZJaDJVXwzAPYSbmFZ/KAB
hqxapUw3ZdFTt6YGoHrUvcSqfhyCTdIHsnSqud5fH9aG74SkKlTSaTULJHK3frukcmwv95VVfMUn
gDLX4SIsvjTKFa1l8PCpYM0TLomuR7JLIrdzvSUcQ5oRqb1CbcUf/dQs/bEuia+49NdeNsC0HyWu
aqJUTZQonB/dvTYsiffJhK7rRK96rUaTv1JxiK02JcnOrSX+Zz0l76JAtAG7CqXs3JWp4M7IZ8+g
DFvb22tR8zogSDfz6te8ieclX8FOXwGIcncprtvHmRbtcGfXI2voC2vlzKfx8SkaJqovqXcT3tp8
sMHOI8e8gn29LKJEF2RqRgSNgW1F/DeTziq+heAH5BFVGkhyhAC1vxW0hO7e3/pRUrNgkqlPC7HA
Pp1sIg36EwJp0P6R8eTVWW3zV4+f6UjaYxMIl+nhHjBwKAfc65IbwLSZgrQ4vjZXpmEZ1B0khX8F
NJiyxGyi1jeY//uqr5i5Nj/SBBaSr+0s2Car06WMNx2xCLR5mi7zSBTieTTnTR1c2kIvtvXH/j6R
5A5+Hs5D8e5iBDKuq9wi7nyg0nZqBXORcP7MULbaMYfzKXqQSvbUKyMFF560aqbD4kScWIvTMULX
UqzBQlXpbKK++B1gppiJgLEO6107wmrG6uMeP2huBdyfkSP6kJfXZOXk4mD/HcuYrlw22p4sOxG9
0nL5e8zHooRL27J8VipZLOSJf7C5TKB0I3D+vcwC2alsAUgntMjiPYhqfjC79bek9NYS/dfTvmsX
Wl+b8KwIf5e1xfQZVWOz4/N5/ht8NvLI9QoBLU5/z3YDpf82V4lSPXtdrOJ7MCfpyJ0numzWHNBe
kfverWcw32EP9tg2gsOZRC6NsNxwryNwwhKPPhu1JY6W3kS8sUA7kG+NgOMydhlIihfjsB/hdPbC
t2K8AQ/b4wd5m6DrfEQbsRZwr8BwJxGiH6x9rtHmoL/wKqbJ27ODg9VYezZwsY2A/AASJysBrM3K
Zt8Dz7CbzcAsw9/f+B2b7FGWTgEvqWxi4/tPs3XGTzCBd6c+Coa9ILjnE5Y3wWRCn/VMG2SIWveE
HEQETlORdGJOIarXF2Z6tuZrGELCUMEN/XkPnxWjo5qhqk0cd+qKg7fnXMwYb6H8mSSDPdLhva4k
Zg+fTJdzgWoLy7pkfK88DCzo01aoMwxfO53laXU9BXO3d8qShJojLTNMzCkSiTEmWnTqfM7dawa4
nrlQqj0490i7dkuM6CSNyfiQTQOkPMOXe6hhshWTauHMH2+pCVMUfflDsQ3O6KVeg6nEJBIZLuht
5MvWPiSpCAYJEyLLqWxJAXrZailxpILNsDVEtC68Diaoi+ureQkTF0gI6dDRAPPI10tHteyj6mGw
Y5bm6lZKFDDU0jOXv/3SD5Dd51Lsdda5AUIJ953rC1fMKKSAlUM0g4LvJoht1NiKjL4VVBW/ii1V
ZcIyno0yN/SbVtTtpsa8cqCff2zNjDbobHIHSJiHtyU6vFDuciix4U3dUfVBv2tlTWi7wRnhdyw1
kTWd6B5fdmWQAXFjTdI5ZdoIAVvmE68AmIw9nZ+3+uvQKk6ZJtx7kbaznFqCQk0HxmKuj3nqX+Qz
zeKFhFtVGu2V4+qxQl9sESp3XIMtBqTcYCVBJQIHYN0jhI5eJiXgcW9Q/3Sv3hDmUBbMOxvMthhc
hGNROVbMvx99X63GH3jxrjxApN7NSNOupSbrWRQ8W3i0uEbUzixAKMUMCeBNtTKBCUSt+kJ86nEJ
Kr6A2fFYmn07kqc7wQ+IRnsIVVmJlnPHwJL3FPORyPcWm3jNAkky9cR4OHsfp7yBKpaFAJo4i2H7
3g7O7hb/st26vt5K1CqxqiUS86zInmqOQ/j3n9BkYoiJhZjtIRebN3BGRiK+tYlXlKg+B6jPH7Ks
2ay17BSc166uVfo3SSItUxbKd6B8oOdiW6iIxfWbxT95lc96xy1j+1bCIhDPyZqQsEQ2vbedF1S2
VJGsxY60LRrDWfv5s+TRFXqQp9e9WtwclpT1ytC2W/Pr1XWZVwBJo+HFWpRsnuDPrd2nLil4xnYL
0t3IU0LEh/q4kjLEMBnDU9+0mxLXMtgbTsM87ms6BCt8WBJg9ZpdRZUSbS1cjcZnPYkDlomzdBWP
MV3Ptao7/B3+HgWyRpFGG1flE2S63RQDcWiKYvSqlXcYKPkD2Jhx2SxMzHtUgUin5xvaMPXf4YNG
9SkjdoP/U8Z8jKsiVGKOZEPlB4N5Nlk4YFZpNNNBaczjUlUJnTGBzZcAnf+QLIdndQHwEfICnoGs
+v0uvAjrqX9wRbhxYRa6yIoNg6u3dt16LBQFj0t5tR4pfX+EoR7viu+7aNj1yz/k8DEKjNzS0uiD
GWwXURzuwIOTZlr/K9nyWjsB2sPrKNZ7dRmVHxHC/oDl9BBqgOhRCuGZob5c7rJAs6J+eBdE6I88
XkdHwp0155nWEl+ggC9sQjBNVF+1HmVfFwLdXJ8nKy+DxETq3cLOCocacc7U0bctHg7tlL3/vGZu
0tBTwLGN7jHTe2wqaoY1208MonqGgASJTfh7j5wkxAcIRWUhfy+skVwyoo37jdC9k1H6FXx40TuO
4iV8JheJkk2djU/vtsG1XLbXY5pfl5h3hHVLmkVq92L0rOXn/uriPAfvzKMb2euCycRM3L3Rlq8Y
/m45YO7JomvY2fgHstvlDcT4oJewWB8nbfI0NdAFZQ8jDCSCbtvC9ybIdzDXNOfUngRlxQO+/BLE
/1jLgMEHfTm0QwCP4m6peMSwKVjEXnjmjzBDkSqobDfkMBC9s9EjLASSQfiXyUhbtNRCJAZ3D2Vv
2f18woSDmfto3joXb0hakTQyjCYxSZreT45hjGjwKRl3IQPxr+qXv9tpF9XFEeImE94kZ8JIqS0d
w2JwNwYnTlACJ2KaWwGGcXWpj4X4Jl/dYDZhroJ5zyAoU4NoPry58wCHkfwJDIOzXBbUjznV/GG5
H99e1m/VUVPPUCe1u5V8OMGK9mZA8PZPfpYDLOoXyhFbVjp19FvNiO7vn+PNLJ6AAqdc91pJq9Sl
tAzqb/d/gJJ0y6r5ONFA7Uny/t43UsggCfPCqrD+GA2belXTpNgfSiQiLnr+GS8BiXDq2Qgqhsuq
K1MwhYEgkpPi+iZ1ZBGdCfCcisZz30JKdDUKJPuWwNwby58U0jpFgC7Dd/G/L8fq0N5icHvM+ERs
4U0hxZhqrXDg1N8sktIYp0DgJYH8EJT3P1oOEexTyhOHaEFNSg8pUPmNrpGS1Dh3EmQd8MHFYuKd
uoConqkVlsAKnQ9q2t5Ve6Q73A/JllM6m8ryL/LYocs2aLDsQxTcXqXJaG4GWPf2aNrAVKkHUz8f
PxAv37xsXhIkILUmEuwBKkbQZ1r6OIgS6QIuQlkSjGr6Z4MG2pR+T25xd4IJYEweeanUMcfN+6+V
C3D3W6OyCbGUxvSo0C+IffLIiT+iRaSuaqLkmUYQsv0rhdE40E0cxHLmBkWhhGW7req1VJuFW5NK
HOCU7qB8GCZ6Vm+2po+R3tSqvbLpMWaNKW2O5njskl/qkbGj3OWEzAlJNXuKJ75y8Cm+96lFMDEo
f1OX5jZXDu1SUM7Nuto/8/hKx5V2KaX0qkWFv74sH+9At9mNontHmrU6E7oc4UbyYoxYfpR/QJZo
dew2bVKWrk8dBIkMr0GVeF68kBLVXQN+u6CjqUm2T1sNNL43079UC4fe2Mc0FZhcx8/2jotcNhTP
52m+S5pOVZ+HbIcK/wkePJ8NfLBH3vq/AcJLjLqz1QQxLHu2FG/PI1eiENO8jpEWnxFn3p8X+A97
akoKv9qclv7ghWqybc6osJeqXgDGoVLoNEcO2tJXSICSAiTlpwyrYONgm25fPbEcc42+PnrGTzrG
ppcwkbiSMKRPMEPaELvPJXPFEThlAe0rZAspLMKs0OCpWiwgUNDuTvYOpQI08HUTEaDEbfwnzmiw
nAtlVjVNhy+D6yuAz/OTmaChmBYne7QQ98LPs1PRp0Wi11qu2MR4NoXpLoAAfe3iDkIV2XYLHjX2
QMk31AvcAtyc4dmQIAPNzA1zEEN4FCfkYP8v1BMPT4szv+yC8o4ggQYR0AQxF2yJOBqoLNpQn90b
I3FEP7i/V8/Qk/Ym4l0p9qX1NceR2oTEach6XMbnmS/KGU2b35l47zTe5Ed/vZaavn7RLtq8o4A0
eaA4oV/HIODrexCsfFjyb0nheLfRTNStAtXpqw6jEVJOtMZ9vD2S4J4XT4dOuTWjgtjY81WGaL0k
en8gfsYuwNhltJ0ZfRYqgjqzU2S0+jon5lmidnr4lnKEdDxGhRKh8+u9SCu69V9jKxSAcbgDm01M
PoFm9Pg2tpJatpheCnN2ywwzvxLSlhVj4W85JGTOAp1JUKjj/f1BraIw8M6sflq6lGJjHbq3aawZ
a27ZAd4+gwqDy81mEEpP+uk7x+pJgSFUEE2k8t1WYPkpNubowlL/NCZ1UIh2vJymVdE04R7jyv/i
TiHa5IVu1oQswg93riW7tsXpUs1GpU/NCTMJFIW5/AeQTwPYVVLbpC61+gKQgSukzeB5pQwPSe82
AOpR2lmRJD08OK/i137HXB3YBnYe/LkQD6RhN/7/Af0iPKQ9s9z35HDRHIkWmCEegL6vjdJRib1z
px2i9GKbQX/2Nu17klNH5Q383FApGPEORWxDmxG/uOrxNCsFwnGT2v+n9l9iW4s+pB66seIqndor
Jg0t3T6p4JN4UDG8VJf2omaXmKXOU+gvD4d2dNUm9pf1GnFgOdyduBD9IkCTFm40mwlJEIBWE/Fu
YcDhP+5tkG5aL/F+BZxeZiP1Deqcpc8CeB1G+2Cvj0quvSgaCo3/JrYMX3Od/m2paVw/0xlK9rkZ
mmo93chXIEU2ROyxKRgOPLQoW8FoAw7ZJc4MQQciL+yHJ7GnZyowSNmiavya+Ls71p08//0PRGSQ
SsjdIQ/RrH8eVxjOYfx2QyWGBk/FqnuyaAww7Du3pYadCSYjVPM5RWnCXSpGbtzWovFlNE5n6jNw
QwHcxgBBKCdp1NQ8BrPOdnJIAmQNAfR0O8az7o8iPt5YwmjlRDcxYUERZYVmJAj24PgzgHe9aynQ
Tzlyx+0BzltXO/paiFB6w/AGUAE8TuoXSo8TH+Rf5AmzkKXM+5Zz/1PEMfDY7XSLFwYNwFVFVyhG
LpDSDxbL5wgCtfm1LEHWJ3Ujk6/9v8WiBEdIm+nfvql/yzZsGy1Po7oTSH4pPxrB3W8pjFb9mURx
Lzoi7WeiKjKQrIXzVXVbGJ+iveNmWwYQobKsB6JKYveI3mzet7VxBLshm0WIhHw/4LO7JCLZsG10
ZYCuCMO4LNs6WqxCBpTuhM0QqClSGkBscwGheAI5Myjz8091jHWqF8nT1EjOdfp9QFPjlrSN7gTQ
ynC1/Dhfb8h5HQI7xBg0RxAQRrUBBW4SqFvHoYt/MCkEndC2lsTwqjXjmb/PdJqfrVv+VdKxYa3P
JwXBd/2gFU1K2jYEJenzRJLrjdGuOQCI2AA0J7QVT8A00QJkd7PG5q/0/jVNRH8Q/CH2+b8FD9y2
GPgpfdb7+LWr03sin+JfFiK6Z9liRpzXf2TnJDS6GFNeY2sH7sC6rKLOS//XkqzRNx26mhfbkWbU
YnoNv5ktAIj6+dk9uScwbGox1ZhNGQgxQ1R3Anq56e9ntS0w4i1RtOyLZhpyQhatFcYOGrocQawV
b63OIBqoxpqpVh+vitTeL2wyQ39Sj4kyAOGQtE1JaJy7kt0gUkG7VI/kGLjNR39FaXR+cOU/Kb6N
ZUS4V0GkdHU/plSN5NMEyK514Dijktd3QLibaP6Ba88lE6qPTHBGcS0VyNJTytX7//ZE3Zc2PMQC
MMuA8JRVbOkOVkF50uJjs2m6tO3NRP7YLK/TXrbR6aK/S7tsv7ALDrXqE0bR9SXsEYjMAu4HhV1s
NcARL0K8oGhW2e/vFy+Hw8P6Dk4FP27AUhapCJLCflp8shbBUxWtDK9xVgTOh+iAOKBAsLVVGD0b
zpLP179AF0vX1NwqzFw+rkJuuWdx7Sjsy/ZMEmX07+EMkD9w8db9+KTEmuu0qdtzBmNfe33QNwZV
PodOyzq5tlRS+kVxWvIl6I8ZuiTNSTM6NB3V4rbIlcg594sg9Exs3Z6nVadieEZGJ1Mbf60FX7c1
qPBA6zAQJEoU/2JAd/jpne/gIX70SefHNNmxMFiuoqprDhmXMf5PDMF6ftdpiDDdW1mDYFpc2XnE
Ywe/IP1cZgpngy48r+rhMEEXvJXKotPxlJ2j7hf5RXpSS0jhd83C5hSRoMWtav4rCO9M/lvFuutM
iJ28FG0K++aRJgtI1IiwjJ8kYhoKYKGaoAnyF77PSDsPd6EsFhBqk1AkFrdOtMYFVjv2KrQ2hiWT
YNPUlRrjWU6CUUKFAmFNUHJdE57K3vgAuHpzF3CPy9AByXdJb/A1rY2hR60Kp9JWmmi2qOih/jRh
z5wncfVjIhDCeXHzdnTdX1jVR5NrjRJU/YPEfRaV3+jZSpt3Bw4Dvnd4B2bPbwE2OifpJ9MB0cyv
JEHkZtljvKmlUduD1mtMhIAC2186ofH0x3P4JMY/icuy+wjFf5bmdhkc4Ld7MHot8K/bK7wx8Q+d
svwdxdHRITbZi5Mxx3IGC0B3S/tw1KwgBdYLVrZpjUORjJLKzcu1Brk7KE6G8zl0KQVsJDQojZiU
v2M21m+8QVyHS07L9VfjuFcqtJEyCZugKMuGOA1yQkKhkeoBi7aCfCl2PQG+jz2vOBJBAdl4pONZ
sAqMgY4EyI8qCn/ApP+CRbY/sWVbAtO+7g4ZgdEavJSk01bxJqgFon3wnBkmT+8qJQuvOvv/fdQ9
0Zktd94v5ZGQp6aDfz+wPkfy+mVKegKbbBQsGJJ0ubVbdi2Jf9skBzHtR6Q4pPctwLE1Vb2GdATl
jqLHA8yrqWn1w7puomfZO1evKHfrcdhGkIEdjDrGbZeXnqu5CvM3VoM7ZPXzmF2SkF/4qmJPe/Tg
x3C4vVxX2HiANxxU7znWw2XcE3aH1X1WdIoh0pTYWGxoVs//eJGQQrynXWbsrAv8n1L2kf8bP65X
iTrMZT27VUMxGlAPneF9+fvgdRi9k43E9hejhwYhfwv0Af+MY4XQw4ZvbHBDOM7wvyVyTe7A6vnC
FpmC8RwqKXtB9/tMfe0Pmdjrjhtr+6RsF5hrBrrhK0DYC1q2/Z+2GxD+vqNTWRzxqOJRMiOiEJ90
0uNCROEO//1nqKbgUJCs1rOYi/AQgcUy7Gv3xwmiRuCi431T4AabizjU4D1Ywr9Ic3yNuwv18YU3
XELiKBI+cZEBkIpsj4SolLiIrdkiSxafN7trXKQm23Rh3MI5wY6qpWHStY6KKrPCIwC3hUnM0ve3
MQ+fSn99AafdBz2eS5YPlPxoD3rMHEmaLbpW/xe7XYTX7hNZouG5Dlc8O4JTBJg7jLy2UXsEw046
ZMFR22PjdCiBnXudvVcJI5PiN6Tn0F6FDeQt9UED9HmfvOF+4/meZmQMEQVa/5CsCwH8QKFI5jgY
ZyT3GsfrmpptwrcL+o6GFEoL0TbjgrgxIp5KJBmeSaFrhf0NrJmp71tEdQlb1yT1OtXGqsFy3VPn
sAW2/c5lKpKNNYuv8Ib2z3XswRjTQPOm2mLo5nMnVc9cFSEQst34VDu+mOcLyxVWAwVhW0/7Mo6W
h1mtXz6q25Kiyhi1RkTu6vDiIxy4/K2qV061/qKJqP5B2iEpFI1pDoUZyXLNB7iadvD7aMFA72v8
JvMxiLyOpEdOEzQ6nTF0OSv4w1C8pX4KAAGO+CLO9K0aG9pRknEKVqlTr98tCzF3H8L0LU6cOEzu
5MRlB9q71a1po3yVpkBbP+OR+YLmH7pHqwkqPMbJOv6czH+l8vmE6z4ne2C/LuqEYDMb5sNrlIkZ
nrzBlz8FSdVuThslPue9+KkOgZh8+/L+xS3Viha/wU6rY3ixOp0U6+53pqm3t4h8sJbQKeSjtiV2
IidLd5L+XUZwaFp0xQsYfhAcCld/ETv05Y51VRjs6h3g9+N8elxhp9Xuf0IfncXq/u6CZ0wKv3Lb
O0ow2JdQ6t/9n7sTQvdSCC8S9Jq4AU8NwZnjjnFqjD8UXOI5b/l48Kr5LOB92ZcCAR6mpl6l2ilL
vteAONs+7m61Q7HHMXAen+Q5IMmG0GGMNQLIIxP/ONPF89vv0Mn5jIyCptMRYit0o3SxW8cF67hZ
8FUnxB0+0RGyTdbPpjsYwTb7hNx6zUmf/TlTscWnX1J02C0mHClSlVdAqcU1tISFwXaa2ZUS0qrL
Fat+gCzloNe1dI9V5/+64DJ5zFu0wezwM6JI9ssJmHTsG/eTRTI+PfEOqh+PfFVR7oWI+Q9edpij
kPOsTxQvCCK0pZwYvJSjoKCzw1HPb0hieRArPxaLWtFO8TCneGcVtTPCaQKyTV9DGTuIEv9/MQfc
AoBApdxyCua3HK9byzWzf45J2VZ9SzKcoPOMAtHaBFQtSV05hTI2MzjQ49rcukByzrWg9SLmMDMF
6LdPuB12MvicRqr3tjR0xMY0ZzqIJUsTy7/9HWB19E9osyHdSq7KKZxwzC6857YeQO0o4wLeGXuL
u5EUQuQiqWW+VtX2nFyDVHC7zJC1wfFPOeZF20/xR0Dep575oKOgID+RerArwIrWRh7GUR2T1MA/
IIwXGuJvce3rqrNK0wFXT8zhA7BoQmVNqP+EzpT1SLi96oVlH1ySw7kJVukU3QBRrg/fcFRehpJZ
fLDWYaNZiuPGLWOh8GyH4nSFpFsMbUWaQIGfDbk/9Gm5i5ryy+A3yZaouLb+hsrVIFCq5nOo8FvH
ewi4CCLF1+rMyU0Ti4B1E6XcJv5UinBLreR89Ax5ht0JUI8iwYfuhPoj0fFcphAPdpIVG4Xqhjw4
Hy9r1WfkQRVWMnVF8gG8I1KHZVsa5HA0ObMAC6gH8MKyWKSxSjjjYcVIpGudiF6kfD3OcA1Bb2V0
C/8saTgEPQ7M6HBHRsiFqU1ntr+1Vnqp2s2SEhob0si96znjmb1OeTPoyaxhsA1R1dbMND/L24ab
LF0D2uhlJJ/z34dWRvtvr0zSszylU8kPba5ds+Wg6QJ+YfldOT47BczC6+N+fQ9ekzg7g513umGS
wHd4t+i9qTHQjaTOzQE5BbuOGXJLlzk+Ew7GR0uJ2n7MBrcKzj+6SyOKrsi9WQ7yxNa6cwjUvCF1
tNIFH/trPseCysJgEqj1J7BA5PJc1VZ1tbyeTN+BP9Ly0lCJrPFynvWqXW62dExsUeaeU1+7eb/f
YFv8kWO2dXcqFTOpyegBRb/+AQuLLWhFai6IHWFEmpQtx74Eia+XSwIGscRzlj41chzbCWKNE4aM
Rl6HZKncvPfanJdfrbduLhtT0B+1K9nv/Aev1k9xMt8MvmQZSigWlqwneFDJtkDFbS0kLXvJTcC1
VcWxFilvgxFcPmFSbtRx/h+34QORW0n6zAGd4c6dCVQ0TVAoOQr190XaFEXBkqdSUdCqBhPeWxFC
b9QcW5813b2mA3eIpeZ9ZEFByyYt09GntpeZTQ/ZXLmAngl4JOhwLLAWhB55N2lsUkGH991o3EJf
eVtcX4UF90GIxIEvX/PGZLsS56bAhqW6WcoxZiuQ1yQuvod7zs7Ajl9V3p+7DErqBXSTBrvbO9F1
yw/i0Lwhbnc2wq1DfxnIp2D7vOq0XIMgsOFuQVvkJKBEhGTWI8JQN9ZrV+zMDa5vvfNuyf+px9u7
u4buJWTiEfnqE5oH7Y2Nmg3fnxPNEkL9V5QegqRxE1wd7vd0TcJyJ14LLnJmSIoT3T3Swh/065SW
D47kWGKcJucrN/Lhhr+oJ3UAH6zzZ3czf1nKgVtFdaKp5YLzZnBCHpbFE7TsE6eCMKlrttaNZqcm
MFVUR1fC56/1icAOTiiZUvtfxoWWatSZ8PA7PSnFHOYdifnhIWkGz6lUAp2ADHglMlZrLOKCYe/f
s0RFH4f5N8bEm1lDQYyJ0MO6ba8FnJZl8SoEBvtP6jcq0Ve+DmGffa3vLUS+DgchurZEHH+8e0/G
zEnYWOYMfSYeJVVzbrGgz6rk7JtmHt8bQhz7xrtmPhSQDXCyj/GlHzt+9jl3zPtvyHiz8Gpq0Wt5
FxCVfA9sl6An4/iqP09QzA3FY94X71hP6i97pkpZadecCeF050LqCkq3Sme4hJYedy+ryVpIOW7i
WN85smkHn3gInCQqMD4jh66U4WhWG1lZQ8lyvY5U+OOFXUuyGEoca8kpZHhr/1fOA1QAILyyyZA0
lnBw/r/qVPf5XyWldnQO3L5U1N0Cbc8WiSdh/6JzL0HDf1cTz/bPjqQXBL4nmakCpw9e4JD9VzZR
5O5G27+iaipJGN0SRoRPu2BLuzeJ8bldHXF7irIzoYKrMPg3bcE0bG/h/kg9124sPB2LeCzbJvjf
XrtZLyVAvGesXML/4xa/YX9qiwY+7eYNMSh2kZUrpBPh/lDok9o+Akar5m86PXY+3gfMxVWJjBwm
kV5NqxhtGTmoWl1PMtP44ZgUFGdAd49g5GdTDnHzaKDbnNhW+5GYuq7L4j3l+HNZtPlDn6hkQ3lT
c6eTlXUeVBQPMFU2Pgsm/s+77PXUaV2iAgvwP4NPMBfIBOxKV68ookdQbj3p++PVUHgZLMDTLWl4
p4V6sbhKA9MIgq+5DAYVjn3InvuafSmHsfRDlv6FBpfvGER0wQhHAVplrPzKm0C0QqQabKkcDs+h
DzoO8H6aygI2pudXahmujF4fzD606Y9dQ1kOqEhGksmLrB/sAElQEd2v9G4POYupZw07gURjlKTy
BGVuI+/TpCBDE5MBl+Vmz9/1WHReb4yiVsIyTBOccc/92cIYCgky+XUSMqnimSEWAz8Bnd/pA6pB
UzlpeyJRl/q2GB0+3ihVT9udjWYq2Sz1uy1D1E6uLUeXqwkTn0ZF17ydSfDXp6ezAY/YtA1p3oX7
zIEnTus46f0PqxFRNy9ns6I8uZ0jEvjJlAhSCRIiHejHQDJk3OhvJ3UkmjoO0QDErofbWlvozJUu
525xmg0V9YouYMsqkEyzWtrgjuOWqODngUFW/lwdAyc4S88JgRYXFevs0VWM93gKXSX8kR5OAI8G
nV0HclJeLn/QP+GYQ5AE9G06o/Q8GRdyKDdTPEquvyUuG4Ykf4tv2qkHLiwJIxb/XWBpAzToJtUs
3RUXa/CvmANnRlqdNiY+CGfidEJCEoashWyiW/XzfDAvyWkB09imvAbvKkKDTK4r/4kMUQVesThI
tGxstP+WaLh/xFttHrZiNKYp/5+NyRnS+qXg9HfNDoWXP1ny03rBaRZDJ+HJ8gV866ymiijT9U/F
fa4eVnet3WZOmKkAzB0GhO1qSBD89fnmYUmZFJmdwWFnDITZ5K3llIq8sTERyx5SRyijGKzS2X5u
1D74bMW56svSoPLzT5VICHr14O48g+qV1ttmiCTU4mHPlLjOP/DfmGGTPlIwkmEzXoXKr7krmf2f
ZN3+EOJd9qHriwP+zv2bFOQKhJudLBpkSA6LSMpBZMm0dMU23PHTyLgIXl3TtFmK0Wv2UmJ3r0HE
/q5eEiwdrfXIyxe4i6/66c1yci4XJTIWKDTkIs3UdGoYLfAjLC+QxUYAo+kpcCFon8Td3KIyKX2O
dqrVpXTGL8yDakOkHf+dUyx5GAPQTrdSl567I/5EGtyQqmFTVjIN+d69NhcC1B5icaMWQMNXWOy+
JN4fX5F66+Xvrq6a6HII2nfIjS8ZnzMobyxBZ/ceIAOklo4XIgKfNZhox/0UENntWATjH8anCp5q
Pouh/8vL+hess2eutoGdVSGHGXdhh0qFwtAPYA8ArN+VTQY6Re47/0yyXUyc1QpZysmZBMDwCkEU
gUK66Ojxsq3rmoRyfeZk2/NXP72xvFG+NfUSb3IJhUp+sWDWof+nCPz3miCOV3fjcu8o4pzCWh5B
00qJQhurOlhqxL9g5gtPnX9L3nzNRscH/Fd8o1kSt7a/f1uTW2fnsmjummxmBvc6MrtqemFxy4OS
fcftulqtLjsm918Fh5kS5qhuUIpRH5Y52O+2xiQWRWol6RLlJE4Gvr/NqX/0uPntN80//ol1I/IK
1wUP8RR/aEJOskrCnJbScxOIunYvbdC6dgsKNroOrmZxYLZ+Vt8xTesXF56I3d1lDFY04Kly2/6J
sW6JxS6Pw6XUtv0fEGKZ1KskeLyzvmUHtf+0u2CPv50Hrg6H3KXov0V8rkvDh6m1UQUAISU3QvY4
sk+ykmxdhCOgnoPEFA/Aq2nMHGf53r38Kvya3sQDdbQrHHx/OMZiDJYT42xaZkQkCYrhsYZxh7K4
ecKNQQOeIxoIVILu9usnWeCzAB73I2xlZw6GPqRDcvxsMI9eMKRxgltCY6JIV3j2rbp4jhYUYXVZ
TlY7TCk/MvrHMWreZNqaZQKWWm+1CXqar+Ajr8LIeHBcDe6qMg9ox4zKGPm4L3Ea+/RNMHFSlJU2
fQpUeW32n2S1byFMSfsrmIeGHgxcXmpCknTIDLj7xAxM1OuKvgygSdqRSzY2xBfOGrVTaK/PhlS6
72UXKnYoNeL4gUGbTR2GNIx1g7xZB6q15c5+09VN/Ec0nqfXtYZU1CN0IBhlg0aLOs13NwLe096K
m+HcI/A246/zGjkcuvJRlp8Hb+17LJ9pm6pvZjTcB5x9Y6IaEc7iwnJbpsZ32RSw9efWGT4G/vhC
80iYgp1Du8rP3BaHzo02E/A9y0jK4CBRmR9837dTB+WXDkDnuSLHF7IfDdIhlTuCjfd/cA8Mv/Zr
GBF5y4v4o/8DTJCDWxLKVUReL830ZiQNskNr+I261wvo4qLaxqePuNBF8WTKv8GWq7m9owU1JQaa
mIg8mVwsU+HWNtqcRjWk6IHxkoJ1vZO6QMRqMmT9FrQ6PpzjVRrq/y9o0P2C/7kO2HmOzf53wQe8
eh0SYLNEls3BaDWi1xuHUenvRtPFeGexqlGuo05TaFtEhb/ROW8X6vM0NQLqRWaY7PVuKWi0tjYO
ukjiHFqMN6DmSxn7u1X784l6zSYiwLOX2YhLple4ZOkFi2/40p5zulsU36WRpgXgkoVMUBjIzexA
q/3hAVypEtYaHm3U2EKzBz2OzQuknYq2mdnfvR2/ix/a27y/DbKzfxCEA05A67j1vuIpcJ44ft2P
ko11PStTuuhvxQgpx3q0i0nkKYc+w3Vb+J/MkCjJdTaqjyUz3y3vL5Vz3jIyLrVgQVhH8fPXD2Qn
wgCXDMRJ9NsT5mVy/2RLaS5Nn+HIIXqeIL9s0RpSGlTDBbBKyB5fWutpBav2QM6MIRVDSfSp/PLL
LTG6l4QCCrfO/PJKs0STFvT7vCF/wCK7+SNr/KHcjGaVNj1JrMl7cwArGYiH9L2ZYt8IE9nNFbUp
wPHPErAp0jBcjsjJaXNRMgo+oOpL1jxvpXbXalt8varBXf5sxcwxXk1Rl5Q6vyIZiRQhc3snbW0H
35graNBYrPqsbToiMAy6Cu/DP2DF/kPyZTK9ttPAMQvrqSsZOVXK2naLr6ejSqnuVSHdrg2B7eJt
ElnMEr1jqj2Jtbp4KbIv+pcjrSt7qx8uRCFJUpwQL+VymigCz2gfm0okxXP4lxeAEWdEP+7BVkPd
S60Sb9lqit16FNg3BVImkA8MJsQPeAqtqRNFREVhOB8Nq/eS7mpSH6yWJzeRKhXnFn/WeWVulLUK
e4uSHLfmDkF4fWLMHbSE9MdVwU2OkIypjPJC/xCRSegoO8RjFw04LdmobMLU+do//FhI5HfgpzMh
hhGuarQmgkY5ecqK+swG7CAn8Tc0SDdBal5/p1Mxy6T4TLJfss99Mxijk+oNkBp+nZ5kumbKiA0e
c4YsAwzuSAE9vqAmNy/iZIUmW7LNEwYpxYpNczvnjuU2IRbloXhXWn5U/m5qFE+7WQWfBK2myRyB
7Y9WN2A6Sa0h9yCTqLnaOeoesCCtUAo9G4LHs8Ph5neUgvvxCGIUqPBADvLSV5eTp7qezg6NLvua
pCPaKgORTXRcLYyiAXT63bQfN0yt74Cvh9JhnRUnXnfOR4UlyYAerGQVNv+9i10HiRqYjswQMtqU
v83eqyRQm4o+feDHxo4fC6OsS/lkLow1YGN3n5C4CB3dHTMAzXZnfBgBCzE0N949oX2LtWhFjdwZ
jRUmqei5qRp3tfhwbr5yI97zXbw+1TcVzi5oThWBJbdVJK7NJR0o/l9GJLsYrB1F+c5cx4vpg+vm
xBjIJmYc1+WyGApNzr1hx65D4CozUY1H7PboIISXPAEpiTydmdie2OfwXosHThuo5cJo3nkhgAg2
Qt1j8qSTjw5P4drps4TBV+nN0Q36iojG6eLpQojGwpYG2YybOgXDQdsf7z41UJKhMTdxoOPkDxOu
YB+OuGuYo0BU16IJrse03LXP626JOe/RKc1MEg+3LXZqtKOla4o+wlBlZ/pyGETQCGhc6FXDYM9t
JKALxEeHLpTVyK6i076BvUx1/jEW+h4QxHUcT4Ny4dPgo0NJEGmHM7ujRgLi+hsHsIcdy55rqwTu
FC+VEVb4BNY+WRxkDK/rF+O6U4oVtfbtdQzsGnn3zX/RET56+k3qoEHX/i9koypOcrMvNlRUiUj9
bsV7+SndEAfrsim5VaVY1nOQnvxnzkcnlGj30mt9rv4z45tjagbasxaaXmaNyDqxgrz0MgmsRPta
ggWXG0M/WZZi9zSUWFRyakdDWeK9wok4mgiVozeDEkXbKrBjQQar8Su3SwoaTwj73eM9N+A7AP4L
p+akMohgIOFKIq/y4MlImlEWYloXO36Zxt8j7TY9cY1mFJsgvHxJpczCPyO4JREZNs5Nd23PT8kL
TKxx8nChAm1ZbxxCtaLfUBS72AY2U4hJ+RFqE13kyOIJ7kjlMyIfMETuDjdjme+/CEVE3kj4aHKs
bENo42Q/uHhA/uo5xMo8m3JfyNgINI/Yp8tZQhjNe57Xe2bYV27bZ2lrjMRMzB0LGGLJEnMaPy/s
AgodazHnxzRU+Q9n1PLnv96hPm2wxcQH0ZaktC1aoN7UeaDPFah/cnCgzrWnvb+ZwrLXT57VConU
yzuuwYQ+CdiKZN0+C8TF/ilFa5SWS55OPz7btubDSdJ9tvKkAqqOnR6OnVXYqtYHVGM/ELb7QrXs
u0KDWxvd+US69fz8fa4wJ384QmFJbfZ7JJInyLP/BDObiXsAXp4E93k/MRHlqilhQFrlDnRxrRXk
/CN299sViqGrnRhS+zeHgGz9WnXiqlZ6p5iuceNbaH7diiyUsdydWyQg/s/maLxnWAd+7yqw0u/P
8Ob6f2RQ9lJnftk7g3q8goh7YOJ9s4SvS3Wtr9CP2ol6JaXETbyIDItQdDaj4EuQpAJC5N7lGXZM
rw4RCIKe7WpTNAc/QN3ryKYWVWZCYbQp8fXT3hmX/AYJ9d+PGENXPBVALkwtCMvtUeDaJjXJ1pnX
Aulu34ttdQM1CZ4mzYNiSQ0S5BdB9FEu5a17vRdrSkMiB3EX5JtJOXOu3rRXEY96yj9D5eU+eWfT
Z3e0wvSu8h4C/M5toDPP5EkBGJCbo9L7WIHLJbgiKh8q+F2PzAqqTpL6/Xh/VkkUZUSWZb1qUKuw
Z17U5FsTpNn2BCntSF0u4tSpL0NpOz1mDtYPffGyxjFpvyxzR9YuOz3CWUviQHC26rm+OqClshYR
CzQB0G7UarH4jQFe0iMYQKrR77oZMDPFdgepnfVW6BAYgLR2tbD5/hB3zKR6DDCWS3gaMHex6Yf0
UcULP2V1K5VAfrZIBPjxtAMWRff21Z/vT8q8lX7cIP3wqSzg14mlIlWQlTcBiuLLzXYiymf8mrw4
kfVnyBZc/DMsQ4rMA3rlMi1supJCmfGEasoISJ5pzMOKv3U0y58Mfe9EDfWkSM2eDJL7uFlIBnLP
j5B5szczSkCiypaMdLz0KFE+O/Q7KU0OolUH4RmzGT2r1S1p84z49pBWg7a93JP8+RGvhrWpnuHC
zAk0qkI39oCj9i8NjMpOwA/hAeYR7B0keRmvIqbQBf75+xGGD7ERfr/mXfwDGWAeVlJi2tLSP6IY
93JYrshBxFeCcIkb+hIxHHDaSPlx2z+WRwJ5JvT2G4GlCGVun+pRl9FCUpzVkoGO7gFjfGcCzbux
jFsuNq4jFc+AGwwfiA4zz0Xz9gj5KTK4A1uvNGw3GVJk21Ovu35OOkeemtkfxorwTMFHtDQk4MP5
pHoFE/15RBofkMROgRpM9BgfJKoEPgxRtuL/JV+2cdgE/NBki3ZOmiICQ85JTSndK3Pe/mNK36Yu
wEDR0XNEcxf1mUdeBpaBU+Q9Tr+YrsTwCotoW98QFhGAd+T1lEwya52EZ6BKdCKemBCTRGmcN4Ct
hnPLG0yJPL8M2LJrO/jQ7BmiG76l9//cH3GxMqUo/dIuL1PC7gploFhhtdmr2FCxQ8hrJ72lPAFf
V1BSAgq53Q6znMM2xqJ8J2bbYaLu8N2U0tACo2PkZgtWhj7oOmdck43Nh01UsQhqEFAGsvFfkMBk
A4ByR+IbcXSLXpM5Sd/SV1EgA0LV+0RAM1FS6UZ1bYiFX0n5ihzsjeTusgzOpQLd46V3PhBSfvMF
5FKckr9ZgiAltJvMKAnrSbV+UpdQh7NJn+xl+ZfFgLmQYqgZBPOxHjTi7/fBZoPQf2Sz29zyE59U
jNYFcPxsAcgHFrEPjWdPWLaIWdQwMWLxjEZt32SKONNszESXqqM+FZLOxX4xq0NFZpeE8faav9e4
lQ/Q3M/nZWuntXMeR2363cxEHcNv8fZoMJ5uSdrXwssf/Rv6cjmmtrAOUMXK4cerc0cbO/OilJax
i970M7RCV9stnahxg5+WWAERhS24+nzRnfvmJgJKveKVt204hbU0DjQyztSx71WNZZflxZ7WA/Fp
pMYTI3gQLStcqCLLGRDLJdgMRL5AWIxqFNdX6uJKF7+rcP4mgKrkvzVL2kraKIaPQX8ImD+CxWOt
Ou33cqHgWZqosHJ3qOdd4e9Kr8Ffv1gHJ/33BCD+G8J02rlYtjbrcdpkJKJ+KymkmrjytkH6dR7u
vRMCTDUV2uQkJVp2CFbUAmuPV3cJ5sgPD8bslEPAd0kl4AIr1bid6z677W4SeBLwbQ+5/ua5J/FT
Gsbx8Whz5aEr1k8lz0PkONMcB6MSFw43ng58t7RuAw//nZ+jei82PKrvDBvx6adHMRs5xBaL/R3h
r7JLU7JSJnRpEImq//l55wxzlATMdOOrkT5h59Sp/ohSycv8zm9lIo1OMdJLBlbjqBBrKPPpwBgt
qAvkd/dKHb620itF+7OUmoW4+mRIPJsj2xpuI97ZFvQgv1+fH0AwQECezGkOkf7blT20MRkttTqa
GPMtMUgw7Pf9GHbfyrXiNbnUZKJQsBigI6X229E/T+fw4P0o0MoW/haXU8yZOQO3CKspHY7V2Ogd
ezIKw2k+TOr0dlxUOOhNqaqoSWYSn0xOejTOu/PR2Q/oxn5ILFsAH+PWKMGGJ+WK7bJULgvxbgXl
k+CRDYPqVFO/gck5P71HSYoxtcMToy1AmgKq4ZgyGWpSgTw/wSFC3n5WtJHNCfNyzT1vhP5ocD6T
7xRgerUlXTjx86JjPtXmFOLncrQh9Fxjoog+U4HjIcLDN4wAWPOZLtx7OGRw/+GAN0EwJT8cQRiB
3LViRSJi69OuYcnpr+mLGKNFDjsyFEFiDf9FTg55K4m4zF4N5lpGZqi6HtErRYhfAIQ3KTaqXMro
oED1s0bCE/QEEsS5tacxkScYOqlpTseyPMRUCEH3+YMImTkNdPKSrt4aUr5olfIL9vioH07b8GG6
gmcK+Sngue308j5fi3FBsueVi7n6LIQY05WVixphFK5YHn3chHQPYR6r59CGFZTQCajdj4xuOoMc
sgC70eVDwoqPkBX3lnxJ0uGJZ619Br5qejt+LAp5fPFELUVfd+OBaWa6upB1PhTHQ6Q3EM3QyCtD
kz9iHCkHn+vaMGHaUXBohoE2G45mtfbJ4MTi+Ov6DDkxQaalbKIkkK2XCPWY1TL0Fb/shf7xdTAm
z+Fbfw2YeKBvM1O7Jt2sAZ7+bMEKSbREi3BX7DeL2RTKdC0bhBWyoUWBfVRSR/O9UsbdcvYAwjjv
udhYPIuQR0actNLk8Kjb4+p5LdNoAJ2m70n/mXTWE4IUT8caYitzupQk0T6kXDx1VTRHgoKcIqya
agWMqWXGFDdAJ+tG1gWfDeNuCmgsxG6QaZHcoKmsx/R4F64jROg/WIVjc5ych+xhuoMixz8iRfQO
Q6+Hg0L8iScikiYRchWCz9nhfXUKEkFjfkeZDyP6dSsPDuw45BZUuXt+hXl79TiZVOlVZ3GXXuhj
L8W0zpDL9KWXYQOjmiy2QAAfGy2SEpyXZPLbvvDQYNTBN7cl4K7W2uRPfn6nYHTaXG5Utuvus//i
QK9LRVNQgnvo/MEGacSBFetGXHeUccoNZXBHTd69geTFUBuIA/IJbXIoF9sid/RSyP/xWPkLPgi3
AcBWJmfLfotZS5W0z7dEcumwzuP9wMDek+zZkbNay5xzdggi6hcQgejir7cbVUOmnuzyCofAmymV
N9cGOVbGaai2Ivk0MBfqxfVJVos4Z3/+2C4WPUS4jMud5QHJM580x1a1tfvuZ0j5wxM3CyeJl+/M
1rRHWvkjFCt5WF+l+AMejt71/3b6SAxx1De9sC+hejZS7bJMKLVcuirtgOwVNBu8Ow1eUAyX3LIZ
ndKzDg6NgeWImI1k87E0XIZqpB5r/tQ8igPcVQOona3b7otKMb5u8w/TPSxnjMoA1NU0XIFOhACf
fKGuK650H0Vk+kfD2XIO9hwABNI/SbICW2J2MXpOhKx9pwy527iQ7g1fA6x2Ita+iivi7Auq4730
VksGdqfgZGxKTdRa4yruOwHBBq7DUJl52n/aonLEhEt71lCy/j36e4ovsQunzckHSWj2EP9SSHiu
HmUUaENaKSiPxsM2XPV9adH/U7eUQY6GQoyRhPAyPe4OOQG5FIeQ1kpIhW9C9/4s18+xg7HHGrbT
r+K3DoIvqD12S3gI/pRREeDzCgzBLC7UxKubYnfCPL/hFxzxnlUxxRYm9UqNyMCxLXXoMjzN8OWn
xc1gooacIB5hHNyofYHlWE6yc0T0QDMJG2O7WPyYhxl85PsuYCyQDhjXI1Ds0Tv1PfNYe+igr7hE
G/iR1c5b8z46EiZkN/RGWcV5QVBR9N0MC1T03lT5w3Kny3+AgGQM3mHp52RZOK+rqzXPn9ZiHVkU
J3Z96+1hJZkDPDnv+8zNOc9zq5VQlz1s5LEI9P9Cvs032HIeQ9911VQVEieqzwkGiQP4U/yuvY0e
6Lpm93R6e1QjfX2dEXdWccsRLg+4jm7C4KENmfMJQmFUHdOoPy7/NdhRm0304EqioPPWerx/XX1N
HV0KTPP4ONJM4EYLcIF3arCVA5fsKJXs1lhigslM0/lhYEwwSW+xIVRVTDydQfUNVMlM+YqxYeUr
BtW3y29H/wy6VY10jWO4s6JD1ByJuuaI8+RZBf/mbZeCEQNlK/ux0v6xuUuJeBw1eahnj5y4VZ9J
uU7JTwH3EaPLSZnrNBMRkeqIueLMU2pXZBD416+9l9d1RoP9dkK+yY7q16e3pHILkYQCOlUMJrqV
/kEb03kS5Lhw6rMTG3QPUtm+vx44XAlXBSvwUPVDdKZZvENse4E0UbMRTG8ZF450aVS/u2+EFEtU
wf23zoWHnumM4cTBwZooywq+UbJ3AFV8A7d5ZGW13Bxcq98qyXG9E39Bw9y00zUr2B91ZIHcoq/f
w+CoTviBqwRITDZjKVPQoBD75S1WnuHUCVt1DG91M4CGJQcDoCRrmI1ubczjBTdH0wS1/sePkGv5
H3t2HeXL/BhmsFrEkfFTch70o3qPXy3KNMFwTlg9AWgRAfASR2ZnGPQUz8uDBMh9HVrTdG41Z/JD
zRM70DGUjEUCgUKPHqbjuptFcFvAh95c0HvPeXpc9Nh3/n5qKC4Piu4I4UKKEedfBSeCvKCfAkMR
KNg/iZ6bJ4JPVcQRZRIifX5QApmG7T5MpZWAcs7VSUemVXbEfSIoAIweJ5ayDhlOOjnNInfiHJUl
+mVS4Ut3/wkR4aCfWbYgB04Fiouswy7916P4tuz0J4acHtWuGhUmcaxHqHS4qAZHaPmNrGfbvZSq
5se8/zVRyPHMOKSmYO7UrVmsaEMEc55KsykkG0S9twwsIVF79G80G723M18bXPpIyhxNrNySoHDb
VRiV40xvS3mtSNagsaNsycUMx9ECO2RUoRWody27Ck3oqh++t6zSite71M4vouhHedEBI8tosWgu
YNKdwZRvFOowMmfZixvY219OLL5/IVXCqgPoYQJMvspljDZ9kvolA0dprhcs5upNF9L5FV52+0Q+
oHk9lA2s6WrulJW+HPifCVoGwyxmVwD3W1X4XYh+9xg4FZs10walZ+csyRC8oIfFZUXRaw3OX/Wz
QYTnQJTjMh20zhVTTxhmwAgE5+WW3yE7ijkvHGpbl05hCaVjY38hQcqQZU1xgkjIz807HRK1GwgY
/H9TjkbdoxLAWpBWLAFEaWBsJ4/sAIQUoEYgf/xc9m1nytRxqdHOU9nbmmdbKlF+uFJCLXXIqNRw
Fk5vBKKRBU40myBA2/9s3pbJOikVwHSallTnzq8X6poza9Cd5uIxtpePbXSUh2fMVW1mr/GwSEy2
RkbQjN4REJOOWfm0ox+kNforaqowZkukJs4qSCXdyu4TmSbOYI3oCLUOFREFyNZy/qxBxp1iaguO
BqFrbq9pUClf7ynjdrjMMJRRGymoMEJN+vcXal2lQUbHKU0h0dbc924zkYVEr9QoageutqdwZSjg
/+HXvyTxGHXGpcb3m4/7f7qYihc3SXXi9B0kjwtDKBKjzGBBAYOKJ9ImaXG8HwApfzT7RSg1Ebd3
ZY5lzKXAs6l69VsCesR3dH9YQFwjcrcQopUG/IEE9J8OCuTT3yinQpSOFY8Do17UCLzAQjbQL6zA
n9tbhNNEHLHbRPnGl/8n1jsDjgr9KH9/TW9Zv79ZFsNV2xmjS+QyTmmo+mBi5JcNSynzCg9bqFZc
SidayesChP5H6zr1iUXMu5sHZmOY7eCYUXNyyEbKgyX5+zpcZHuZtO/yjviKyPkq16PR1raDowHZ
a+5Xo3LjWA2qu5ibw7Ym715FqfkcaGagjdWYSt3/o9T0K2DD7v3caoYdE1SmMPTME8y2lJBeK7Nz
GIjM8vyY0kiYbf7jvDkUYXkKC+8+rglkK6fJfsu/5ATOI5U8I4Myivk10Q9nytwCl6DD84fPfWin
7JlxNID1SAxzGEqP1+nK69KTbJkJ3LbHHR5x9aHJ0bjxlKc0BkTdF67eIs+JgETM3r5bBis5/BwQ
3SaWyBk8nE33BslvxbMHM+KizU3wgoG5ixkVcFBdISlA2Q0oVn1D08a4JqorqB8ROuixHomjO8DM
otjigTewvRkb3rW5qdx3tlfNQ2KfOy7gOOOY8Blr0p5HOwXSMwSdJBBHnX5jC1s5qAk/NG+PhHUc
j/kTju32RHzQs8KTKMGv3Q9P2c5J0J0yWfRp7W++4wfPrMKqbVbxL3insj8T5ApDTIfOKrDrXuKM
ymHSBuGF2xuKOg49kVzJTBSrxwDZplfZ7X1jpZ48zPHUSmWTpdVV0v28+SWwRAeXUjzTkcZiJHjB
nXfATadZFwGqsUzKXXBB80vwzFTbzWDdysyJE4EYM/85/fSGlcM/i1X190AGoxxRM9Q/acADolAO
+8MyXQRHPLGFEFy43U7P+n6/mu5++5vC6TtYvzrF/ITNVnvkS338ByOVFjHg8xsMwxc9S8fiL8KJ
a5+NAbNtPFj4muyeQ+p8+G29VFL2w+E9MIJp5FqcSUJX3f2kuy1s7z8f4R2ki+i7yOH4HHRaRqZy
C+OsdyDo0L6AcQ5mp9UZavMd48yEi1ZnPOvhuoLUzC8sAujh6X7PHxxkbrczY/hSeRS8zna/1DEs
5LJ54Giaat96hesViDM+NtlpvBWXqJwHXjv/42nUJMZabnRtJg4b0Gzj/N0a/DGj41jADdxaIX9A
AIlW+chNAQGJhlksx7WNpewVVgapMAkBi8KjsZuQtB0c9Z2ONXaBSXpvSDt2oPxN/bxAVumFlJ0k
180zjodUY3nIH/AuRQWChXL8ol4hm26N+7CnL1ZyypmtSEsWsuzhYk1vgzDe0bBKtcEeAeZVBtHX
cYl3TPjwo6Yv6yiB2jJr8M6fM9sRcjdioP/OeYKl/IcAZY+xwj1uOg4C4Ts/7UyApLGBAjZAk4SH
LSM1p3Ru6LoOi1IPjZlxK6jkEeL2g0dn8kAg3m/GfRloRkXa2h1R+M1skTbAYkY2geRQPLMefjwj
JxBz7RK6IU3LVpguNm017icnpSTE2Ix6ab8OcjFXLDae8oJrf8hkCgbwtwcWVT1xiZVxHNj0fpOg
ZVKOr9Y2rcmwh3or0yHoVbQ/T5WcLI9mddNNVc8/S0H6up8a/sx4XvC1mOXPOxF+Bg1R3OHRY4Bx
yjJrq5k/ro6NzAOTuiqGOcxGYnjrp4kTx51ft4W2G+J1bP0nLp7sUyEiKpda1eFhsbZuRdOCYoXo
TVgVCkYo7jc4fModgvYj3jzBtONF5DvyICgjFwrCAVhXOIIq0dqvgUPiUhMnGWeZQVHmnwWNUU6T
c0RxEHM1C2laN0NEYM9GRKDtQqv9+fZaweJUfS1y695N4T3131L8oSL/kROjQSrHpFGXsjXkZQ5a
IYh13leWGnlyvRc0nxQ3Btp0FPDsLRLjMWiWfOr6HgCxh9xcLfn+A4GPwckd6OaNF68Y6XEAAFbi
POAKvHKMegvbQcKzhha94ITIldjBfGBLyaAz4dY9D7Roy7eUnTfShHkCZWUauBfQVWILQ8P+06SJ
F7Uw22l43flhl/jGUCHlHYy6kSA+PO31W0v4cc/NJs5PNygCNqsKv0WEMq/GyZpzK6gEevoRPm+Q
qzzJ3tYSpb9895owxugGRIhfgJ3JKYw9nCAx6LW/WdzO9eRfa6wA9Etq6CeIRjJ9AvGAsYd6Y0sC
CGWHnN9nZX49UijaeR4NE1ap89wdprmvvcVZQslIymf204uTD3vWAIqtM06DMeqEEZdnWa//9isZ
4zwVOHLrKpuHou7pSUohMIYPfEN9eDJjfAcsH+/wvF+6y8ci8GScooWiqywPoPU4+ATwHC+z9UsF
lS37FMhr13DsNiLyPb6pLlDmULSj7P7CfaVPN/glwegSbCMnG8BoHhO34swZSinR/sbZfTugtm4s
TEtwxSwlMXaEgG/BvagXcZWIHb/ErnJGViKlebIMxoywD8rsppgWmVPXxRQbX9YWMJB4Pk9RJdSu
eHcL7p9L534ONkCw0nGMybR9dYa/TmKxEujMdIY8ikAC9YVntkr0Ec8D/HVRasOmN3xOFFUuE8pX
H9QMsRzlpXV4B6oKd2RdKKtYWWkPSB+A85JtnSpNEWIoWVI/sY8ynJeMmfnJJWe2hvwergg/ZSrB
xuNVouzDF74ixZgSoXTEoR9AOXQXiUO4Pr1soXLiZob150CWcRrkMRxc6Lbj4Q0G7uFWS4U1JUcT
x6P1AXOBV0EYD71c2LSpAF00uZlV7f4Nd6uh3Injn7gR7nlAw/CIaRSEPdiL3deHpstTJHBlRe/4
CzXLwVmSRZ6nJjetLHt3lKjeBDdGEzX7niOxL1ejJgiCYiJQ/vfQSZ8zcz1w5yYQihZdLYmknXCz
uEfM1NFINsyiJm/6KbJ9qk3Jlwq0Ztt2DPztE2/aU4SfmRJBxGuC+uvlWsxf8OKBShdxsICEyJQr
M7bxJ1AKyvaQ8K8SNb0OawO9M8gGryYFKOkAGQGDAczA4jsc/7GwkrofFJyq5tG3XeNGiKIYl1rd
qHvwD9I8l23YWDz2uSvJAkTVKv0GV5VHJMs1pkd2ESk4H57SPGmNJXiUpdxphF6QFh5JrD9eaJRR
U/LOuHguOYZqV3TdbIOtv5i5Ic5+5UKmKQ+NF1pAs2LMkxizixNX9lcvSd6V2Lk7vEZeqAjD3Xx+
6doA4UYqsqj5DrR2YAvKW1ok7iaZREku51HBhntXRXeBpGiBTZObG4gTc6UtjOYxHQPZkyFqF/VI
eeIcEb8yj1goiPNLR2uUhyGMwMJO/lvaWjIZYsXvIeIhjT0gXza9fXJ+9BPneTIYtq4GvY9E7SIo
kxhnMpTAyuG+fyOfKQsJ03LI6cEP/IgBAjyEEnSaZRLN2BpEtoKW1XRhyV7AnWfgJfxTOa8lEv90
0OskbQCLgkIR7EljWRZYFD/8Hyqlj/tpUaMVOGfeMXbcWVcsrnVzyMyBi3iPGnocRCwWB9DZuR4l
vguEnHy4aiZ2l/GnejDjkuhqQaNYc3Sn6ARgde9EchSO0D9ScZI8BD3sy4uZNJAH9s2joiZonvib
kZOFqOioJhiwrxdNzY8g3zrGkJyhCY/xIicJFSdpZSVr2Gsp17btJJCeayxVJj+VjjgMYT8bvNzS
yQQRmp0M94aduTQf7aYDv9wCx76k26I9Vwm1EnDE4E8WpFuBx6SkNMKS+pvErjCOrhOYuVMXUIjg
NuKHbW2/R+vFlQyEGf1ywiKjg4eCl2IE/STWi+yvCMn5gTIgKp57F9GAzrsfz2wLMeMqUvA8VjIg
upcCNaaMPx6pvvfuMv93+k0dysTbWtj+DfM9aeLz6sIptmkm8v5kPdBAeMyZxColgC5afyx7qXsL
1cUCn249L1MbX6mGVIbhodWv5RruKeDsN5xqHtwxPJ/B+upmCrcTAYdieFxv8zEuz0/e+c4An3St
Sk2MHi7JvTzOxlMQBzggHFUSHeReigfQoChOWZdhDSQaO63hZflxDky4iU64M6rOhD0YbNaj6idL
UNq4mmmMJDr3vTmaH++OA2CNUJxnEj0Kxzv24iadZm1CPK2D2p3fyz3AD1/5FjerFIZJXiYeh/2O
zXfGPdm71FVnv15X7QTkqa+2jvvgM75eHsOdpy51p72mTA7nWZPu2u412vefQEr/hFASHQEUA71s
xqTpEhu0ePmVU/Fp1Y7qSxxFE8FR7VwD1W0Pl3PhBKhxV/kYBqkSgglL/ugWtY1Wjh/C9eSCm48G
5QuP6LLpTKp/Z4YST6zGeuxoG/H//YSbZX1Ny85EvG7cXppBDB94bnZ7UAvOQeldtTZy/cPbtnhF
2bDhm8N/l/TmgqlKg4/A+6Crphe6alwD+XibVqA+kCaWYHqO+aarw5Hsdwe0eMFBnvKQrDGtBXCv
rof9VHCB0nkAUQNaTPOzo5d41flVCLq0YXBGJ+NQPeq5JFhn2LdrzLydz7I4L3d2p67zvhEixwCV
b1czPW7mzGQYUVmCNZPMFPHIdyk64nV1V/yuqHAjdeeTsaTihIZI1fnTYSoVHQ2XRJ9emBsSvZPn
9/FusRdNHULZTOuugnWNZwajh+txlzTXsyd8sRqZguvTitUnfDGqEs/XvdCAGKt0aoSjuGLc7ZTP
+FQpi+SgZ1tw+x0a5XnSG4AU7Alspc9a3GyX1bOCVAkAtuDWMMliHUQMmEgipO8LyZPF7ZTBGOP1
bwNbJhFcu/YhkUdjsrTNteC30L42UeJU5e2a7BBksibXrBWZAXwt5zHNYhNxXwDeNhtkc8ouqJFT
zXvPBZl0BcWlH+YQ506lbxyeIJ8YfKkeeZi2qaFBFjo7wX7r2dzcL107+3LzSHoLPelY0XwNKlTv
uYXQJakvYLa6Y3KpqOXtv0EyBRq0Ap25UpRK8yF9LyCguXvimtM1DyXm29ahKtMwsnw9lMVsBUDQ
RS7PSjKYx8NjKc415SfAzuu5jzaysyNo1/zWmiGN4CW6MYXuqwv00a32F6FhgmftCWafYFnlIlWq
fAacmyddQKaiaOlju4JsGlnQKjiYZslYKKsfYkqzpqPymi5CE9x8NYU4MIUe7kFnahV3ayMgLtmm
H+5zzMaQ/+a58RJF/nrQioI2oFagScTCMH/JPl7f+ScOx0bYmQOn8mX1AGwzT0pBcGbdUWYS7H5g
ZLQEz6JqQNKU0H1dz+hLlypZytDuQ93Dvz3O3cWrZxF2zb9QD8PdvGIwPowUGtZvPpP/TlscgXz4
jJub13yP2L1i1JvbzY9wG+1GBzoRhtMZ0P1vpxmB7jkT3fAXzPIqCjAyI+qmHa4i2G4vDSwYZBYu
E+gEMPlNUqtaKH5yNigJzqe3YbFdBm73AX+GMgTldWv15Y0u8dE9W0UsYzQiO1yBiYXcYTEYHIGp
Cmt3i1ZznAugXSPIcVryMsVUXu2c1Bh6+bBRuK4X1H6DlyZEbK5PGsVqHDB3ipUenk/1+FP75BVa
rOTsxjEV1UMqtvzGG3x5Po598W5tYam5ZVrehvu4GtlV2aj7LVtFErAxIv5RSvpYshmIueh8SUJP
T/9ST4gSjdjpILn3uUvt9KJmFtuQysyoGvtAAaOfTqO4f2O2m3C0aJLqJR53I/Sfpnf1rgQza1mS
M8lb1V/UZ1aQnNrjuwxyGJ2jnSzHgesj0frc1GB4veus8rn4x0KsVOQZroIyWldub3VT+gpknUvg
C8I9+mQo3EwUnGZhGd543L+MWXfS7fHrJ/iTA5OXx9pP9r+CM2+W4BglWEHp7tflEW9vNf4dOCnj
Wsb6hV7pCf3LEhPq6EL7oXw+0dy1URfU5RTP2Qi9x7XErrSqqdt52oiL0EoWHVMqD6frTjhV+VA8
gHdUcBLf4gfiCVkeWLfTha3JQ9d6JX8w2KEqtyhF0utDsR5rcj8dfjMNQH65iUHm58Hp95fONdcU
LoV6jhGZxbEYe1pMHsQq1x7747X6W60xRfLhJ9wMUGiRi/oZjcV28oDj6KKEb8BBW1Cj4L0LU8Ec
x3dWc6Cw06Tw6Hi70+Xg6L1cRA4Aw99BInDAYSFW/eOu+7Vt/CxqijA+AV6BBHobhUul2zFcDteR
Bhmzp5A9DCgmH1mg8vEqWf1oIoMKc2PqlcpVtrNPp91/fTeH+eVVjKZnuCCM6xZ8FUKLJjfXuhUz
UytmHERjfquE45rfsSw03SL5XG3zpkROpxNpPZ/1a9a6DUtf9yPgX963kh1AjMaMkfoENFLgQ0hJ
cOLwXdU+9ZzSlJ+0UxnLiq1Wg0U3FKNlPHJCfL/yHnXKe4K3eB8ugO30bIFEXfoPxwYtfddPLDlR
7VCcXzSOVZ/04M0AWm5mxuu6kydsDaRbazzo/qZrsy8Vu2s5MTCFNtouRsAZcyTC5ZLgrkv5UBU2
xhYKRVkezKjtIiSjYIf9sx6ij/UeJmiBcKMJFObHXSWixyZwQy+cG0P8ReMTleZ5bWh7oszFostJ
G2DxX6LuzljWT5hnRHXlh26G8YuB0rg4blsiTUJSz6r9gNEWNCnY1BgFXKL0OTFyde/FKGxs6lO+
xYFS8KvW70xvW4ce4fX7CYkX1SKtipi/0ypp9QzKz1pcvI4YPH3cRwXPgAifwmjdI14UKKRGpMWB
MRyQf85RUvIq8CvBiA2cbb+LFnxf9DeNxLBpMYVPtpU+WF+JSzi93JvytoSF+qR6lpaP9MZT6m9T
crq+OvJxBGsqSgaf7qUfPQsF/+/NLcKFaFK/zzN2UllMQCCkEP04TfXoSjn3bS67MQ99A5KCFnTN
bvROUrq4uhWgY2sJs6H16LOppEumujZ3tWp/eP+N4YyQ7k+2OAeaVpvWZs4FjXcCcYST5xRg/iWS
ojkAmAdFBMHMFLpS56U2vZoMy0joi3eYAr4u3S8/5bPncPVSmi7gaizAyQ04njcT+YaaVpGLq15B
sFppD8mJ+6m9qRy+rPeIaNtHUrx94mKtGOuVvxYk3cRPiYmGdGxsUFm6cEL+xA3gc9ZlcEUt3I0E
+aTvv6WKPgtRVA+vUKfV4dwg0I6XyLyGBaDj8F0bjlwSw3pnnlUoCUp4g1Lum0qBajgW9e9VjVQM
zg1j61y1b/Yxip/np2t7itZtkGKPtT268yu8GrQP+AInICtDPy5NS+RotbnlWx8o/HSu57DIySOX
lK3cP43nyRIljgrlODzLJu+NLZRl82O/lHDmJRADfVnVig7DSis7MX7NtwKdNhO6MoqhwZYEJOle
jOzcYVKTYGlR1CciFghPM3x4A9VRignIFcnCEKfbfyfk4WlrqbSkHDRmo96HOcLpgVlLPMAj+FTQ
SN27r1QMCQVpWgg/aHdwM6OZwP/wxefNnsQC6tluvqQn3McA4Ksegh0/5LS8YB9zlC8DKEH2V+Dh
4gK+0BBiYUZ4gNeluPlY8EEG4B0Z3YfZi3aV0VxdtCpZUzm1Azisq0QKRc8kl8VLI6EOX5mh59Pc
vq8h/7MwWyX0Yoym0c/CHlhbxSOntmhjnEwwx1nYNnSBFoXgSbvsdtnjNRliDieaIV4JQ3XVstge
yl++X2OHqbv2MBR3VNK11wErFfopRDfjnLkKzDZPxsHoTc0GjX5Pd66SxQQqLuHlVkdcwP+FIZDV
8U9din1vKfnodhCy2RC5Px4CwiE1inV6s5UBX9hUI3T+5KNtX/dBk79MYlJTT0JHzq01aUCia0/Y
Hh9bnYxQUJxRzM5l/ZVFZNv0m0TZUPtbQCB0kwRo0nA37yYS7RX/QQ2pkEIv6WbqLrnkhgsR7Trk
X9fbLGspY7h2AZrO6+tnanCTTnlNkvaV9a7twSF0G5W4GX7ruEQzi6yoZ8EPZjEwWhg8sOYlA9u7
+6jTL3FV2a7340uUkLn1SLgiB1gbSv5y/ufCLXXmA2BSywC8SDywjmrj31FRNgMwwHKDXnfo33DB
9lKIyRZBwgvfSYZ7umAL2lu0tLczDNwwR2iZGrxILUuyPoQHHZz/HCwJiGApXHCD9mD8hG53C5//
N/y6dDg8ulSpQitpKM471cYN37SiE8wX4UzzxOTweON3RtLNwd2i7mE8tzz1j7d7rwpCjmLVzZ/k
D2HSLctzSV/05J2WuiwlKCwsQPk97NBTaX8K5YmBCq7Vimn4mEPn0Qlv+nJ46SQiXQ4tBGvQsTqD
mnd568NY5CQucDzzVHnqyunSrVs4SdWqdPoEn9OjjRHCL22+CYC4vT961Y6Tv3Bd5T7HRp/Ueb5x
PlqlYCFSXTH1kAph8LNZdU5RS3JvynFb708bziwigwJZA/hC95HuyT9Cupgi4OAi8bi+L7W+nmf2
kiPHvCK9+dmF6iL4lvv+5JXjNFrE62+fhtNIZE1NJ7TWveIU8VEw1lI8EFguKFlAW73Nd8b4gKDD
QaXsVODp/UkHry7BAfi7ekx7iC/HwmAVw9LQWZruVmMR+/pUEbAupDhy3+HI1RdwiiBLtDwXpxof
u+8jp/EgoaL9bM2j6Ctz6ApmTA89cPkfM/earyyWeclexP04leug+WyXYh6x4AkZkhZX2VDGB2aX
owp7bItGW3ZRNNpoDnZ7FfCFWmXzYFgUyL2/nCNUCJjPbDmi6N8rYf5QFAElof7F2YF2WGRmPksT
RlZ7Rlh0Uf7X/HYFzk9HEf76Jc/uIalI5VRnRrZiRFeMBPGXIS5cltC/yj42hP8aameeHIvT60mU
LsFIuQHYWv0jYxeushdwU+WuRq+H5iHGh54ZnL19byd8RsA3TXpFJVRWRZh5CM33tlPliyxnTG3F
BMQY4gV1A//lnCBCanPyXw4bjEAVhLWK8LL5rJ4ahKTSWT/90abOIvn2QJOOjBJHgUUPF9cNBxvD
alzcKD4cR7iykMtX+yIemmzvj/E3Ta10BzxV35XZVT9l/BS4TMGZez91gSobYoHHTQGfIQ/iQGzz
5LIAjqHKqeREYg8RJU2RokZxHjEMVhSXVKLOoadEBJTwYPE2l9heGhUZDjb7wJ8SFtThRo9WBYrY
3ORupckXg6iOlOXY9F5YXEhlynkqN/skKQevgafp9zj6i0jZMJbJaZEZXpMN4IHPr0+eERFC2Bou
P1dYcSi/1ZqOSE/5Ejt8wLywzLcxkFOfxIy0PUpVFQHpuL5aFOA0OOpUeRzVCGKMGh1BAYg5GM1E
h4nXuYgFGB/+xE4pv2mtbLct/4kNvtfU9QfR2DfpIvj72aFbzPP9X4cGRCtDvAsdDWMOS5gC6YbT
Iu0Kcnfm1IkrJT/lVx+vnAGQ1LOcQ9tF1l9Amw+w1L+s9HGWEu6A+EUDcGir4X+EYgW4jAd3n6UZ
UIfOGTq/ZkFADrP1S0c9AEtZm2QHzmuXkwG+p1+Gj+tmvBmhRkhdYnqBQVWZxoLQ0M+iYJFXEvG4
9+UwJ1TnEcF8UNG6x/VeRRQsd+t5BJVqwHeHbgAqA4kHdiOZl6laxQuLw6wq9IWmTP+1JEVsTrzn
pP/YUtbUEinaxLTa9XHMKR33ZMb2EhIg6JC3/dnrX4QNXyM+wo0GCjDdDf9fG1pJmMQ8/ivkBaVy
3X1bTepHLxdt6xRyrOS22T1mOGQmnOVZSuIUeDOD2o/ZSrfB63400iwUA8kkReV3y3fgt277vFss
NbvxfZ5gBdmyc2SqVW1Pj/Vo0QdZ5IjmFL9xdVea3UVkGphYGT1szEcuLjZJQwHoL7iU21uo1QK6
DHQbYTzkOhDGQaRq2w1ac44QS3bCbmK88cZg+BNaGpsR4YjA2qfsz46gHpcjRj3CvdT6vSAjmT20
PcEN/eOuLUnCgYbCelwsYjPWFCIMkXrPTsW2bPnodghkTuPhwd/rvZGKg13EP8f8Nk5xfL32c4Yj
uTstz2j3dZC3Xi5zBV9+v4m3poBTWVfC++7BLMKaE9OVyMC2UpJh1vBr7o8VKPSU4Y+GLBARIu82
cMBJ92vOy7TfaSXQeA9OPpRhie61oSkLQHDvlTfRbNNL0ygg5obXa2MbVj2T+fYH6zqeHUjNJnSh
dNH9dgI+yLg0eebqjtHWYibHsJNTKCfu4gqutxoRP/NrDSo/rfjRsSa8+crnCyfe3QJ6nZ5b8JM0
wEh5CfE+51HJCDPjA+IjWqBSOmRrWfe59jo7gFcoaxUKuB8rQi6ukPhhViDgGyXy3dzvoG/7x5IL
dYb2M6y3X6bjDEDJXcyE/HGoZoNesIGqHeE31g0UATh9E+RtZDefjm9DiDSZbYCxBQKPrYly0GZQ
H9xwzcb/mZzxG1n9sFekixTqJuXThRWZ0MSH6tyyemIXw615vP5XUpWnv4Ug+TOLlHoS5QxiyJf+
cJp+ZMs/f+xN26M2ukQVktYVujeLcuZilRpxofipXs0MYnCqGu3UBbHas23Fp3WUXZkhJIzJYdQb
5MFQcUFUVjo03DzaoBxIq0SNz0PvtPIG/NUv/EHSgLqlEG9fcPPErBuLG7kpPYSxQX/PX6Dkr/p4
lGVadyf8Okwy2hHEmdbqLyfUDhU//SbMbiXBQZjqCQR6Pt2e80d7PiiBrMtO95UNn4oRLktmrW6C
gLQIiVs0e4iHym62BRVb/eg08sjrOdEVGYO9reg5uZTfn/60wpZC5Kkfvt8U0pc7bRJzaNNJojTL
iIkq85pGIbBm8DaljIpPfN7gjIh/qryNTmP0Fpu8rWgteQDl8J70boRC3DFYKbopqjBhPsmgiDf5
RFopYs+Uberl1nB78Ifbo6uhlgoLpKeaEjG5ziVL71I9KMK7vnap+Q5t4VWIn6fx1jytF4B4B39/
LubjrDqvbZEFB34r4bfmxjlVye7OSB0FnZi1UdWrefOtQQsZ0UhRMo1fqG97FV4jPUmHxqtl9dUO
3JZFuXVkgYiBmRI7ehX+1PzNq43kYuM4aEvionk0vMt8w0zkoinYq8cm4UVb0R9Hlb+Mh4FUfFih
hg2YxtZqIhTuWV7zgd5Oj8d4/OTZ2lqk9cHkL/nAPyRsaanCg7ahsXQt5eT4cAeC9J5zdXy+ftAd
H9Yi6dXvvmXfjAdE+7uls9MQgz0/eNl+kcfo4n+bWRjbyBXvh3FJZztvuuRbSShrewhlSfakmEaD
VKim4Vx9SjWvi0LkYNsKtjzx3aocTphotyMxzichDiPyqIGYm9bYsSKUVDGXJdyUe92Ru2b8Kkmb
iT1O9klbdFHTm/V5w8cnX8Zy63HjLqgVO1OBgsePSVirj3LCmlBcV482F1/TiZcJRWgsstrhvnPL
877WmKfllz1XJjG6jvMrE1V5in2dp8j8uypuqvpSbru93RgDOiLBvuNnLLOJbjfnXGWqi1JQkxjD
U49JXE0QUctQjVEK1uDwFQ4iP8LJLOVQT7E8IFAaoqTdVuzBE8g4CpR+RliUfXM+VGQ1kz7Dx76U
3ZKBVev/L0dwlyEhbsictNainYvwmAkJX4LEUAG+BTNJS3YFrSWAG65/tZqIm+z21HHt+ueBaJ0U
jMhFPuAbmp1M9VxgGSlyfMSX6X+bSo1GsuW2TmKcl8qptYsjqXGROQFX+0tDqsCId1IYrRfUUxIR
0+IVnYpB1GcxlxiEmnmsSBh/OyW843a/r/zQdSDH4z/geev2xA+iYYya/86hdLXoGKGfexEA/VfB
bNVCNAHHp+tzvJPQxU5nmPEto9+GJavgNhC1YMBo/cXZS9+jYQ+pG3NH1KwxH4Ld11ZwnHcIbkiu
GNM9/sZc32UwT8kGlqgwrqWFY32yA5kcRDGxT7vMP9q+fB7QFZj4dsKZ+siLB8Eetn3w8nR6O5pY
lDz/D7IyBcSxH2R9lIhKwl4rP38I+ADrI/yVgAKOSVCZxAxMAjnNBe3z0wmP/1529vJ4BiI/nXZf
FBHa8/RZBUygzrn1xwbBUhwzPdySv0C8LbhqQomTLDPg3CnFaHM3A7m5rMHLwH+qwIUELb4YtCx+
ulXuGMXDUiDGDrs2n+Tors29mq7WcUF3Gcz231qRCOIwC8xporkx5hghsMFWm78Mzm8MP4uU4cLv
VYlzZqU9moix35ovzH+Kfbh0TzqR4Joyb3MAUQ0e2UReA3fWH6W70t+RmMcm0UTJ9gj/7QrRH8/o
z71VgkunDsD3fQUl0KjS3NENV3HCbo5oLUBo5QnKY9Mvb5k+qKESaw/tI6dpClv9D3G3fkk3q/F9
CSUvjyRdN1Y1mWKpZzlMkMyKGAnYWxhDy3XT/c87aACEoZbl8ggZG6iMMK9RPa6bwl9CKAD6ZFp5
6JYkNNB9JHGIZKtBrEO52YcyvpteZxRU65dyYXON4krzj2YRSxqUlQprlXBEYAusSKwsj2XoVitd
UlmmduEKRp9EW5qWDlKs2xx8mxYPKLbu9L+DJchBDqZj6MEksvNSyixGoiDpkdz5biRvrMMKzrHo
OG2RwGcXOtJ4ip7+FtsR1IKUI3pkyy6O7u3KhiGQnQ1eeEYM3k7qRVVWlrJ2PzpidjPA5v6cuM1f
WP03Bqx47pFhK0fZ+wdKf8n8iuisMHHHJBieSGD4PezMrD0pMZsrYU8iGgf/PpY7dZO+/+LdzCOF
3Y6WWIG+C/6L5/xfNnl1EKb6qW3iM9VB8vLLZG/CnhzvknI5FyvEsY9prHysyw9o4MQUmSo7NQ27
JhqGpXXGN6CH4KKQayMJkTn/pnyrUuVd2vpX/WY1d+W1aaMBxT4fOt5qLA45sRcgi1VS281vMbIT
1BfD1HLwrcdvKycclofBopcdPY2WchfbC98+anTvhJNPhnNafqaSsfNknyT6QYKARQI1M55GWkv6
7wm5vmSfA91VRwustkj2qAUbVqZhwirUy7D6FZ/WLvmpWKSupFU+MuH2w4lIlxuyyRLJ4+Sb+oDr
CwXeQdJ7no1c5L2YydlnkYQec50V13XPUpNn7yGV1wsx3yuDghWcvRPC2ShBfyZ4/tNiVEvSknG7
aTVje6v7cfs1MJUnXq4G0dvUYQ245/3XEuVVqBNkZugvv5EyjLJef7aunsx71PmrqGHdm8F9Y9q6
h4yMklANYTf6P7NjsEqlU0krfrymgopMbL5dCN8l0yzXupTr+NbsOaSKrduL+H4bv1jgfsIikoSs
S8DHeDTgT0jIIqXoB8qcnkhmXNzDqU92A6RT+tz0oXSNQetKIgCe2SA3S1mv7mH/xxFf8i7xkrUz
5e0kB40ieUmJ0uDPs4CmXuC6UPU1ZjsmcsQIGimCwp93G+jnd2ePUjTHDlJnmJSb//ah31/28TjA
egtj0UgoMZumeZxwOU3WY3b01gn0qR1nF3t3Jm/x7KRZXCFpk9KK3w4QYJkYuv5dfG90qU1uM0qa
7Sg0lqE6cP7E4mjNxV7JB8+/MfnWTca98k8JHmkqsdErd7PRjGMO4VcxdyMyODX2UYzxBXi8b9jZ
NvtSFQr96VgdcePWj6WS/NUckQvjM3bWt/+CfNcxMpTaG00J5cSwDyPNSHTKpkj4QTzHbbb2GRfk
4vgjJdnMroilvVZSLcNpW9UktRG2OWMboIyvgpSWGHDQhHzvzTdG6jk51HdXvop9msL8BetWHNjj
Hh4DTZuJykReYmd3m8UMgTPhTzp6eYbXAsnCo9qQGCmkV+/YFfdJpfPQKwTBtv5uviO0/2//KYeY
xzEbmGutDuoO+E2I+9afB8ZIt2QTIkaOYxNU0KzL4KSv37YZMej+yZR6jBW1pw7e+cBO/YACoSgy
yg+s25rljTNraM1wstABlXZJTCwpoRwmWRhVDMlPKoHlP5NJ/2MoBrakkfPtBWTMyNH1UGAFyGlw
A8zwPaeWONh952IFTeLJUGwT0RV9V9+AcKTJY1pkMXImGjL32NL2obqbmwo+BN2dq0RMOt+ht7tw
MoECvqpvp09zR+AroinZf9XFICnLx1rWRcmQL1up1gZ8jGHaQHcra0NiZeTSl5JozbQwEvgrKLjb
7fxa073GLlRG1oaK6yT+XsOS7IOxMY5yTjR2CZ5neglATa+YJfmlV5M5BHAQVcrdls7sWb+FonVw
ugFaRWs2oWt+q+BgINvx1Dsi+3iPdsPB9BjwLyqLxShxiY0Hg1WUsqKqM0xs90lI+wwMS7ZApmnK
4QerWAK0F956wnoBqdBpSrunELOIdJi2hoTpwZuUdibElUzJo8cQgBktwh3fVSf9g+63tYh6naQi
VPclzp8UILbOdSe5AeYs3Vf1dSAVxajBTcnU94ymOfCcVtmD09z/Wp9KIuNegl2fHMikbn5Wn6o2
cDoYcjlhW16Lm3ZdwC36jKyW+7+TdrMUk9AFMugl/7T5xiRNiIpUPiragZUtn0OCYy1+A+cg4M//
K3rUFJtP/dByaPaDRMx1FLXAnu8K8yiz6qDlxUcmK1R94xArmroIJ8gXybsuCb+d+bKyd6e5g+mS
hPrbVThjcQtbuE33JOA/FilvDoq+iGRdTmAFo7MdPigQWS8D1mTZUWQwD0g60WOL7MXVwHa2kBtc
M7e1SFbzR2AunjIkEui9lv8EcXN4nk02B6lv1mJj7pyUF3GIlIxtbUwDf3SYuAzjJt6DsndZL82l
9qOvhOkB6FV/Au6vqyfL4iUiik6SoKr9jSCjpAE9zrG+Xq7p6R17dTDWXhWrXiCkfjjnBe0yVgiX
D8i9HfRnRJitut+pUVQHuUcLyBme/vLaLnbhmqjcr6/gAxDckeROIyQ2kTD5ExCMhvIovigrxC3k
4yEmxx9PqhXHec1wXGGZSXpQtArlTmGQUgI8hKXPmpYz+J+nqVVKAfq+Nf4nQ4T92OudXOZx8Qw6
CA6C81W9H5IgjMATYqbpRTRFHXTJ8zcJWKAgcZKCgwIsUl5jTnDe4cJthl0zs8f+YgGlkuWOlG0N
EQnINJmd7KDRcHZI7wa8YlW97kwJLIdVVKyatGyLdmY97VFU9EkmTASjNoFqLfSR0G3is8VrFo68
Mvn8oFKnUaK6wCtR3CaJ00S0KZxBVHJKoagVnezbwWA8ZeIMSZ9aqekOYWF210o0V232F6pUW0YG
aD38w99adF1nVa9oV2Lg4MMtKmvsRNSVoKXKLusGY14zKbQdzESNQmFa1HNV0uFWQcpaAVIVaCEH
UTGvRXs+jPI2X33l3E5ouWvp4UR3wXrYyMfML4jWmuvR/Yc6Znmrz56zFIZ58vyqPU/7qiwdnwFw
VN2DiovluO8uJCjX8f8gmGDftgFefKOkQ/7qE0aSje8BO670sNdm4W9/t9B2cu4lPp4AUCeKSQyh
Vv7JljS4LKi+RhgcHrK1P3K3MVOiZ9z23rhO3TpmdfV+j1sMI9/5sqTGZAZvkkyI+OODfQh19s3r
SJkEL43B8ehivJrMWOGJ/DHH10m7/vdd3bBusQIcCdEEcj07HMTqPZrFOYJd6+Vykg8xKRWVUgxx
vgsPhanmNUr445q/GcBCLgXYsBeY0sW2Cmmp6VxSK5Qo5vtcvDQ5KwyMgi5SXF1GGcLpHpzVHuB8
ZzDJsS1mtif+7Hz4RA7cLesosxJAjZqcJ2ekGQskA/OeYxT4BR4rUhyA0gJea8D1xhgPn99sr+aY
eZmF0BcTe/uF64uZqJRpSFZHOGvrm+RZKhlJNQCkx3lmnqd62tXC/dNU0HJjK5R9H0Zv9Fv4esKz
ArxjSEjUVyqQsKcL5FA/j0m4RxdI1PmwJRfo92ZigOGtMb5wrYBHkeEg4mhIv+8je9m/JFh0L/UE
SimYPctUrYyT/P3vTlzx8rpa+e7wJ/5lUzM5DhBe6BRt42KRfmoKEqtNu4ZDAQa0SOItfo2vDVbP
g7kXUIh8f76hElK2wlRj1UUgCo19UGI/qJoI/GtScXD3F4svMSdjECR2ha6q9VC5YMBlbYHEnXSg
sVZSxwhkXYQwLw0N06dRdiY8nIlmampEBH9PHGcLsBTdYFtLtbT/7gX8ZHv74rExdHrmN5lhL3Qr
eZ5izyi3ZqiLudyYO9ypQLxTOGVONbosOPqFiC5COy1B5sbXrB9R/BMlzDRlNgGDF/qdzozcpS0R
NDlpIaxyr2/giFkwnxnWLoNTyBoacIm7rWLeffCy1VgXB3BmaePdKNIOOI/8D1jyM/b6oqNh6KbI
K+6laGWOLjLzUkI3nTLRb2wqgARb0v9JvN/RBDAG4dGDvsH0ZzsX9lRzVHg9SNpyx6XDe3YO8u20
vS4yYZCdGfuDRjS8Y83gm54AXmrB/OeUYbI6Hu5W6rmHKjkLbpMOeL3/lP+98vTO3HA5eUPelTWy
alk8YUsKfWBo+cN5TRBhxbRJ3XjbMP5mvuhA/omUkkqVRXJgB/aY1evCOqe84iWa1xVL/m/eDspw
fbkAR3ZKyMuXvnHVS5JgWNTiIS+G0iHqMftwUuuV3013WX9CmLGPwx43LxPfl45bVKBOWJ+t9GaZ
j5Gn4juF8jaoyMUVNA2Y9HyyD9OqZ8cguP2mYYLY5pzy1YF+Xxa6LR/lAKHWbkvCoGLFUHobEaty
2TEzoOJYzmmP7wejb0JETNlowVRf4/JzEnN4qFZ/0K21pOo+uplvr7Tgiy5xKbTE3e/1lCxzOLp/
69lyMe08kX6H/WRIPmu91/ePMU/DCpMgHI8cT1Kb7cMpTzPUrDORva1dsLDZOkcu5D78JDuAWwx7
tFaCCtCdUu4DB43766B/d5dDaek2dMAAmGyBZ44C9yKy0EhNFB+gAptwsRJfPyxRaLE/rmxfkJl5
QrwoSZNhl8pS5BrnIO3XlT5LoFhyhXcD036/8YF9u/tw/Y401S2m4kh+L/qu3TJYtTRgRQKzEWY0
l/cXY4a9oFGZyyyA0IaVu/z1sMXwht+8d4AB5Dfcz/28PoUR5V870XHh5c2R0plYTvx2zrbrShHa
7whxlz4MZRB7h7ytxy74al4e8GLVW+n3RKElf9C5M1vTpXrnT/SR82WAgYEaJg0LftHOdFFhs48B
Qb1sRKndSy18ANDBFQSG4VgS/JWiGq+NUcq/F3F4O05E4Ls4NCSBgkaCSsgY0OCffJqLEVogZp2y
9yHz3mfUrKC/ezeVCi88X4k/tCrF31Vp1/4+vOk7pMbBynOPFDDE1rA9cE1+lf2gzitNOHWPQG87
bfyC5OGB40SsmggsYN5Qw449NF8wyzXQ4vxDTJ8DVPU2zaR/rYt/TX0RYd9XYBt7y0R43s0frF8I
/3JbJcEF85An5ESeK8LGOOfYKYUw7XWbKI7a6ou6lUf/XhXTQyi3htFsFvH+XIs05G/dwcbBM3pX
uHIfqb7r2MnSPc8h4pv5OIuTnI1Cl6zJv5hStNndoxS6Xg12+A8IVqOGKywuqu/db915lDI7FbUJ
kbRHjRqf8c3dfMYmnHFxEi27/BUQbgDd5H3cI2ss+9/3E9g1M22Vm/YmUZBcwR9A9UTpKtj0sWkD
lLueyEHQ/zJowoO/7WALRw6mSM0nr0HV4mCDEMlUQcu5KjA9r1NZPe8sRm3kdEFw7wMWvMrIMDR+
Zw6axqU5Obro1l0e1YIGPYnEEW9aQd8D5PmIarDGk3o7gLbE3zXmxhqsx0I4+p0pzu1G0sNBdt4H
ylWQTt+/Xt+xkBs/d5CJL7KdQusvzbEEchucM1806vDzM8pTZZYMt+YUPZ2NnoHWVzA6KD4Cf8Zy
5sT7vM5LmqDwvO9JM2kIs5kwD9JSAGl+Lze3aH8ja83GQuPsoSEGmAY/o6jA/oCssLvOSiExbM/7
TE/Nai8nM/3sqVbFGTxzFvb7ifAka3sunjGr6CporWBUb73rbvTwSFPVNnjgexIz1E65/DBQ2nVb
mCR+/n83/wifNdu83V95WU9HhwFVh6zRYRGjvSA86IGUcessE24J4c+bWSBcca1S3DT2mEucWkad
PT4DUXb8K1kYpDy1DGme2RbJGZBqK4gtdenISbs0xu9cblIRXvnnDfBV1g4FxltNyK8twSad6yho
F7EHXY3Bs23V8XAdDvrAd6oR+37M/9WXAqIw8qsMrGZv88SW+9FVCVMvlD/LDhKtIDUliCnBYhwQ
ZgeEBncR4CXthxub6XRVvE+u0eJpRn4LKHTrTGdBM9ANsmiUEXSm+/AOKfPliutQ0sWm9LAEdz79
SAAgYIggp/ajt9Em+ikrzlr2Z7IidYC8HFl25mcoMs8J7EbKieXkLjgo0RmidRFgoRJ9/EZYYKFD
zYhD4GS+3rYkWRgFIOV5LkP5qN/Z4yWzL8M82RKk1zQnc9egmzhycExU/sf3bpNFXFEmgNcPQ17A
TIezbZI3OjRzTOUb2kyM2YRKAckhaZaEkGTxTu+E5nyAZ2NvZ2mpNEl68aG7kxIkTR98NkcAgSFy
K9erv6g5XtSenPPixor9pfEr6GoHBpV/qK4MS7J4jFRcm0qXOXiktAPgt24YljCE4Nga5hLh/DU2
lyjFLIESsbiwc+SGoi3xlN8grbX0RCQoiaIVBN3YB7Vy0MccZNKlVAA1m2wfdoA8qYpFEc9H9gKW
KhsJShrEdftUeis0/pvqDLj+uua/Fg603SNPv2gXsGR9SeHnI6pUx9Ks5xg6+sC2+Jica1V904yJ
lCkA909yipdfmzpZDrtGklmMB43mo4clONJdln41KKgdGLnu1s55k3XgC90CT+ghPODJ8jkd2h/p
bTth3EbOMMYuI0Oi+Ky2rZ6nES4CYlFkVX5y7zJmPTPkZLTpLi6Rri90JwbbnSXUQb5dSDGP5SdX
EH/umsGEV5o1jYU7+MxYYYabaHocmbe/hI7aD92mb9+BZ34q3hhBxV361J9rpcFwnwenTir3UEHo
uVypzAwLGX2yXjykG4FNQNLMZhhUr0Cs3P1nHNOm1Sx1Pknuo8jt/dzNxTpariY1ejQYWuvSN/CX
O9mK9tf2SATRMdOs/rzrb5tSU/acBFCFJwyH3e43yLISGVAMKH/p/nT44MWvRQAvVQ//6gV/vtgc
8B5+ZXIfz2Ubqn/XQN1jql93Cqjoa72nz1tpKgSRYFksNYVljHwrY1PJVvd1XJAiJTJU9enVBbqK
AvY0bmVFBgBNAxttWO+Ycl2Wy2JuqKkuHjjtEfsoG1/O+H2W0kVsZADQKszDBVsfYXv/kY5z3Yct
NyWRP7hkSkgSlmSiAO2xMMMGgS0/jKQf8YKDK4niXtLBBK6+iDRqlBqUpUsTsAJiHobGudhsYypp
gaI4wFWW7zQ0Gy8NRwf/hV4SQzYXUtWZn2nQ8y+WT7PYUsfkV+19US0q2Ak5292QvnHayemc9jGQ
+6E164NNPz7u5zPzCZaeKeqLZxceH011188l2ioNu+fdULjyxXEFNjzxfd8FF+8tOS3ZUiyI8BrI
Rb/ShmqEJ15blQSLvoYDYgGpKvt8wsLlMpel7YPhg24qUqIytmJ6Wh88recMHc/sVJG+Iq3uLNp9
K33Z3h3nZLdTiVm0k6GvD63BjXp75ShCO2LQr7fr0Y1Z7x33VL82jmm/ILDcDIFa+ZoZ5ZrlNua1
MYOVts49A+1OHEdid39X55cvKR5bGnCAqHKcxsK431d3y3fCrPMrddxq/PGUs/N92M1jOxV85CNt
sgJmV9RNDTOSmf+KR78zlqaupYucgiCE4zK+KKEvMKTzCGWEK5Yq3N7MjzEyAFEQUbFi5OQVkkRQ
v17Y2TY7IjkGQQFpCi1kWr0Ra5TBf8A3jt6MxblNQJUTNYyoPBZs+gRFfdq5sdAJnHqPgbx/QuIS
W3v67SDVfk+yEEJwzTipZV6aPqu59ytr4CYqqiPkR9ytD51jXC/Lj2vkBujOiTUf+Sv5ou+qf72e
oQjRaag4kU6tur6ZdBle2qZOald+S40LJ4j+Qv9qmyOkNoaA1YYTKSwRODxj5UJ5Cr0ql3a3x3kR
cL4q2cFB41BvJ5MFn27p6S9NsK9QKOvklOOPomN92yt3tLJrCHmOb81IpnK/GND1yYNJzoD5YGaE
wq5u44QIpGxOhuUVDL8+zqEG2dEAx/+Mtj30MSBvevTEPmT/dsgZeqd6MRxu6KVPLcluL4qLH/Ow
OmoeEzVuAzR33DpxT5HN70/YgZZ2I7r7ksa1UnLfWaqjPz1rpCMVV7v0Rlp+x3ev1XH9cEgSv4dU
o823iMcLdJeVvhfv2IlbDTaY8069KQoIGVDRkCV1sakobsmsY3uZbX5F3WxERn+gtEPX99daeYAC
G0n8QtthysE0JvIHzNPqGf8AcrA1ddiQZM5mehU1oq1EUVBClhm+vaXDPqIo7S1oHW7WgrOcViwN
XsYZnfORdr4Ig1SqVKRn7mwWrX9X8/sOM87pjNHGf8porqNia/WNTbrTlLbNmFdB52d7S2cqZ7OO
4t/u/JQg/eWM2s4/M9SN/r09bBiYAa5dez8tdG5BPLj+MUyYb9VtCUlIkR2N8bj8L9TsOI74v/6P
XsxF26N8cvVghGSJk4TK2JxYTOUApedXCPTStw5vqyZzGfDfVoeZqwIocNS2J+pnZ0rv9YMBByNo
mtZJqk4sGJIBnevprVW7bXMeHemy7GjIB8JPP1VKO/U8q83+5CNm3oDamHUT1KyEs2LI06jDFyNy
mxpFnGaVSM0cm5ymr1FmFMu9oU3swHzy33pq8/luUXJSIkPzYFEuiXeiN70/k7kWS7A+wMK/51GF
a97mAVXWJmv0mDZwZMBrCfB26p2x3hEw4FBCYEuhiX4XlzKcVEp0BrXc6G+iftnd2rn5iW0WSt4y
1nphNCs/KzPR0m6ZlVnErNhRJT62Q29ypi0XdNCDwSfIGf4nTOuDPLNRf10zRZTmplL9qC5tYlHs
p39DAj1PeGYDKCrEKIdXmPj81lAfHkR+mRhg00W6YztbSPz+n3/fqa8qAytiqMwsxdpsDp/7YnQB
xC35Wz/tizM/PVYZ9V/7JyG4mjorEbJP0Q4CEuXboHtpJA1y4Ct/Y79Yh3qICG0bNxXrQFEf2zau
3F0xJ66a4fnnLikYB71Wx7yFxGwqx/H8SFnPPdV7HvweyUdjgsGKPIqEnOUhg0I1UB9ic8vYGMfU
u7sAADOAFTatpxim9+cOWBvWb270AFqNCVxMvfj4gMBEtiAKoDbid8ried1S2AWjeTLuthF2cMeb
pddHNW1CC5JpCRR+uSttIZsnc1VvLW5qBV9IJP3d63wa1/dP7QkftZubM6jmGIsO4IeZRJZc7erg
ewlO93jvvNg2xdIDH/IcFUC+fNATZxfMPTfhMpLkFISRzu6Pm6JdKZi3uqv5czKmeXsKL1lylXln
Lj2eTS3aJsjv4dFod5vIBUxTNTctiQRDK8m9ASLdv4kJ7o1EIfpbDLBPGrF90k+s2QvYNXE5BE8w
BfQafbZ7r3wLdWrfY+BniXQkjNzbUZGrW3a35r+Yy/Kp40G6X2vn7QgDo3xfg2d0Jtm5aNHmKeLG
dNjxeWZa0hQC+WqnB+4y2a7MY1E4lUVcFJssOvTs1HhMdedKyrGepiu3poZSDjslYgSeqPODkEgi
QR3KQm1ReIWroe6SQcBrUJpJVicdzaj7WGpLVByGPtzUAliJHF4kmeuhtV8FfJMTSIjQS9p3ybRn
ldQIn8npXrFPe9W0gMWf2OKhmT51+Q4gM3wpDITZYDHd0to517v80iwULaKnhPC3dMr0F6dxbDFk
BmgPqJEJmAFKwN4aMxKWPdyH4MMR5zq7ZOWU9V7eR8zNgvZ/Xg04gT6mbgw3k1BKdEyOI+d3z84t
Ft8BoewhvvbzvzW6C7Dox9xTGdCC5PZvV1Wg41mFPjrIoxWH11WcDDh5Vd+23eI0FSUtHfZL0nPr
Yph2nmLsIWFn+l87jcVmU6DXWfX99Y3orugSjO609H4pg5LKwr12c67xNmjYz7APwtl13YzlHpHU
0YDnQGbn1klOsavaXJuUXw5LGQVkSuYSj5jEyH8bXP46c0BYLCa5grl4759/XtlAvX5PSseS5QD2
/Vnii8wMCHzH/aixwukFIy20wxtFAC71WOCbPSNQ6Uj6sDmIXOsJbL6ExZUchM2dQCswDoGVYjid
PJLwTdFssUACdubKNxjqXbrhVKsznR1Cc9/WJh6rlfvEPpOtUV+9bViFUlqafzNk40gOvcgz8Nbq
BQ4IxFXm8xEYk/YrH5I3LVAN3TPzDvKpHUHx6YVds/T8ohrwuqBLQRALR/uvzOt2BmTBGM5GaFtz
YZt6U1Q1Ri1XQh8422oIf0qKOXRgubH8dZLt/vYUUsN53I4Jt2jjc051nSsiIPG0kYRWsvxWHxAf
m73STk7S9RUnPjQNsKnTH6kf1I1U3WLIfyDjk1f6ARxsqBMUS5JwTzakKfCwxReEpqVV2gQRHVOr
RtT1tPPdauZG7+E3qbIkXumSjRRP4a4rDF/79TKMF7l9vMUv+1juupRCZTm9Wbo8ayI9RhHu3e6Q
uhFTvYNxpbQaldljyp7EHJPQAzvgdq3yUrK1wYcn9CHlwg952wPW9VVJi5Ro/47skUwcG7Z4Aq8v
GCy22EIm1Qfb31kCVPehVPj7d/tiUGvntMUTGjE7Pxf4ox3vp2IabAeQkmsFCQEX3x2yPwtq+KkV
AVWFBA9reWXQWbgXjMG9xm9D4M+I7uZz2bn/uYAluveycE4ZpIm9y4naPjYh7FFXWsKoGGu+usJe
pQePVhsq4sMPiBrWtlYyBe9K6IrqD4quwNzaEcQasPr+eCD+JT3cy4DPszyTjFXBe/oMZmWTCXUb
26ItS8muwvIMn+HTj4FVf0u/Y5SC7EqWzihVuG+oN+N4bu9nCmM2Ze1ox4jpC1kCiYSGloHZmlcD
1q8+uoDb5KwBU20uxeHHsh55OylJvBH7cnXtYQf3QAz6kQMA/uJdnkO+7HD+DX2T+BsyZe9p2r6O
E1/UO6ovJOMEo3bXZBtjosTb4r2pRccdin0APScbIwmbWEfZ6DdW0rIbLlCrp9nCtXYDANX89umy
fe5QzoK1iwY518Z4IEO8gLwCNKLX3ASNv2KRZn/oii6wI8qTy+juYMkZ+b5ZvIPT/8MoHfKwzps6
pMbF0/qCaRlDU5vcUxFmvI8qq9sofg75PLulZvzpPJcmZoe0bLAK2m0E748bGNx+eiE6FGpaenlh
Ox4VOx5fGDokkdnpzjQa5G7tmsaWsXesdMfj8W1L+pD1d8YBtC+E5474cPQ6jVmAoRPcrUaUEFZv
TcYjJJ8jqnxwcpjV2zSa5LaQMSZMMPoTYzX7VnUC8vKYQ3JYkZT215muRhgucVwQhSp2g/PL9LnS
WKcHU9OW3A/5tAD6yARJOl/5RmVCQkMAalDVQz9NiBBboDwphnXgBjeH6916MDnJw1YdVaKqc1gE
eWl24R7yI3zLQrkWNALRf26QDsYDh8kBV1S9Kx7DTpUIuSyiVnHxmfjlSYcoxKzp0fwPasM+ZlVH
IE5OfUphxhCWVpE77g01qlsbGwBGnAxXfa9ONUuIJl9HAOhGgqj4ElFZUhillf/EYvtr9IoCNX5r
zvYupaIEXLEUliZNivJcCRTNoVUSBiSXsQ8IOndSFyKREuk+drVZZrZ6nQX/kWnbIBD0Bx4FuAlk
OSHBxvJE+TPGIGedilOCllXcWJQcUvR8gMZnndh0mVcdFAsjArA+23ntsYdwGdmWcIS87qalQFcR
K3hIyWxt5A3zCo8nWDQOd27+Dua3SUla4T6U2oCi/yAdPJ4U5QLpgz6VD6SGp6Ld51iV37SKUKtm
SXiquQallaIrlLV76IaX6QhYpitUFfmb8lyGPATmeauVJzb++ReOyc2StblZ2QNb1J4GxQBDcJhc
cV/CYfx3neFb83k+z9zTLS9PvXgY9U1wghZcQ+ZID3glCJE5S3PT/BsIySulPbcxKF+h5qrh68Pu
L3Nbq6MVRM0ZqFy0KiRiIDn0fwlttB7Knuo9yfaDO7qiIctVCr2wPXNAhxXtK03Hd6XswXdpUaPv
mozwU86VVwUkBKDY18osienyhqMdk2riXRLqeeOF1tI6EbWXeAppND8uQznw07d+y7FBdcVzT0mb
uz7mNO2cHFEJtJJV+MERENbRyHqbQIsuRobfndTiNvojUuloRWXf0goXSX4xrM/VfpqAAV36nbAc
ZGMohOZezzRfcTjZxmXEjPrJrIF9sGKbQ10p1l6DC+cBmdB8oBhJBo6n/YF4ShOUAUGwfsI3IpNS
n1h1hVcXVpipRgm9JJXetM+4gr9d65BpPRmlrPrzHMOnwD30ITQVFURnYPA09BCvBAfqGeippOOA
NDSZytWvSxZXv1rVreGu8+aD5vKID6ezlfhwD2L1d0y+AwgJBEPAr3PJLaRS+ggql76iKGIBarap
9SR922qzl526Rj1/6SMpT4ZgjmdQ9tfbXQ0CAkNhRk7lI3iE39iqp+8khFnReBUJzbdqKMDUycfp
33wi5NpDNHmqWH9vs/avWYFC90Zn6IRAOu7XXjH7mj7uw4B4WUvQlli7I4RPVQhpKHSIAjxZ8dgV
J6mkYGuBWA9UBKPgWgk0BxlXH79v6ZDptcg2y2YdosCABKAmrQhfVIPUrBjPtmRtpEq816ht+3Ud
mpPV8pVdmYZNlWXL/dWv4fdQLaerWWsJwkaOuSfPbKq0chUEdpjTz+EMsCqI3lcNJj2d18iEhZiZ
ns1PX1zAb+HjlMRMaCa07BB+QjNPZXVAAypYd/csyCv/Th1KncWz2Vtbsv1znSqNw63B81gWngV2
2Y5SCHaOS34wWqcfGLOQasgpVvlLv6J9guXmrxlhlSrAVhvtcYU4V1039nH3LkWrNVECK03KbZHx
/XrnlqA4IDux6cBzowCaDJguXLPg/8s0ec9TeuC1Jv8Hu8Uvz7gTHlsbJRD/iePFaqc8AmJBcSin
/ZWFxuq55jMQ426AyNupRZKYFFBsrhsIrcYJtegDFUiRh8FTVrmSU7h2F2+Z/D4mLeLx9kNkARHu
Itb0WbYDoJjyNMmuimN/7d6QXZRi0gf3M+UMNhswVxvUyog1ZypWHklr7jiZLPQyZlFaTMpgTBUW
S1OCAfF0Ghv+Vs0fUNZXs8nNoOjz6dncls5tLCGmCV3R5xnS0J3p8Jxz+9yjpoFpWch4T0yMGMSb
KfDiOk8zYQAfIGOF/mwrAK+hoWOIWyXxtolQuB8LGjFLvhMkjw8BYlw6I+uWH7W8J65JIeYRdWEl
5jusrJR1yJd3AiXlSa7XNaf5kRDh1l/tNFwcG207l8tqi9aaU/3md67lWa1FY2xKU+NQ6eHenS20
Sd2PfCtFZyX9FbnZ3vY+coltHl0HBeaMqqknO/aHIjpEqQCeXEbmk5GvlOGzMfc+2zNSoyK/Lc/t
2eyE6nvUFCesysqtYm9Bx5wnemysYS1SgwCIi9iqG69boFCNCJVoUX9+zfLbRY/yRKFoeGR0dT87
BNbAtpMVj0oM6CPI7dzhghtvpAqzJaR3PMlmTX8JEZ/8g6sf1c1VA7rlsnD51locbEunDtYxMHfM
VSDp5K2aK2SQ1eIFaYUK4oSWJSi/YAyABxqC3unUDg4Hi7JJTjkppkyCImDJgpQc+4sr7+hNA06+
Upy0mjbeTnldKl3ytWNE2rsDoqymI07geMuaAZssbLaeTU55sJO+cHWM401YNaFInF8TBcYyfKoe
U25hRwAI3aSmbkVTkWtqYfyAnCxFQoH9AOwboksaacUnKZ9TtNR3WLnaVP9ABHu3Yj2GnVjf/v4p
ZwjWblBJO95ye+Exep2G12J6VTpPRkH6ArnJPfepee5F67f7UoVmSsfxM9Y9RXp9mAF3u6CxUyac
DasqZSsz+XkAU4x2Xf/ROr9bxvFNevGIUm50aovaCnpd5NJIrgA8u4DBSxYR7agdGVDHQT7yPVRX
HYL11hUOsC6f5ZtN8640husot5A0FKcQKhlueu5KmzfM+2GIZUemjyb0Wqf7t0YHkLXv2m9fGuBG
4PaepoLotlRLRkiQ5pXD9MXy4TtsP2WSV8yvZWVFLSbI3hFydxFHQfcutQkKZgZVTqt/W3AaqCPP
acsrK+5y9t3tp0DRivhqBGXfZBvmljUCXu8/hMW0tAQIEL6+nqNe/8DmNDS8bZ3FxY+Oy6Nh7F5R
kt+ZhO+mR5ktShgfvqdS7J/NBKTmF/Nz2Tn3v00yc5jI6EbJfYzgypHhC5mFTAVRQQhAp9FS+Ak+
vTgs3WHxPMoAlj4FTogx/OwV6FyXuMHESREsIW6omSFbl5TBYcENEbiGO+kXibj5ASjg2NWl35nN
sCLFL2SDP50D0mUrX/6lfbjQDlp6wpjb9ycK94UGSZnsK0CwPd9eTM9UdeVOaGDiieUl/xKvjrYb
rSw21PtiM0a0eFT4Zm39LHDvTM1fde3UFdfH8nQ+02TVJE2ELK/YWyJNBtvDVlrPl13sc3Qlf42T
wfFGGF2K09Kl/AymQlqZ6Fb/DdzTIgtLprbSLm/Sg5PgiJBjCWmMV1vZLA6kGRPfiuY2pGeQNVRT
Drhme3uS1fDRWioKZ8qI1f24knsNWcZ8DvjH3ZQ2d5Azveu1jEMDuQPdq3YiphKEvwFlpB4qX70V
ClD3nClS54JKzFvXQ4R1g8VMfqHw+Udnw0KlRGqOZ1De0QWeQtMvWFAhf6cbU6BondniYCABr3nt
JxEP5r+WQxo+N0i7ZCl+X0cFU9UassxM1mmR0VY9lhYoGtyhEPowQEOSNAFp1mupM8eTp6J6vOy9
wp+Zo5m1EINU8DitAv7/6lP92QP7qGRfIEpaJhXOR8dF4BSZ9oB23VM0p6gKxNmxUl81ch3F0ruV
7FfQO8zPspdYkqxWQcrMOegGseWL1T2itnFuzjwGay6c+7tbRXnKWr8/w4xtTDkMc7Ie+YpQY7BH
QR4HTUwFqC5lHkvUob24XP2zuYga4n5MW2SwcNAGWM2MQIxT+QuruP1k9ogY4rN/bAvlfpQpjTEI
rhctptBQldiPqlhvfI8Cq1FpLRMscqqI9DJtRGeqHbTI6E6lvNoC4fOdU7CPpIlbIUB7LCNqblrY
O0EqMcRBlPtFUgpKmzjBmPyGGcevwE2aIpvVLwenwsikfvgh50d89dMreqS6pZPJgGX3lIFJp9wH
Ni6UUZ4nGi7Y11CLsdr/Qe/AnkjpSnk+h2IGUkB3gq4z5RaoE4v+Be0Og3S/mccxm6sLTvTgVepp
mxvkh3zS6JtNInCPV/dPff9d/YemnPiEW3IOKiN0XBtydfC2uJ+k0ULZFHTEQuTQTR8lH0khOVPo
ZQmNsIE0pUtI98/t9W0WDtgn01/C6hJmnFhqnGE4PB7scDE/pp+6gpUnOEOqsgQVACJCM3Prl7kb
1gnc/iE7sK6oEdufjcnGKri4rQ7qHCZpBMfx2r8SZNLqFWNxQDa3QotA8SFRQ8chnv24fsemvinN
6OEmyMqSWkyK2XnGhbWhOsDRaktBP3mR72QZEQ/F2MS8Qe4ikR7amBSx6JCLlCKO/3FINqCp5/pg
Oo5/HNR1FU2JKq/JlgaiCp6azMwffRT9LHq8Pwd4heacb2psR5SJ2oPg3H7GBcWxvOEq9ERffSkQ
SGNeQSfpVZ6Q7LEGeKncdx1w37U3OIGBNzmePCNxlVqDGVUX1FIR8dFetyPPLYF6Qehjd9dUABTT
bvgTktjPAFkd36u3Na5B9XgNcZ5LdiO2WPpvZWOS0BcxFilmDgoMkpLPH564/27vKyeMfC0hccHH
jCMsIBuiKqUupdOaD2XrHOiAujTx8mBvlaUUOUJo3tsit9JTJ9llrmKz/dWHEtv6p2Bkv5nycdeJ
LFTgsQISz8oaozBiZ954+tjz+XDQgtREiLmIMxyMgcPK0I4RQXIBBcOOgphcxDzVHrDoh6aKCmFf
y24MVy9Z33CuuE+MuU54+4x4gdhg0MPdHUvnAstl9inkGMHc7bgRMZDdXYe98bIh0C9X82hOSxp+
Xqnnn+/mII66yTWiguHUnMxKZx2b99SIfO4+B5GrRPM4h2M2il6J0dXNjlzTAuVHhGR90/lk0dQe
LvksNvxTn9/7DQJSuEipSRsv7mwRNEeygiPkB0jOzUMEqSitCqkZG5QD5P/8444V+YMGSUuiw9Jv
GxvHdlVIvzsQGTFno+H+OvihnF6GFeIWVPESR/FFMgJ70HSGs+QQ2Up61zVdMbjO5kiNlpLdDNXR
A1vyRlv2rX7LeQYu8JEpt4V2HKYySWRc8uvikxPsxuLuFpOJD4TnuaMG54syGLIfyjvLxWPuMg9H
H8KrdWLTaF6xpf0PQ9vbnz/kq5DHMoJ5Xwgd0wvl5eDUZqWa5xEo6dFNUZXfcyjTYKE+LN7h09wL
efXunk31zlz1uRdHJM6bJhkTFXYvtIG56b4WJuyfW/A+q1/R50LcluMPvnIC7SWhRYRLOghvcK7B
FriC1dvCRVPDYKFSCnrwYjMsV4nGbWve0v/RcEd1y2MTRKAjaRTdoAuNkJsz1C0o8S3MRugAQ+oT
yD27pv6pXwOXioyuk0XuRL6r+/1rwLx8OsHxF2mcemV2h5ZrbcnqUN0nwIxKA8DZEt9xgv80fTP4
+hQCCdkGrL3h7aIjiVKpXO3NW4vZgzc1bWgrsSwak5BetthZ5t9pjBTuff4wKH/JL+NoD2QtiGve
8/yqZUribDCQ+LtHjt+7fQ9MpDWMLJEa3Zr5RioWanuRVujCqHoz9w9rt79PsCNT0FqUT54FkdTI
RV6Gyw/ExHkvCmbhnRKM1uddODMYSEziPzhPWGen86HlaL9qlHOMLqXrMmTt1HdE4jiQSMrLn8Gv
Zn+UJ7PlDcyvvPB4eulW3qp9bDzxdO0vWJRacWR1K1F/7k/0//dhVAL4hPOpiVZQP058TEIYjJhF
fczmV0JoNUYoQ22y4GQc9XINCNVLB2lAet7xiPu57fnsM7q0P5WKyvGhlORINi+S7Kwp4ELBlMf8
vK2MIq3Pqft7tuYwKhFdNSwhzOgy06OSz0AXfNt5VxrlImxpVXo9NEkHkNzhSFCCpcO6wWTAIvrj
qW8ZfrnKboB2zQxitgV/r2HE5q/bP4NcnfE2UCAG+VuDSZZbC3llSUP1eZFJyUTv3e+0BvklTH5/
HNgX13tK+LIHn+N22tEd9kWlc3uohbblWuxONlS/wmgn8gokXSKLvghthie+H3YWA4i4j9TUak3M
mVTJbWxYPo9p0+Wr6XXxGYoWhsxAiA8hbExSIkxau++lquDK45wJlwf5o5CWQ/gZsuqYFh9+kSRD
1dGhuRRET1CRbSDvSbEnYqZrOSQwmNDGihEvWp7xvJ/AXTBW9yaHMjSvZfJrjQ0J/kGbmRd3Q9Di
SQOfSca5Gk4JIWZJV/9rluZTpoA2FJwarL9glovzbhSVdhvgjew4uC/WEcqu5YT7atBeMvyRsSVH
TZzRV4nXZAb8/VqUr0Nxiv/GmDoSoBWKrrF4GmJB9HIaeaYRVj9FC+asH63Kd8T9NNEFmqih9Bkx
hcUhINojAIgtU4YideqzUHF0tWdqNkMHM7hqP0ojlx/H33pdYW5q+2iiMbFQ9RnsMSzJKVIb7aBz
YgFFzus/THMmKxFrm80ZaDmeVxBFco5RC5bFBRoLVfRhScPt55aYiNehivg71xLUdf5HG1aFYJ4Y
yDxBZMNHTPDdur1sJEBPD9IQUUm6MjY720O6tu1JnT4AUDwaBcARxREK9o29dJemLjHozBHvsdy7
C/k4loJgP67N629GBdYgbBWfzR2o2H/2OUesHNvBLkv2IrkKSUrNu83g63xVJCbsghoSmcWstEQP
2Zou8KX3PQmrzRB5f8jA2awg8cxJWdrPHCqxzUGoUUfnMJ3a0ebP6XWag7R+uqsSQH/C84ztGIjv
YQjt2DtXk7g9Fd6iNnRIZlhuKy8fS2t7MDVHcdGWI2fsM65J6LjgaGqufXsQtLKBlp1nJ8V0/9hD
s7kM22eZBMICUzWk0DzMZUZz9Oot8I3Kxg+U3phWP8qtQXCczCo3UUqtgnT93o+BsGboCAXFL9+o
0LHkMwIvGI7NYY1IOwsc7fSVnd6H9hFAKT4Hv1lIxKp/g4uFQ+B+DSxzsqMXmdNFepuPWolueObj
eCjE5ROusuU6zVXRfiUXwrXc1GtM08EAfTacEFP2/aQd3twa6iD0dEEXDXXdHDXvenNO+rxuZlIS
zCNKsLqxr6HOo3W4z50dEPElNmVhaH6MLzcRMmksuONw4l+9F95uAajpAXkaLMAerC7IalYzcYKS
Aiin5vxk61V/7pPi+Ri8HrIPVqoCJXTs4MqYFnN60+JKLHfjNMY+2szFL1dfDysyl2xRHsuwuCdZ
2YVSULw0r7c/fyrVVom+yG8+w2eMWGaXNjAA7fpm3iiswKCBJ4uxHv0cuNH1kvQifqMmqOM1kP9C
VbDCF3jYwql3iqiabdLTl5Wka2drgnayRx9DGYbt5txLoSE9NNWQ1iz5tpCEFdZ4vdl/p9nNXYke
grRduVOjg+9/nH9gUGUwUU2ZxBfbG7XXiAsJRRfDMVz0rvQ1SJ7dT4XVMTXAbAO1eulNbMtdC/95
mCe4EuBWL6i+FXpm9Eb7V3H09XdXC0+wgfz/J1Il/zf5kmFZK73AVykp8eg7Fzqw3Rv8Gdl6EmIq
7VyzfVmeqQkOy5DoEYjfSwoRrwEMlBns8Z/mRcGck1MolQ6esf/ubIaxjOMaAlsMojPxv1Sx0yC8
cIHadTT6Rsx6NXIsbj3xWnu7B061CGjB5QMyPvX/1ZDoAU9UTsfiyIIOctn5LFsMkoh4jqoXgX34
L2oXhZnDswStooe/12faxi9JeM2aO54tyh0xCxbRJvGtA4oFDkBCwRpP1ebgqbZ+Wrvjeu1lZbCn
k/Pg2tLxJyo0Q1pgMivZRvNPdSIUBKrhAo6+7X3dxSSU2QizwcLgaYHwyOoeEnS3wD9wUGz/JWZ6
rpC9mT9f8RaU/Qbt6EosB9sTJoMoXQrTFiKoeONC+0Y2G5vl7L/ubzBu2j39i19dWo7wmVJivE+C
V00NJEk+cpUXUWVtctu6sQqkq9lZLlm7mnY/rP9Ll0b6yoa5aFS5dvO/Vw9ynfcufbVp2EySnHkL
FGnFQC+SBivggIJ22Q8LP1koH+rsXmC2sDXX3BFUudyyKnbPSPaL7Zu96Gu0r6XyO2hR/xWWD6lW
gQBHMposqRuKYOykWdamzsJmwy9Nex4y9UJHU8xj+4FMerlAlZNxICeJNYNC8lnQduz8GkQTYF9I
njDVbZ44kskWfuiZsDRTBExLpGpbn7LR09kfEjO9fmkveErgv7vZn5IdmzGM0s9fmFdLIczMBsym
l9mFOGk418b7kOrgDKETRgRl535ejDZ4CqCFl0bR4rKtof0Ym06fqdlU4C5mKyVOk8pwiWWWUxuT
J87onL/tVmTjIgDHTaP/FRaBajrkR2c48hih01V+Q1IbCr8tsyEB3/GcLXM52eiLXax/QIT54dpX
/PvlsT7eqag11hR1Vi68aKnC8DI+IrFdyf66aU6HCwoOesrpMIUyUSqoEeWshuhKcGc5yOoJkoMM
li/D9eEb/R5fuCmtQgztlhlII8pIzk3l+0bJnZ6N2aocT2bs1W6wpiSmiLYojsqrZbGW3Hsg99UZ
Q4krk/cYQk3aKlUG3yStpxbf/PvZd+hSOSJROlMnFlRmdipg8Rpc+37e5BI0UhQ5pKP2Gk6mnyIP
SabbB+4LwvMn+JBKyUCjssGo4+50CiWyraWKjx8Cs9r8nkI+Kfl65gXYrWhd6Q82pcRcyDPftARB
pvXadeTXQg5kFiysm2D/u8zP3t4Vwk8dlaEA8kbbN8RcNwGD4PWV/pDsuSSEtUX8OM2Wr5BpcKtq
umd3P2sVRP284RelFvS/6cLPKw4HUgKOeKofh3j63gEfI5Er4R2EnexPeOtWz63FD0c1Em1eqiCe
6JZU3OmwlkuRMBjLdj6nTPz2STzAl4s6v8Sxtg5piLZmtsYZXiyCpD2VHxqd3LQtX2IUQXYrVmus
0Xnsf83NCDmHdXoG0BjVNA6ALNk64kxu7PeJwIskvjsCjffMxN7E5xgkY3YmPEhnd6H3/V1v8BcB
7vM7Y434m9D7StfHjpTSW7no45I3Ja8TeNKcAbzBREUC4TjWMBx4pdcaHs8M2tUbShlb7xJohN3R
r3KtP1rN5T/5iHGaQe33EyR3S+qgrtKssY4dmGgPE5niSG07pO0LqpSyloXx7m5kkcM6i9gqp1sX
4NpmbA2dN8ZHSzJoz03g0KSXlrIrzKtcKH2iNJR4mvp06zNLasZuUO/Ov2Rc9tge1sdBoc01+u8V
hm0/s4Sr61ZdYyrXr9I81CTSIRXpBdo9W44o11VET8E1M65lzCQr8OtJ/SlFGi8yl5y2UgI6tptp
SMJ5nIu5zBL19gqkEYmJ2inxwc29cw9gS6afhwatGcLCOqv1JWIiyHyvK0Ou2ADvfPeH5DcUMbkD
Z7pED/jmS/EP9Xlo47piGHPS9CjjDiw9OWj3VUdtfhAeOvSYFLgJfMLXyzCy62DCajT/StGgKzQs
WtIHje+8nnBuWm0xLTgU0QhMazoySCHSFgf0WAIjEVUn5lMBzB7ea674x96BpmVTeMUVLAcTxYaa
zbz6TRHZXWhqax4Pmo8SITjtqp/QpbVKFNUUQBKa4w3gdUkWydy4TG0GsaXOTU9ddI9l7C10DrLd
0XD0LuOUJRbZd3sjijuNvSMtwVkRkfdO7R+TibjjjBdFDZtjDex8usbhLCgU2bdeDKOLHqCFWxW1
ums4RyKFarWQe+8mQydyzggTb/Vv3xIzfR/SKwRsXkiTmnZZWLDvmh7pef/PCBdd9dYCWsUyYxTg
5fGHqRvIg5NyJFjkBPL/VItDVBGYv4J8+7G/qnw4kdJEXQ43ZfTskmIck1nud09u/2wO5PC90go1
1DNxHkByEzAcSpqrNkEWQ0vW6/bmyIOzcQJHX9le4BpAYrEtH/QVcs8iHjWzO62kIiMu33XZZWSy
2oJ33m7i/2XL9CwH1BjwSxI2YAmO0mtgmTIVSJLWgv9Ir+aVja9Xwv2xoqI4BcttHAS1gHytD/UX
PlUcd3juWmdZbCwUCnONvXvdjhsROCAu3+DWTG9hFi4L4mBPdEqvzjeftd2zBjI/f0iG0JtDKLn/
6XVFpg9aYSzLxENPTxlz2a8D3bL2b7mFEPwPdX3/f+4Wj1t4YsfrJ3pijN8svEnXHyacTeZwjkVL
ohH1wQ/SnoI/jXqDNifJ//pvr4s/RN1mlGm/gngnPLqgxA1518qYY7WTUF1TkYzvpYPAJNIOOYKy
q/6Uj4+RebHpCGmdQkWreGhZDWxIYg/OHNQUGBFIVlNeyXC7izoSoQzGJpi1G7VP+pR2v7Wvklb3
V5ISHsOTHPV+x8+KOwkj6UMVLEOM8EefMIKdns4tlg0Rm580xGJj00yuxYDWFj1y2r/ZKSVkdL3b
a6lsNN8l+VL8tKJsfSxyvDm0kMwkuWdq1D1PAqAo1vnVIeu5acSFVetfj+wGQCm3S733ILnFBf51
aDzxUclm1Rz2QQN2h/guMBUZBGXMAgzJweqSOh9cWNMIe5Cd/zdDCAVeUWVKpgX8Q1vsA9PXwMyV
KX8kMyGsj5+omvHtJx8Bbw0gKhR3pGECwYM5OdSZOgbMOIJjCrisrAqvH9ppyP+iGaAWnhRoeeRF
DbEbCVXd5UlrnpAUfzZ9kNCNUNwRJrbmmpR/xR8xveHLJijnbhbLT/yGFSqBQ+LNud/CTl3tkgaQ
Rdy132wrd8OHon2z/DAqZ/R+QT4h2AjLqRFzi/MNS9ctgrFpFzE1oFfulb0FaUWC0c+hcHIZErKy
a+JCMAj0fgqhkopK5PslWYacMQgGxn68huGPQ6kp63qBBbp9sbF2bjQDSr0H3BczNM3PYCLx4niZ
DYvgj9f7n22BnKh0e9pG1D2GLeRAPWwPIn/yQlRhj5Y1gm3qAUR4jR+R7f9fLEGv3bW/26usOGWs
twBrBjJy60LE8uYLSwkRarMCmmPX2qA+1ZlM9xggMDKl9Xa5Bcw9Iqa2bAKn4cAyZZtoi5tGv3OX
4QmPayok11mkkPaW//oRH/EJCGWxrd4R5LlHwab6vlRyOmbWD/YHFyowy2755Tysm4rxPU4kesNq
CoLbyvu7xCjUPSekvDTPuvhE01HUYizk2QyaTruUsRnEfPQMNMa5uZhgAnmEsYQ+RW8bJEjf27NK
vdUfxVFcg+Dll0hlSARGANkdHrtBLI5mvSFDjHUF0xdtyP9c0POL/msJvgDymNO6BchMS8qay+b+
IdzXSuF1/uTUZzu5A8FyTCQqjOrU3WoZCNb4muv7dP5uxq4aiaYd/TS8ENO4fhHcVpoGm3LRxi51
c2wDC4dxzK8xBI7/6M+NbpKVxAkzJGx/SIoMeFu7d136hgMQvjyQiKXuMGyTMBUofAl3cKegNKzT
qVegm0vAcN1QIB495O2WHDKJGEUF9PFfV0RaazQ9uA073hzXTV4X/rHLQEB0MeSWtEY4kYoVEl5o
UoSI13/V4uXZt6Q6hHxjPhgNRyIo0vIhnFJBzPKponjbD54detFeozfaXnfdEWPalklom1bNqHP3
hWLQKJ4o/wURyzRDxkiWGvEDv3RUYOsG3UElu0YMaV/tNJG5uKfAa9vGSxp90A7nqQjt2TjokOiO
sIY+LUJnZSkeCV80iCXPbajnJsR+nQyvJerLZdKLynsG7b3upPuPthBbKSHH2+OZG9J6PBZdrnhB
biDbmcOM2yuqsLsymTDcm/0fcBW9xAVZczTlxzD5Qt14SHwwsdbqt/q1MEOl27bynhBFBOS+6S9+
JnJIhjsLeH6qKQzESrRqQhzHnA1phB2cJuH8M7ynYVmOTJd/kK/BJh2qDzfJLavIdwd+QUfdAD0h
A06DUvqfmGWVln7R/5kgqKaMIoxWxQXfkzuoZL4Z3nApcUlMBscf2UqmssqNE5titudo+toFU9R4
zI36H75JSTB65HcZ9b75rwoGVQGdFhVTLzZRTouaBwrrr5fMpce7xeyZNKMN8X7rjJ7NydstKmDX
NZImidOjKMjyjmu1LSedZuKPiAlJhicxwak18HAS0HECQnZK4mbcWjM2PXRPe45lZfGSDtxD+knf
o9ZNUdWbo6572nFkZbVs1vA+SFgUMcuQ8AA18D1fx+ujoRZby+imAV6Aman9fiZA4vyzdUhRvxFj
nVYvDyllu4UbLeF9ySva0/Z1399h4q1Sr9G9wO4ira9KZArxA73JyI9kTdm1iMg4/ZcO1OQyDfJy
Tkdf2BDHMiIbTTSuJ+Er170BE60PZRKyfxJ7iC9uJ1uUgl88K8r0ndOLdjdgUT/42zb2wfSqiR81
rLKxxAgaXGDkphcPelSFVOUXZIDttZegZve7i4SAGybg9Ll6wcYsoeCRZqgQMvMX+OWeDpiNuuLg
FcSOtCg9Kfop2C8kvBjANwQ6brgbqIwQiBplpWOJXkRTjoiR+RN1E+lDfzfbURygXOG0YWkpbEsE
hu7kuLBHKBsqdoQ+sgP4c48+GeaxF+NjfZDB6InuGghWGH7OCEwAvFRa0REsccEmOAhxuxLbHvs4
KUBuNUja0uhVz/GHOFvMnZLIqgRAVfXmseFZSejOgcyKAQcpoydZQpiwhfIVYPF6JmUDfeiriDA/
CKLq65xqgdZMyh2WKEf6U9BPJ408HKo8JJs0fC6VfFCzUoZMey0kRX2Z8c0Lrs4nELWraKEeUdpv
P28SYw1JHxIXNoiGiyl7IftkH/0LbXCqsy3VoB4NGc5qRGssH43rLXbXN78GW3nd65zj1KQv1/5i
h4GIS18lG+FZYRDt8FTzfejdoev/vGQTaG0JFTn/yJpwLgGr+yKhGXVmZ+djDKSMW0V0C3hS/LTE
z2+/fozJxBpK3b2J5Iyf+UIm+7LBc/TyAgaC46K2kdkmb8re/EkhZ/n+jdNB9k+sJJGBY8d9SnYn
7D0bz3WBlaEfXdPeF7dlyn2Ns74v7gFwCTBpAlT3O1y0ZIE+MI2pOnEuuI6vgrn5pXn3VMDZW4QP
ikyUeqKoQINlMYDW9QgsSup9oTmuXIiDOgOyEyyZZZ0eUy+cdCbyOlxaqgeH9A+rv8bYp1CjZfHq
34AcA2yK01pYid1Su1njHLeYNhwdwUvRX996rFFZ6jymfPtELPPWiPvfUYcJbLX887oi4Wjihb1a
UhE+kEGMQH60GUMrPUYiZUM+NXvYD7xp8dsNzJ1hQntTq3aCPB9BGOsApJl8KQGDRV1qFPMgztF+
2j7RtA/lvzNA+G5y3pIFn37oWar+sGaoBOqAxwEalSGNfW2Ygpbt5pD6rS0WwDxj/1FmImPGYl4t
9uz5b++mgvq/KtXNkyOnHtehjfLSB/NvMUzSrBAlFCNdMbIBGYNu48SvlwcAy53KxeC7egK0xskS
Oh7vlWfgIBxfEcrk7v7RlIu6lLhORUt/FJ+6tFpVn9CozYdcgl0PjtJhvJChtWPoi09hK9pX8oEp
viZJh+0FJ3leDLZAnL+d2xi0cWFr0qVK7CmVxumSaWek9Qt2fguoJfyCc1cmYHe5ADaSKPnLNzir
9xWbLqZc7Iy2uDV6oIHDCf9xKjT01gG8IB7UexylvDQvihKdcvs0L6wMU3eOqT3hTW44cjippwm+
RupiyZ9CDEUjrHpP95BOFw0KbPRCyi3akKSGcTyga29NeqeBCuAQ96hoMZ29QBkhe5ZWWNpqQ8rt
hJ/+YaF8eG5jlA0pwfYJ20xo2SIMxaSdRPZPn3yF2z2WzvYU1ZGqRQgdnIDNv+mU1RUyrNU78RwQ
yPZDcUCJ2l6MQdVqF8i/PjOA37kl2USklnMS8d9NzKygPEJce3WKV03WBAKx5qwYdcPoWRukJFqN
L6m4o68xGCUiHJP2rTbr8PPQZm+Q0QGJfKVoYRf1v+q8w5BVxs7O7FEdHMaywx0asYkfVXoFw89k
yrcFrI7z4eWWGO0/zvTIc+AFS9UB/Y0ZtIbgCXPIogdWT15efLj5RC5x+k7fHPUqMGiuxGbYXofK
F4c1wXm2dtb2sAf3LtFrzaymuT8AeMAp6v/c2fWFX/0UJk4pWJcoTTmCgcVQLy1nCbJVDEIs5OzS
A74yYLY9S4S5VdHMf0gUnCkFMQRVoUi+KKx2BPRTFUqt6WY8h5pZLIJrtsf8UEDWGjh7sQBmqVIh
8q3gre+FmF4BB0P+wWVahhlxsw+vMcEBbLilMF9txLNCbXayUZAkKjXPHSgdQJ9/p2PaL9oIQJWW
CxdXi2uO0+j9gSOx2GjAc04+jNRDZmKLjWnYKR0/D93KFi2y66jmmswsT5mBCCV76QhAXY/hmdky
FAVDhd50q5y9sVEQbNNWB3y5G6ZdoNsqLT2sMPbP8+H1Skyjh+RZvXcX0OpBCVdG5I04iu2qAj0a
F4Iy/nvovhKRCn8W30dbp6ZsTi7f7muzFidaSTIGRr56YzQtehrnbWN/fWFoEHQn+CQN3vuU9tWF
EtBlE9DYNpoaIytco7n02wpIaxkNrNpQ+Hs9ua+a3hnpxV0kWp/UAC2UhgEPE6IlqEOfTPNdtimI
edXqcQcIIrmLPNVIJhCxn5hCvKoMik+yl66m52vCpLPRKdattNz9dJdZj54LWpotvWLh5Jwsh5ML
rqfRRiua6oDnNyAGfRCVqiMAseY6+28lGOT5i2B3SubKJNm+suO7RalrjkjH635CfJ6AONk4NiXe
OrHLZpIjKUJZExKOkaLVOTK7jZNNWBxcLUbfEyDFcShiUJj1ChSG7BTYLSkARnpEdiCHfCnjF5c6
jyy3pnACTvLP+JBruMW8E1udrmu4LOrNNletx8PEOnMMgc1LTHcmW4Yh4pln5k0UwYm3eZhEPc1G
4+PJ3OOveNt3daft3O/joLxLqiExkxWhLuSsuzIs4pk+6u8KgV4IFXETmTUpGZdbZayuSS6yQ1ig
sPAjrFFF1FiyTx2vmNw0HHojplit9wRTFgoLUlPFYd0y0anExfyAE37oS2P181sEpmXVxgzvlgEg
afVZsDzUO+fgie9PH6syvgu96ID/yLDxqPth8dPlDAbCQ7gsN5sJI6N+opc7cKsxdOK0YF3DqpJa
hvZiKsSXLM8Yn9hZHITUbmbBv5+/bcWuqWyKlc/jExl9DuVe1z3Ao1pgClBYoXR6SqfgM8pR7D9i
7N5xZnZ93LMffIdUcOq2Ge4Ip7ewVCmX4QalJsAgPa2j/VZep/fCm+1mLocShkCpFX13aYwVlYG0
lV5gRStzLaNHnnHQKT9T3ukwFhzY4Y1zJQI3VwKLrKYYLozWuLNTdjYaU/gKPnYxAI21kUcOGUl5
yOlyQ6dRPrulmmhrg3Kfnzbu1ermpgWuSnF3qgTxYuQB184ABNmR9+SOd7XuN+Vbh1CPrjNP4z/c
tR7tXw5vqK/oTYbyJoSoGNxSFQWJkHsBH+be55z6xfX+YNB9wZLtQvp3JvdPhweGwOawreg9hDwm
PA8FBeletoxJft9f6RtZZ1CLIBqShUiehJUomvHjtIWPf55Hwldu/chBRH1ZfnQEA8mvRQvNs8Cm
j8cbABGndUyRA30BA07nbMCUJfGAdHyfBDDzKOpLIsLuoZ0e+CvXbejv41PcqwGZGxl+zwiejfdl
8O3lF8MUKjGceZN+G9aSoLVGX0jG4W35lms1E6D4LEkLDzRDjCro6ZY6msvm96uU8WokXHOfvp7T
3ShpeIvT/mR5jn3yIj259EE4IA6BFE1FnuIbKkUq/c7X9GxaBv3byEnAuJw+nWzDYPMZUhcHnq4g
RChvyzDs2k6irhRfi67L0t4ZAgQbIsgwQxheU9TC1pY6YPJewUkbT/axyXIalb2vzwAQZmYW9fVY
GFgzu6pbwsLsuZBUYq/usJfPdKrEdadekVWAXaZTVGsSbavR2mTfMSLZpbt/4DXgRwl1BuzH1C0Y
pzel+xGjmMyUA3Zin7KeTWkXAaTAmiWpSFsWR+xv2gGIJdYLT5mtjhlQuFziGbjYGMJbQbJwwEEZ
WHYnHPme4PwbYVKC6pLh5pvVnbqYnC1uLYD4XtAoCPWC+ZtD977eXwaS84A4rBD+Z7G7mjomQOPN
u3zmpyunRAxqRIMSOkzNRdRKV4s7APIRWjocqRiGyEofwCCyIMaTqNSqUcp0rRNZPBnWov0CY4v2
8JXymFkcwcxaKl0mXDkmT0eRfPqX9+/7Eir0lkkvcyzNAVtWpDvWgM73mBS20TjBLnzvNEDaGJIg
46FFog2NaAUP8BeIlrbTPCS/N/19Gn9FLmqJpMuv/tQVhakjjze8R7SkCH+bQg/PjIaH5wVUEJJN
7mUMJB0s0ysSorusVDDz0OHf05vtJKMwFIDSzLcUnc/Xq+ro+Ufzi93weywREIuD6b/Lf8gu2sqk
o/iBJ/seXc52ud1kRfVNtKn2egob9cI46A1Sb34qfrHuZnX9SKx3g+jWrTFf+KNGWsDrnVYlK+2w
GveyhYTnvohq1uTyiA1l9CEPO7LPhxN3SYcEZM0+oETzldtLUbmvTm0wzKi+wloYRUqXGwI6xiFL
emQQKTvd8Epj9IXygb9e2RF57cBTgAy9gSZmx+zUaHz8UzsZYrUFkYTlORj0jsayNVwbHePiU6FM
qc0On55o6gcswwYnomyvB1ybe9aAEuWettBb0fJIwSRAwkjHqGCT0Pjp8hM5apEaCQZh3Qq+VIP9
6NGYl5zDFGDLk49go+oThZYMTpes0ogQClPYHt0aq0FyHeNzWByLh7e/FhX7DYOQjARv9dhCkDX2
8aurqvWPWqPF7da2HkxsvYl4phHOwK0HjKDHs35AlUHX9bp9Moa+6x7xU98KcX3wbRnuXAF7qedJ
QqVCDsq3A7RsI6I8oX5aUznLR5SFlOZ+AjUiDBjVpiGj4eXdXLJntWg5X0jjTZO70G54lzwczJvZ
A35uUsP3m0UrsbvV7kDlq5F4mC+vVPnlmjSPNc3XNaD45uyc9c397P+QL14p+DsTRD6i2FysQJNg
Ep14FMWfO2gw9KSM/zex68yIFe/bK3ZdgTeuF3gTg4j8ogcxdSkZKrAgSXwMApWr13iC9Gh8C5Bv
YFWkkGlUm8YV5o01GNVfjIcpIJ+e0TpasnycwNPF7tGqFrzYszLHJQpLB379roGS9eAcYiU9Sw+j
pkKNHhXo8GblRpV9y14t7wjbqnAXdlxvzs6nx2fX42p6pXQGHY6BfEdpT+Bx4/Jz9goJm9hAVExI
j0N0uP65iMwfq/WCXeoXvA21p/3UwYDX3elFKDjfXB1ReNTVMnOhGxwu5z5mtIHHtmF5P4DWHgrV
Yx/5hV2eqe9tibgplmgsCT1vbauLJyP+Hoz8Ut/oSs2IVYeW21VLyMtJvjIujRvGotjhFp2V1kMI
A+/v0eBJjSDQVMqgLf+YjQKmVAfzs4z/oxYwWLqqkdKCQlO2zGuc+qbABnNBIflYahwt73sv8R+g
TulW4HE0NqUwbnUcXCDG+Y5dSOryXljH9uHm07BmARRu6Zl1cB2jE3pHmscZrj6mKQt9rcAIE+SE
6jkc4DEqwXzG+k9qCp2Pwtquv09qdjDdSR60LP5l+Rom07wJRSp5NaabcIO3D0t53n97PeAmfuLk
itmQf6qS3IY/PWAFIwl6QMB46E9s2JyMcAqs6EdbNjzw0XoKFGfSvg2+RDJ2K7ryEqQ/c5FC3n0B
R8/YweieriBAxUVQ6m3scFY7NXsU9Za/3t8W94KV9oBGkEIKhn0N0FQHqR1nmx7SqwJ0WfCfq4E3
nrXjBkH+7mYZQ1PmhAxfnIIsKbFDSrK3KnjputSUAlMHJTvyBY9rnaKaruzOvYngVEFMaunE3Eh8
b0koWsjMKC6majTPSKfpYzM1bMPSZrKSI4+n4/Di1MmdgXcYMoLs5RHQ5M1xDLNWxRnXs1bq04Y2
7iQv9r7xg0xadRCgFJeNsnMjH76e6VSbjt4qYvtAdanpKjRiJGgtBONhKMog/XBtfdKztYFiHr7f
f1K+Dd31E61huWS13IDLBWP/eC7msyFeQldnsC/gSTR3EsMrvAnqf1Vz6Lcy0qI/0FQFQDe0aWRw
+3V2wk8OxHbqlaxkWDP3+udNlNckfZBUHCDS9TIDakQwQDPCDfv65Lb1Xhyx3F1WXvbWnpmZsu3s
y8V2Bc43bJxXXOySgSNapcxOPFvzWhMDFj0HP/+gNe8HMlf0mVYE2K7666nX059lFkMtwJO9sLHU
y/AfPLCFur5Au3fphTV68q1g58OP1xbMN5LVhGUefCaAiKotFGXtNBZQ9DSrXhaqm3fy4YVAcFuO
l2aXAD2o5xGfSG+wbPuNo08CQsNEFvq+a6bg+aVJXsOS2x+HBJaPnk6OjhmesYhDg1boO42qgBgG
KiTYe9ExHQ/o0InLxhz9psyGB/5vZDWQfO3/9oIYXkF/1qUmZZ2g4BEuomHVx2Y8NXh41uoWWlLm
JOYeh9zjQhL0j84EGDg8wd5p3i1Kq8C804+BCJPO3PVeNRzWeEP+ek3WnNiCaosoAXApSqa2MkvE
EBlSjtdz4JDsxugWTRHjBOIKGzBq4HsS32wilSHhDx37HMyUhMZ7IQiXm53MrdbxfOntHP2Dp7X8
VZx3XKBaOEm8dXF1t1jn9SuMvO1m5Sa5LBhGEXfq6VNU66t/dzLpJQJGcz2RHxGGCczpL7lwsV6B
qcQe5Tg4EqF9PNTLoMSfSX7lbXJjOfxEm+5aAsIHlKL/7qavmi+iYQQ2PLlRqRMstDdRne4e6tqF
xk1n+x6PQxVO/D9+JJfFK8mETWUxJZs6WMHI/bMItUJcpIGkkpGkCkq7WXTk0BUuso/E7JbHhNUs
5FeEB8f1SGlOIm3yGFv5wIQKQIaZOzt6/euBhZ9lI4fPK4lO/r5PG+z6Fr0cXhkjy5f3MIqjdj/k
wh9rXgVi2fSjfiykgJLxHOboCY4/yBOXV0p+0lm/LgxSWHlDWMmzu6KWv4pIld3Vfb4PlotYc2g+
8gbH1eJjq4vH66lUBk6Y3wkQJCcOjeW6s4Kj3hPYs3hSuOJeho7Xb2N7vzZvBsHk5qnEtz95deG/
Bs+Cm4fvg/Nz5BgLLdlO5xJf6nLHnLaZH4ZKpgWGV2rK7Kobbi6mXh7LHUYR2l/2HIt7ehYS0bss
UaxD4xuBz+kb17iBX+Kz1aB91okbalvMIc1EFVytInfkH7p3HAF+5GmCh2+iYQwLXj4cgy9Wi/Uz
poeYLCuSCPlBNL9oPtaZtFUiKramLvbAx2TZTeieseAYmCdvTUVnCVPAAUZgohtljlvEUsy1kmbu
jh5JO4ayBSmw3ZayGhtV7slbmxsm0E7PS6KpRn0JyWGahBVBizE9ZXWUicrMleKcirdNKDNJhQhS
dXtg7YS7Pt6mfIV2eD6OrXTlwfXq8Kur4qvN8JsMBqiDjW1Bma98tuYe+dMY2Ske4kpf3hl1IffN
dGRmRECFSJ6nLT1Yh7fyNIwuP4BNLnfd0w/b7oQYi9FP2ZBOiXpnUqPSL2hknC4fIj/q5v/S/jTW
FQg01E0894qvnMAtbYaB/7+mhkaNtSTs1Au8bO0GGeEFheDGW0PftG8dDQVPpCic8WZ4Zryvby9b
5gfTM3zp2+PxPdcxR5jw5dIv9O043f5pzejq2nJ8YU6iEo9qPBGAIVuZIKJfLDA9NW9uk/WhBtuV
+f/95dzcj8BN2Ujh5axH7pmw9ik+jE9PzM3fPbiEjUAo0071ufk9kRJacEei4ivyLhZWZYtvM9Dw
mgUYY++vN9CDlh++5UsobeMqEtV71knHVRS/ISzQRZGdUMfdyD0uSLIVKjbXcDIQbPaBoL5Rxw2I
l8+dU97jCuMwbPHG/u7kOP3VCgrIUkx2kdpG/etwT5a8TjG17g4DnvUC6vBB/ZUtpNuAtJ0Hdgwe
kVzDJ9uqS/iqzjhJK1zaXu+0+jAy7GSNTW5wf9X6COuGACxzY7AqCe8StmbvT/+/Jo7mp1I6EirO
xQZabCUP4dAKercuDLcmhHDD9NgwvjbAUgCcbgAwF3XnNlIIpNketMCBtOZndpCuiWu+RtLqJJ7m
IopBSRlMYpd7EfQaKefgQd18E1m1gNhO1wH6c3EZ3LOe6wyg3JGqFNOS+iqkxBn1CWRdFpndnAiN
FEh2Jfl1lUbYTzTcy0eh+5TITlL04PA18b4WtwPy15j2UQp/oI7dGqZ8CeMrqSaxFdB4GkIgF0OX
Rs82T5gtqUpkqOezFQlgXQRufInV2B8esH0gCfHSKkGBNaIGk4ch0zOAkBq6Oxw09KaXB7YsF+FX
HZ0riXLaIoSioJl0u55yItXtqqpMY0D2RJzJ2ALMJ6u4NDHfju8CB6ZKKUt9hzIopNwnmOFo/ul/
HH7GYB4axr0EOrg+WO0YjaeFsPsUfYTwD/UF8DBDUGfv1HacTVLHsHsQRGZtcwtqo0ksidfRuwwS
3EkyxlouQNCxR9oBL5a/X/BaDjiXqX+JDvY78Klr6qYDZDrogVvBM41h3xvfVDvmdsmJggXwEi8Y
GWDbX3cCdxtJC+Suy3lf/+bJVCXCwkV3WVRPD6dEdyGM4VVGF5mwTbJ1+fTJJHFISoFDXtXIHtJS
NZQ2veXt8Ip+uhgfXhLibbbcuuRymIhE1UHFxk7OvUBl0dP+GJ1g4KWMEdxPS7XUjFJnbnBEDCT2
pF2aPk8q0uzkgeA756Tg2P4SSWb309hAHzNr1jhKRfXZn5Z23qNFEWAr89aV40b33eG9ZgD0CINB
kfIEPAwE8nnLCTPOXfjPLFnwGCRFO2/b3UHv7wnh+HjnlikukxXrdBYo8u2y4IVdvL3d6X3y7TIL
k543ZqvYCRyiRuEiA7r5lAl5sS2U+ElRMV5Lpi9FiyrvYxqM13h16MlFJKp/6Lvmt1u6gfAGprQR
mgjBfwG6WerBCyqnc3ezLWbGziOV/9gFhPzd+cC11pMYOPluZ5y2Iawg0ACdeklSeX7qGR/7eEPd
aSKVSNOXPepuVxPz3HFgerHkWx6r176Swcdfstaagt1sVU5kbSIJ5sccusAkMITZK9t7r6aP3kFX
zyQqQE8dgabkSiHi79G8ua/+H2scEI5KAGhuNgVksRTifkzlNdILufngdO8Ges6qPOB3yYJHjmXu
dGzi4xlWXqTtJC454p5I9PoM/4CkZgrfpM/PXUNd1TZaH26HH6fb+3Q7pmYoaS5cbGk7HZQwM7w3
/8p170xjeWNUQG6ml4RVoq2lFGbUdUZJBGOJp3WWfL3wkWTaB1CBL+kTGaHtR8D7KV99HsYmyrcJ
MmM7K88/BfSgCI3LOk2WkhMZJgcjoK2iyWFcHfa+gdoAWLTMWfxwmRFHtRCXmSEtQRU4kz3PXXji
nqqU6l8k/OmbA2TH3qIVhjup+DR69t8QpE6Hp+LVyHQGOpj03yDcz5JaxSWK5oAI1edQpjAtH1Vl
FFAI/g9MIoq/p402qU7NNfWHZu6BqVkNJ406w9VxBxCs3SC4qFMsmOx80kgxf/FekMLpLSFRSBYE
PNdbvYFnubjFfkkGdK2Wtrwd8H26hOxjgTC7eMfm7sWbhqfZtCN0nTzI+iclOfHJEqlB7Ej+LPCW
L1zTYSQ3prbo/br6w+elGFNvdwkMy73DbXQEIS/48d3UryJtq/LEJOvaoXOSShCixvstPXoLe/Kf
AK0BAvQl1eOD41ekskYaOPb1aYEk1vZPzIVdjcxMksfQ6FqSrrKB6EmYeaWoH9HlWMkvgrd82LEm
cMkW58KTYbfGOkRqZokiiZIz+gJ/kIoRsFvLQICE6bMwRf2QGEs0dN40sVeqGuQOo3Od8gc6halK
cx7DWNi/2POnNHytaSK7xq9vgCEETF7cahMWZ++M4w+xJqm2MKqWWu9Xv+/pg4S78iQ1R6kMfZ1R
ce9hfiiQAhjHwKlqVBU1pr0pSWDPNDv040DFT2CgknDhBvK4qvGnC34EHTiiDHLW1qyJVykDzF7g
78H6r4I1bcggCTtET4Sz5kKHTWg0eebxvx3gCjLhLa4zzKmfGkFCbXz5xLbUsei429CWUihjB98q
+NgZB3DjUKZwstGkje2ZELv0Ev2LNsv1tZGQeWeQNMXUyfUbMMQHT1L+YaJuszRfmA1dH4FicDjt
XsNoWBzR2C+0gvy5eM04ILDwExWi9Tq9Wlet+RBpDzHcZ4rKOWPBee4ZvuZBcyXZqqcNVaaHtiUk
ZF8pBLoXggPS3dVTN7UJN5A9nK7jvWRmCzqbuPx9ABetCQm1wilFKW7kBwZrduxHciLvqGcqsyEs
u30lYJCe+O//SQzJ3kRMjfMOcWknQUP8gV/D0e8U2rcgb04Ke77YzJdQxmoAzB5/qDjiwEIuJgCX
0a74vlY10QUwVPaeHfPWvdoKWDsQ/E0o7PDPRKQSEWG3YYEA2mv8jl3+sYXpup+yeAHLRYFxvvve
EW2m9GILJ7wU1mh6plF+Elbz+A/ZwwQuKSDXrOuEEBrls68xNj8f/tp7AgurmEVNQ7NPRoYi1hm5
2Ye7ju9KKEtIZQVlQq2RQQfAdvxU6d9fgCzjkhXOvBjJaHwBEcATblAX+/3lnUKymhU7jl8A2lZz
zf527cDGRkWr/bbx42v6/QUscPbOkuvTDAERMAzQIjMAnlhS4o2L8nNYH/4IR80dsK/DPzv+aU8u
t9NBQdhTRDM64vsiYjaLfx7MZLVKL4zTu3Wo0vfC/nI+VyvAd7GrVFBx0jaPXAfNjPkZbcb3DdSQ
A4MeXTJkc7cOol+eyuYKXL7kBAabaM7ijseZ963Px5d4q4eugOAYEH2073//i0unZy8QQph2sksX
G1nApH3JmbdXcd5vchCTKhvuDJMKoVmMxXSWE3Jv1jeJoIdaOCuUbpjmX5M7McT9L2JAuq8EaNiM
8qIXZ45/OnC2ZtGSanaxLfL0VStDwAHqH1UjnTSeRTZldrasA1291u7q2/fv2gWyDT7GZyypJi4P
1Xck9yZ2hZ++po5/RukWVYEme54Wky4XaaT7cJW/9WnQT15DSK+gVZZGGyd1kj5yGH7IaRvbycGl
Hb7zaCDcGkiUsaQ6ACMPmvxaJbf2GKY/rldSfv4+4PApz2D3h8CE1moauKRsyYwGQqOyBpKPPwxa
Zk1LeeD5T8fXa2fE27UwNeQcbYm+hmN9uAlRgFW0WndsadjCt8kqIQCK9cIK4hcytyfNgKrwb7ZE
nL7uetp+q6RnqG7pph8AyteJNAiu3ZOiA1ERKk9hVaRN/Fcf+QWU7nS+SHmnVaclq7YWPlUDdFbM
2ho/yhoKG/3EgNYTLq/NjqQSZoUkAemBLOyZ+s1FdOabfgfF1/8fYspM/2LgyQpEeicYgzGBfBcA
wQElaTbay8uYu3Ag+tDC88sxGUyiJgIG1bbSZpmUNgw4w9fuKVJmJXIqpzrb1OR4KCNLWEN+qWvc
Kxw4z+VVrAN0l71TuI1OT8sh/GGL9NAxzU2xqhB8d3O7EeCDGgtlV96Ye/cS2mnehAL0vZgqDyaJ
1uxrNhOnbqb3sUb7el9q8NCeH1Z1aCzRu/Ho0HteprJbbi8HaFIUqSsXVsgdaeCj+ClefCZZezYS
SkRBwoa4L5TwjUp28lzkga6nQqgP8mtc9u7/9S8l0lc23nxCstTvq57Bw/tSBhiIfpL275E/Y5ir
kptBKGH0vwIXiXKpvZ2UTKEn4xZ07j6BpH0rVyOzEZ4PYmGQjvIDuMih4yGUWtSRNLa25GHGmtSX
+3qPDwiM8hBdj7+RlUq0alPwPz4k649rtmjYusXc6CO5/K0wU/R3FKyI3sTBfb/2TrMJxw0ZcqzL
OGcv/I+DcYtvDndMiyVUsatwiTP/OM2o+meeNIG5OVIClB+wv9Ptx4f2Kt7cwDzbk6fOdgF1w768
i+Pj8mzx2Hu7h9WdwbQ45PhfUvxriyzvwrInwBdLBRCAE/n3ehVk93bzvz9pZk/ncVuKg3tCB5i2
BSqRGEYDmF7h/VTroMl+WJoToIm+OPVpVYaOd9vGAiZ27jPesY5Q5zet68xk7otQzKOoKyzoI4pD
yoiafNYF1bdzJxf24dcwp61CeqHGgg7CWHH0bYoE5gaRWFIHwQZs7j11fQvs/acNHelC3/Sc3dFV
6WOrAC4zoQrRtUNbGcqOmZWZ/lAaYWO7CK1Yu4rHb4RG2L/a3oW8qnysjA6XNU/HlY/f71WsTA3d
034R53Gtqmhwk8RSQbKLpo4ocqnez3SWDTXPhW/EQRJUybp/ZEvOmWjvLJRCH/K+mAheJI6Eu4Ep
9v48wfmrGOPGJa0g4p78U/YR0mIIi8Xtyq1+kGyVGwctcIuPTrMNV0RnoUE7/gIjMm9/flqHbHzI
ADAVcbcFq6hQDO9q/AGnDwxmczCU22n1qk7CPe3VfNO0Xr/4Iqk6WFQVNKT3BeJNPx2EC2md1d5r
hG9Q4Ftbz2JPa7TC/THpzI/Kd/tudLD39AIfk75iXD9cJyZcF07g92QZhrm1hy+RCYqmbdl2f85A
5KR0U5NtrBA6S0n1e3oSxYBkz1WRnvOMm4/ZUW75NbhVSBntTwYqUtQdfzk5eTMBexeWocKzI5wV
CYhMefRVJREUvoBJUVrepgXnaueM78i2iC7SHhwaEZAZ4Bh7xgPF4q8eBDAAHYfsIm6USGm0JwDP
4nvdiOqHPOOoniJMSZqOMH2Hk5BrnZ3/TgVl0RdaNVSM0I8YC8DQqUL2dUM3SIAC1f8I4KKXLCM2
i5Ebd5+ZqPHb6cQNlrFutd9EhX5uFSXQgqcVXaYLByGqpPpVSYIky54YkERr72/OUl16gK2Kiy9n
W4KTNbYwSzlkxZn41pNsb219pc5VnOCuBp1cG8Nxb7WF/vzFn+SVIGg7QSSkcj+DrIAw7I/PgpCv
EKrvJTk4ZwrGB5vHgl6Gcg4Z0Vn07sO35OjiieUxxYLxFpNRsa2QxK7Qo8RomrUHr65RlVGo6ZuG
Lw3b3hwifYa7PZr8iZqZhsV/WOZSbF9mVgwXZFYoWri7lNLyRkprH5XZqtuRaNZyjrLtXhOEsUFW
9fdxu5LbRrPy2EIYis0xw8/SRPfrk6rMBQ2hTbzFiWvQ8bRGPE3nKw9gCLsFIfQXtiDNoRG9zxiQ
ksTkDqdTXXxrEvUmw9L7NCMfwhbFVeXK1D4ckL+/FOqnQ9xYj6C4CyIv9iqw72Sn5Ky3iVz5aeBH
5nkcvQIas8G/5ZuJh0xX9LjtYga2OTNC5RxaJF0VPOX2SfdlYg4oOZQq1f7nQx5HTBQ0/VvhEyXk
pY9trXBH4u18ivD2LupT/ifooEjgc/cZnpwYq82OYt2ktG9P11E0084iEjiPNFTVANNDM4F49ewM
M+7L3j8H2SG/MSFOSQKwv1mHXXWYNef+bT6gFr/qIMJe2aMNOlWBEACuE6crbRTcKBWeMb20jDSB
KPvuO1qdBTYgT3oQKg/2O39+8S7bGfBnZqdSzkkxyhNg31s9Jyd0E/qPv8wITAVO5eKVvADTmofi
oTqn1+bt99gVS2s8pfW67koKxFAowxT7Ws6gpjLD3yjEgtJcCt5C18V7p8Nl+MKd1oHRdqFuTnhT
9sn6ULjqU3G1PiLOwAubKbvlYsOePbAvndScUKZVbt7IS7bQ6Wu+Xy+6n5MHioNsHA5ZZT79x0eH
fhtQGzH778gLOmKis+n7zIUZqxisSEu9HDIxAKvimgqZFhr7CqmlzwCIp3f8j43f8HnSez7Me8+s
JzbDIaeZn0IflWOkXwt56SAPSTJWclgtk49Ioh3fxBu0espnkAtuWcN4V3JcuWt8B4BLBU7y4khJ
lQ5y5x70my36cP7nJIw6JAVeNyEkoPpuutc86T5Fg/gK2nSX9QiXVOl+ASx3ACewjVifRIpXZohE
tkxYrTN8qfNM4Nrx0GovRkPvZKA+FAMCZJ7MyZpglUIuWIRuY5gkityQiH7ttNkqe9mtepRxguOX
ail8CnPgSOzCAIfwB6lXHWlxIirmDqyFdDpB9U48/hlhcU/nNi+skQ7u7gnM5jQ1SUl+Uu1np7UG
AtJQpBs9sRDGa9N5tuuRzdjH+GAr5d7BIsd5jjc3HRnyS9Uqxi/6+zQRuL+xNABdxcFxRcykRwAl
eqS3Ok6TlgGJC9vgZKDDtU3Y2dYwE5B1yXhv7kyFmW0NUvUm/ToZZUW6RJy3JS2z7gxQLSRCC0Qw
JmLfPfqBZBb6ky3i82sn6KyXk17n/Q1GxJBwwrzueoDMKppTWhO2UTl084jsf7fXqwsG5TzLmbMb
g8uNTwkRJpzuGKLMBr5n2HVxOIGmiAvl2WtG1n3ZUKo4bf5L7GMT++/xI6y0xtmUgUEC7iFISlyO
/+Puwmrc+yvHlPzJZfvNyINeMqlaTqKNjj03RZ686sPfvM5n1E4Fs2wVF072EiLJ77qsnKRzQBV3
KiVOQDXwSwIJUKjqk54K4zFmz7yYsGagkXMazgv+pZvLdI0F/URhZ1QOD9CEDV07X3zx6mNs73aD
1jCZ/ily69Akt77FfWemu/GR8WV4Z2OVUbT6zZi6rwTWyahz/AcvIwAUJ0rPuBVxMeQMYEGrVBtT
HJNu2DSx5W2B8RHcuPiOT20XIgIUAjRVHaa19exDhwAyYrzlHkad7OdZKPgQuLOD8M+jlX2zp3wR
I3qjeHFlyj3aM+upg/rxJH+yGlOnpMSTAX56sPYKk/alh1kIlHxCSJ7gyiPlh4Lk+jmdDnrl4k+T
doth893pIrzNJcEAWB/2c/xQcLkEe6SFhIy4arX8YBXctwqEzC4gUNYS5rhegIcUcVEfafkFPkQF
29WWBfFuYlsxDKNGJJ8nmULub/raIonTlfuxAyBVDp8+4ZbaQakUiCIY2lhtVI/RutTEZMiDQYyJ
7TaDBeudfX5cWmHHoqcRvfAfJS2KRz+TIiciOmNjtQO+0CQDkUNtA90AehClfzBZzJTS6OFXIFyx
470Vu2VYgbTBLj5EstUPmQ5XOL0Wgou/8Lxs+aScfRCFwsU//AyZGfIkSYWoO6/oq9tlo2FT6NBO
sVRgFQ0ujiDM5g5UUby5Or84d+cZrrI6KcORwv/h/uy4NJUJwOxmnyQzInYfjf+TY3JVqkUnDeje
RR+T9PamCxStP1yOMjEUz+ByUHi4WRjoAD54yaYqpqviIvp/wYZj9QUH4qXOGvGqyQutMJh6Arcw
jSeYU20KjBml4dkWxBPTFUrkrkNBrAoUy2XGBamM+kbqxfR9x8WITq6bhA/PP2dNyfzOi/d0V7r+
+vAewGwuLLpNSzqp/QrrKn00t/TY40OsGGs4Vg0pzYmieT+iG67yXxFDlK3hdHV17+PwHGtGcot/
yI2ybB8amA306RzXvDN3bXFIjVJhyepkL8XSfsrUIa/un8UWT08SkI7ZOUjsG0mEHvuaL/k+pyeE
hRKybHhh6fFZ3+DB2Tn4qtOVJ8On/y9H7s6ACE+hcKUnY+MpS0SxKq7f2orenR8O99yo9xTd1qN7
Q5rSJNsmytEnSwWBSu3JIPt0CWHMaiJelfcOSYgyAksr0RmFGi7uFtjEcKSqyU+aqKvsADqbPR75
BHMV8uH+sto4SbEigstGj28gvvWo80y+VJKQKYUpHVxbrEyYOd5di775pS+vDfIT/AsswVUmaqBv
CkeZkeywYK8EvKKlcTQ4y1ZZOih/yjwfP8rNnWN4etmVvipBQ2IyK7uAKg5TzJRXsE7vG7Pb749t
fMAlH+Mroy1aQcLWSzGE4jWxILdOYgjP7Q0UgHjc6Pvp6//BkKKy81M053zrxAi3QOiB6m4kZtO4
D1dmtg7ITQixPXAHbEhZVenC99ROq6hKGm3KZ4Bn7jm7raLgi5GlrNudJsN6Lb4kY8OWilGnZVMx
+qe8EeXu+iBQKsy4g2qJ7fHVt76N/KrVj0q3qQwnb0tpOkGd2+3b3C0zaZONpFgREsZ+CMIot/RI
Eol0c6G0c2Co2TXnP3sPNebEc5CDHySRNlPr2Gcvi4wxqT30DImpM+lKWBBnA59KJZkMchlQHBU2
dQbU6MM3LBQALstzKjKdsAxwNSQdikK4E3nYvOQmv432i8FvWNvZIvZILvU6vWhOl1o55n0LCuLP
JeT4hIL2dJUAJQAVd67VL7tA6KqPvnvRjn6Kmy1uI5gT5RI200QV9a3djbkrnjApd1CgeSN8wF+h
6ycTTvg+JfONLoCETxfYyR6Fn0N0Ch0CX+MWKQK1bpQGA9WK3LpL/3Eh15gLzzw4pkoAKGXFu84e
WwBqyDaRYr+MN/zE+rDI7PS73gAqj9wz2C3LMyTWe2S1/4KYOH/08T+jWcOuDhrv1B/sEOOdQuDQ
DrtzFMjYNVwdDZ4OFvaWBbCnoLFM8GZ4SDUF+GgFdnAQ7dghF6hyfmogMzC4uC0Fx2bXj97yaUvg
crs+l337blM/Zk10QPBBxAQlvO+qdXyRg9Mo/t3upfurGpbl6TVdFnGhdsd3dd5zT1Md6/8UFaxh
1wFlR0xMJnPvqUjjJWp+Dxl6GvvlQx3Ep5Nq383lyGJrcERFBcjd5qGM3UqgvruErAbCRmmTmnMr
rwnq0A9kRCFTFF3r2TJ8qfIpVy19Msdhm/yIn4vX3a18on6Nwwyi/494ZOcj8VlhPk+adyPIckqN
GTDvQQPUb6V6L5rXQqh+Vh8hXvBKm3aZNkRis9/5nXQgSqTCUB/3ICC1YTeP1l9TDdoi0B8E5AdJ
jCoLsy8TvAXKbof6JwkYrcpOQ0Nrhp4QM6oFn/aihCsKMka0o+B0Yh2RFhQhOE/o6EgrVEOkldB4
S1LHMsNP4DRdAYT+0QaxKRfYIIBxKv7/jOgBPo/QVkf5zwJNMfXAdMrshw/ygiG5PV68Tlu152QQ
/Jd68o6ZD7TgUGlp91h379FcJk4QARcpzygYW34qmYUdsrs1+bC9aYFd3CQ97WZgwHcmDHn4fSi+
i//Hmb99ibI4B+ijRV62nV5tJJqnxCNdCcVigQm5nHprOOUq20sYfPqDifrDSA4CJoZ7VTJ799vi
TGle4e9syIDsq51BoqClB53c+KXu3a5Srwabrev8HV94rXGMwpxDurBp+DLW70O5bROjcDwQX+3H
TKYNJlCsmyVl/ZGZYepVhozK0f4qtHuxfuNWAfrGOIf4RvPLKEGRK40BrYvdDJZnMO5rF9X+Nlvn
nQ9T8sw90eMWwexqfj9szwja6DIB+E5945MGJ44En7eTtVyz4oqjycjQHx7afq8S0ThfFCu+JO1B
P5RrK85V7FVEllZOmc344WUG/b/RuKC3EETzxWMu5+Eu4uU8yGGL/ZF2LLczfE80nuHu/U0GTmPT
B4def4Ynr0nkkqFpP0mQHcaq730pBYn/zWhynglGIEeOQTSJQFhagFov6Hm2SRH35SHQ6FVYB4VD
m7XVrNI4kcJpb3SwEyUhuxj20x3AgAZYkW4yIe0yRfnNK3053Fr+/PDJ7p6SCAU5qkWT58JxqHwT
nubLi1UStfS3+A5Gr02O2T7tqwRkVxXeSV+3KlBcF+cz8GoXWd/YmRqa4ualfjNunzxv3cPRSXHb
/OrGG3nL2p3duCoGvSoYh6MkFuyE3c6TihJrL+n/mgt+apKFa2CnZK/P3yJ6rZXLOaC0xdhV+ZNu
vtqTsO1URZ9zZ2Rg4vGHtkhm2XZU1DScrBNZt5DaG8lo9GHvrP7780jR8E7LMCfQUVB1tOAsM+qd
VPWmMmy8p4Zgl9LDXiSwaqcpAhE+hrtmhJti8Dl+2U8TXYDMFtH5kKQSyVBnO51yGqqQwzqQAusr
7vbgyLrRln6QBGWNrSGW+72VvrNOYXyT8cpfqvWHtGc7vuzmPVA28Tqdl7GLFH4OshS8w8bFtYJw
mcsP/KhGtSPdQrhEsxecxn2vY+gCE48to+PPPzGjEq65fNVVvmjsNnb8+OmmJnsslws7OWGfFsyu
DRmhUQeFB/OMRyJKvdk2FTAVQekka8ao89ywgnkGvBo6o5zBsW3NOH5IhwMlLhVS8023/UtrtMwO
ZkYguzXNj5w8V3T7a70jnZ4wzb7q8ZaOzSlG0J4NwzsZDdUVegSYUyf/WRVCbjeZ/Dg0Y1DhaA8D
lE49Y/PQ5oLGMXif2xXWLXDYzdi2Xog7RoUzxLg29xGz/b1UBwZlqgUP5FVMI1o5lRrowHrdr6r8
KYNlCJHh5m/i4YXXoLvCVlUduxni7KrFYtB+v5XHJeB3c0DQdVK5Lss1iF4vjNArhAdUC2cBS84g
/8RUdqAGPYmG4FF4d3gNmKZkYH41fsMsAhkOiVY/cND/shIzrrrIhp5PvZyS3JDasaBOKBxZmeZk
truAp0ITv2j6Q8iMKxkqUqM2hpnnhsN+K0zT+U1dlwnkSG+UvKZjOmd6Td+n+Yg6NV/zm4zqUqvK
OgC7644deWLFR0/pcvvqyu+Qb7PmuIcy6EeugP6xR14O33GsQ1K+Tm+5vMPdqiPSgfS1DpXV2MCY
RFNEAlYn1khbdGbLKtCzmxZnR/wnd5Nk0VAHAHXSDqnOl2ZBMdbVcEIyZFglrmU2QpdwA5J6hcsH
/eSN1Hh5Ebd2cut2GwYGziirYZyBKFF4YSQ1eWLITxikuiKkgtFIpGVJmHzQJ1Dkc5OIXkPp8IIl
VgRRmp1vZsbDDVAxMvPnFI6PfkmxRq4pR3pd2WLEd7FwAGkoVInWM74PqJuZnMK3HyfMLh5LS93k
4/UMT0q2C87qw6oXN7WiKSngoIiAQ3jvl6DEwqEQybFPr8McSp70746y6prbJSVc40kxki+fl2ib
CcJDBmcRypjO9vJcTG/yq2IlzqGwgESr9u+cVIjiPaUb3GgTszu6Nk4w9tiuKyqTnewua+xVvAqJ
C5VFpaqUyAIPaaPh1GzFy3cHjMRyNIKC4w+Z18r+0BO8Qe0reAFxeMcwPBj1rmWaR2B23/b0c1uq
BKIU2SsSvyMv9yjD12h8o2ZKEheonZ5AGMHjYOIVsWg5hL7+ikP3azfsA7/5oLgmfPvb117OXMfn
BFArKV5AG1UE6ot5gJP7cN7UTvwZEuU1TZohdIMATiV7AqNwfRQNgouVG2OilbjTyEF8eqw5wuN3
LPTAN1gaiOQyEf0VeJTRgfmZZTy6cNfP9tiFhqR6NJj+XaEjQqz66KeFRMVo4+FzMvZK9J3Q1lSX
Txo0TV8Vt6hzsdM7vBUPMvYo5qNLBXHwaFz/iBXj///42nxx/QHl0gOCvzt1njgNcal0bxcpjVT2
ErDVHv/8Lv7M/gaopciARX+d2RsPWBo6vyHYsz+RdyNZ41rKSor9wKf68YnYVv1SkU0HmsUmUcGW
6MHv6/0nPLvCGPYV5lyG2aJnxJI5pmplgwgEnCtI5bpzJC+n1ygDmP+ol8OX39afYmAFNWCkMWNm
g/i5IBTsV2VdFWciJ/fWPAPZAXxwog1UB/vc9zfPpqnRFrhMGCN34H5/OqNtO5yMjgZn4z/jS+fp
UdcJwR7daatlcIoAXejN24Z/9uylnHmdfHmSLixamT1C8D37D/uy7JIY5V0N2zGiTsLyVVCqKtW9
anjRFQ0LjY8jMES/UnDjaxCAucrTT8CfAJQTQLEMkI/zK7Rxyu4OFPn6tL0A8ITr2Ecj3zXeZ523
thndTYOUS837e+ByNwkVZsF0j58uT4rCMvuF7+Dzpv3Q2R5NzAFEED6AjqreCDp7xk2xnzHvkded
xhBsBfaOFXFgjUxRkl5O9P2ZtDngXr9PZ8eDG3Yzfpe1cJBOrvCH8Y/+FS3meTsEzTcnpI00/qE6
Xy0b5TXoFnmnlBaqjrP0oTxwQW7rqVODion8nXeivympBHXGo4ld8ExHTeiwv3Rt5rYeI//9Sr5h
E7dRJS2/PFaE1Phpmoh464j9sUh5yLN/Bcbzva4NzKGPC7/LDKZCTT6Yw+c84F1vzpvmHLjqcoTr
92vryUJJpI23XZ3690uJEpLQZ5E96bRf47gy9d9Z2BcvFPF6tJGCbpYcnKrP6C90HBa737Y4VWjN
+nhJzWZh1MSpRSUql0WZ2+8e2Nb70D5qOvYIZBQ6DOSgvhKI+FyQ9k8I6/u104VyNIlrQI0jPL05
hqp8l4uhTAOsPz3D3ezjTgik9+uFyPoiHOPXYYNuxNRxfUbw9wVnoFqNIy2MNazXyySfP3n2N0NG
ejSLA+C0433ssWY4eQc12+SqJvtVDoiJyIV9iwMUZ2WdOwNGITXGA5Qdfr5CyBNxlB513XaFyuUP
TAqkepkkVCgde/v/TNOSntR7lXblwDSvWCjje5Ff2zV1TNtEfBDocJI73ZKVkXB3zMc8TYYzOPJQ
+vrPSwEMkx0opmqeZ8KDN2b2Llko4aEgnNQaGPoOJJTZ7bWzY9ZwMZsQZEwbtk+M3DH5bhVdwb7g
UuRLVHAG/mP2J1kor+vwF/1JqbbdV8biCv39Yn8cR382MAucVtg7iark2/HkQsUCuQduy2c6v+G/
xYlLokunMt24OdA+uddz0tnYulkcWG2IpOzgf+cugj7Pt0QVm1DNA/ckyO/xr+/9WgwVsMIJLpP9
yoWcgCB39IsRgldJvq42fstekoqCsg72GmMOouL4ezUbFTo02PVNdUeIgFPxNQVvEWdqK94tAAEH
CBCxmM01aj2zbYp+RJ269Q/0vTHCgC1OsJj6wXGJZMNblxoZnjGRj/14DQamHCZ1ksFwHQ0qzM/I
okiphQH1K3I26QH3hT7L9yh6POXUdngdB1oIFbY8i9xXCi6Y2Q/63or+qW0N+IfHhKhZgzEYRGvu
kTuFw3UZKOK3s2G9CKSV5BlXio2VTS/+0U1yreN8QojN3sPkqRqOGDgkKkDDU1jhCIPYNBBpg8LS
lSPjK8Yeasr/l0SB5qZNkTl8XtqqpyVxxrzdcErQsTpxvt/sMiWfGZmPREp4qZp4us6xHUJZ1WkY
moVGlENl7X8iHXiMGNVhgzMiqb3Po3ZO1oVUQ1zKNm9bs7ZKR44iJbi/4SUXRBsHlx8zxSFMwsnk
/L/TR0I0Z/c4hCoQDn30C1FdSIAZR++TcyL9vqODQVc1xytvV6rJeo+wFVTknjqHANqVLeLtW6UE
w51OkDZg7m93euzXsA6N+1xcudElSTuRjZzyFBsqvuelo5TPuHsTWliVEDg+l7OckfSmpykwYaBM
APbOR+4aTtsXCaoWCmVS+P80NXyjWifcaZVfjqNIyObJCn/A41j7EsmFBn3yqLBo9rjCpjRI/cF8
fZFFnbv3Wfx+2ezmJ1GPeB3YPWElW35C6TIbJ+lycpGLQDdECFGiBInyS26bNwHr5kbBAw0SKaRC
SFXITrrlPVngcUTyCeBo1WsKth+NtBv1LiaFDW3XNDJsp8L/i+QaXefj20cWUZxC1hohqK3RDIfy
Rd1xyQ30CYvNLbci7LN0cf6NwGmQ8UP4fcVnTh4febsX+P205XlS/aqqyWZMKr9ij+oEWzpnqZUa
2Bbbmb3NcTH7WQlH4WsiM9cWziip7Cbo5elvffnIl/q3Y33UMCQ0dsnwBkF54PCeMMtd28lXNdS1
9aF3xkXqgyhd7K5tMCZEyHLEDTUqyqkaAi9hGeMy/u8T7KISarPqt+MbA9ejeug0jPbZu28uMdZ+
RHedyGqBA5WMf3wvZzUMOYiYLY+A8MiGl3CqXp5A/J1p+1FJlq066sjDK5nnMOttDbDglUe600Gh
Zinm2orxUMUrfO9c9PHYHJ7GEOZbzIRM8noHvl5bSqn/5SG3hMnp9/uV6acqhSG6cK85u2H6ioHJ
/sMdYQfmJ4lkReh0PpUDk51ZkC/eUrjwTITF47KfPQZHC5mrybn/eFIWzmz8Er0+6agg1kQ7hnkk
fYrUu88InRVJQR8P8Q/SaMQ95lAaVPvJEyBoal4hmE3/RYp906YgEVhWVqILszY6II0lCBNHwKnj
OgAeVlx/bquHDHprCeUTtvDTQsvVvnA112xj+f9FjaUKvl7ev7LoM3W2dvJqJmPN66TcfFrsQBwI
ILlXKv35wcm3bQ+xQOg2s3Dy/x8FmrP5rURlTIn/2LJbVm+xF2mXm4tt6PHM68KloqDGkqEtVv1M
BLdv2f1DQ79sFg0puL49vQy8QAkqTsIgaLEGr7q7G+Xs7oRd2S8mC02Wdx6ejxorckdZo+EubWZv
XXPcZRsV+OQrhse2VQgMtPzqbD9DSocp7ycFeEc0I64ElnzSTblAioTc8whBiri3BDA7dH+16Wi4
cpB1CKXViIHKO5P3R8xnkQ9osKVVPIpAyx8U1JHdQR9lNILwXzcX7sTXDYNpufciFW1cPjBuXrZr
23sQUswkxTwEqrqoZBIbRXJly4U+Bm43A6iXuwgcc20o1FqimzxdhSpg1Bvs5MwO3ImYKn75kTB2
hI+WOadVu4AOINlmlZFlcYmNJW+ZVtUSuiwdqcGZ+gj7peqmljUDS/0yYnfGX4VC9JMoOHw8016w
efYrBusngH1TcGXfy37OyH1EfUU8+do8DX73Vxysb7Cw5IEV56Xjb7MwegFun+kZQU9YlUJy/XXM
VRO7C7LtVE1cOZ4Z0h8QodV/+5q7/g7CxdT4syYhtxqpt7Babx7R7bKhHukr4I5OJvxGhZ21zUBG
z5TFkeHoi4TiJdOwJiWR6ZzPuZd63xUZBnsMfaHMgLSbwnoWDV9Gz53Gsi6QvBRrkkGemKmfqfr5
2jnsxm2UkswqfLSOSnGhvkKXBFZDUglDYCJyRf/XAj+3bQ7pgTFLUTAjdapde9/c+85ZMn3kdBd5
E2mE30DuInzwSAIJlB5FuxxdKAyYBEXgF7gJbJjmVILr+0MfbGVYYR2OAfRWfUIodw+czirZHDCU
LWTh5I18YQ50A9f3dA188x0T2n/XlGX23S6SQgKWgtIaYAFU2Z6g849uc1Gg8z4e+oH446kQhlad
584+ue5dgirlJNZwX6Of6qRLPdebq9RTsuNADIjGWNwflW5mHDpn20nvi30TNXUJNpZyRBBJWX2i
JTtEPKFpTyhiaM9nvxgivLQyoKZCoBMJpX211OCAFEi/UmfiSXne1HauuygQ5jkzgplFfMmjP0ob
6kppZWmviDKuqtMYKyZl/nuAtBeKOkrQuKb8+X7odv5IBVLw/fFmxzQYSW5Q/xh2vEc4e9Hw/T6G
oHDVqTH1dCaI/ijaiYiBrkBtAIrkej+DzupHfG5USGWAWyh1S2aJrW91A4Ss9nVXMqx81/+IosHA
c4Tj58jcQZ7XsHfpk6gWurTJlqgVPXe9E6tu887Wcm6oFM66lW5ryt46tukxgVNrwq5dblG6kmRA
fqjbmabJr5vktrIdKO7prY1NguwZn6fl4Gz7ersuQrg1b8mjin2XzrvpjL5+1PEUuh9YltIjhsU0
02M+d5rga1OsfwdyhvJzTCrAkgW47xJbxIcMoeFep0SO5RPiaJNSiynqEvC13nI/yLkt2ixdr6k1
i2JRuLMieuktYXAoGm54mHkVj2SgAx2FKZx4Dl2uRc8zyvPDfvAsRo/VQSES2ZjbRksJDhbATw1M
Egjxfd+8FHG5NuNRscTs9KMZH0ssx0OvG7U05SM+nkO2huQIYzKMahM2PFrrrH03/7FL7j1yEAWN
fGG9twHMremxnY4eMtuAebF282FKcHUyi1nkJrV1mO5vs70EH+OUj1e64Iaeoe0YsY98GXQCNeQx
4kdLNnn+X89fnr89kRxQ8Z8+GsYcF6WhyIkbJS/O2hkJSJ4M8H6JAjcf7mRlnt5KceihgzEnOBjw
HI7R6rjQppYzKXx4GPJKlaVZgcrPl+IwoUMAGdp8v02hsCzDthsCF/5qBf6i2s7CqthaOXrGkJ9h
WpsLNH9eVpdkX8ETe/G8NtJklyEw/isl8h97cDBBYHHwRoLmm8gtN9sYStETcRPsZYoLxCoz+jOx
ciQ8IcdFsDyo6Hz9s99mziJu74I04UF9Aq8jvOYTAgIfDUPV633QipcllgCEa6axNwe8NmfaGr7P
eC0V5XaSLkdTJPgwDW561fVxbRh5HP5nMpePwZOsWwPpEeh95Ow6iihkhNWdQS8F/0AONTUWsJZG
vcsW6ysboGxBnLUWYhB03mdumO2xzwjlbQ71FQ2D8hQXckxqjaaCef4IW3s9NZxLdK1MCXb7IX5z
lPSZwILrUC4CbGQov5ZgowcM5X/Fpfeiq6Q5jFUxn5yfp/eijxpio9LJ0wPmbwpa0IC2vmGj4oPy
B2teBJmbZ1SncjIfncGabZt88aCsGF7JUXPFKqGcIaJldc7mK87BO9yXofMHmx3QaAX8JxGtqb40
WdzKdIOGmY0DPzYXWgdoZGO1gPhtXv7+FnZGVMKVn+qI5QffzxpYuHlKkJYF+n+usLRRl6zgeVBr
EKLz3yRkPoIRnpAA6PyKu/fTcavsgGpEaDBmk699+1quWPMy1wyUfY9x2F4dHpE70VM0YRTLI0Y2
bLnwq1ig5btXd1xr/2Cbje96M4NqrMOyd4pNGyu0X9US9wFq4FOWDCSCAViMU5jMdVmpvn42M7G4
G9QrV6HLRuDn0+no0iOvw16hV0jgdrLaa7/oUzr9IWuGJhtL2TPJHAMf5dUBl1yiyEIcvGBInU+g
Z7iCq9hmLBG65oiJQzXlk6pcSblr5izaGBNH5vDej61RDhVRQnKC5+cBhQNj1Nxr+p8jXRrYafHm
CZD0XfKGqi3JE9cBdEeG8CQq4b2jIzUg5mxzPKGy4R6Vy+OP7qUcA/+CEe0K8HWADA3Rhwt9l95a
61b4XDHJTpMigEO9yvh4UJPGwF4NRKo2CyFtE124FScFt79BvBw4iCsSpk6D3qXqj19U7Yg60rbq
7uEQ8fyt+QPM32T4C3A1gTLfUwZz2JKkYyrIaO2VAh6KxQP3/jVj75RXaY5LBqCSJMq1oqm7UfQx
kN3qXBvQElQS4OMFep3GT4v2tKvvhz8puOlExNKGA6FYEUKR8k7k43g+R1RT6Us81vy5SEl6wWVE
2JD8/1mCOcRVjXa4kCVzMOuh1dSM7FgSGVX1K4qGNU5/xj1AB//U5hpeUya2bmEU3b3RRLAX6L9W
PWTDo36XZGr3TQWK0GP8GOc6u90O/t9Lt4FACqKPmkZQmNmCI2zFxJRFUX9MimGd95cUoRXovWYf
3jazY69KSqTMxqNSeY8CqF+JtlFKtsyh4evC5s1UUV3mJZPTEKyAL9zypFe5LpMOlXOT3SWHgDjc
47PtoSfZoxDgsEsy4W1N1OXKESB9xEzPSAdGswEPFg+J6xUsFgeaIL/5FiQw3BNRJMpJ9Oefr6nq
r/19jn8PYOlU1FD14STRZS0r6mvv/ArZRXNqP+7gwi9BTgIcN2S40MTJv/LyHIBzRldECw257bup
u0blqNlDKdCUSp/smE70Q3p6dLJQOaRXIlREBhtifCQx4I8ctKyAzkGws5NICtJWQLApcReyKeA/
XQQhdM7vjdvpgwio9RzsYuq6i9o5wO26hFbfW/FhbKBnmjj1+QrLzsYfVkkF1Xdj+Y86ELT9X6LL
apDX8UpG/tPmUvdbQb6ODZYYe0mMhjyx/BXFCoVh2ON/E2YL7njX+wbeXs9MPsFSZdbcdLWHAgK2
XkvG/boSpTNcCTPY8TvPoKe2SBx/i+egWOcSD7trpzsyl7kN0GMi0EB0yOLj/YA2JSlQ/4z6qy/Q
IH/S83NdxWoFoNDAuoskGHR/aYdEnFKxQx5yTr0WA6nhaXOoZar4rFInePDjpQe4Q48x8rciFI2U
Vj+TkltpOwLtnsl/HmAsBBVgajf+uI4mC074NMHJh/QU4kJzfgNmJBI/+juA7xOsftZ7hR/CQL/7
vy+I+uTC54MdsJul0NbL2Y6Q8j2dzzvZvHDMOrG2B/3opBlznoG9C+aVDb+PCqabdMKcXPN132qu
axDa6CnGVy4GLuUquTzFDf1vQ4423e9mEHE7zeNKqI7nD0TRDjk1W7Y13LIuQu5ICjt9CCJdUmKd
ywJt30FtMsuiXKIaqpIWOgF7sDZNXoGpKzU/+NPpj/kCzOxAjj70uWHlmkfMwtL5dl3fk9uw/Q7p
iJ8z9EyN6O3CuXY0XrzV/mf/WkFjqc+DbaoqtHS4EjUEJiRwQR+n4dta3EwEGa9reHj49vcJv61r
klls8UfqF3r/Nkcybrn745fW11wkOsPV4LO5cuzJe2kmTSh4+Zkn0xQ0DfKIpJn8RZMYpL5D06rz
4zuOP3BIayiCIKlJo9tY+JbBWODCQM8nEvg6OPTxhvfnkOgBC+6PUCbFf1p+yy1hRXoGVaXTVHx/
+XEvdXcIDd1DPA8wnpNrLFtf4M9PVWKT/Mvwkw0f/CjLPOIDUCVid9jYJ/UgW6wbFzDhftkxjNQN
dnHJRksFwLPU2JNNGlGJmv4UnT7PNIhd0pKaJhdgRD3YURZI8OOvjcKPmziIPy0NxmkU1L0dRnYm
ET9cjmrraD9JW9lL4KF0RtgunOmKVTBSAqYa+QNPqTYk2KmPxmMlTbiOFNYFCATuN7KZQBBAdO8p
riqYPxaV1mQgqQ+NFA1Pkcz/Tq6ewnVZrtHstyRvcVvcyLG16hsjrbfGK0O1SxaJVLEZh4yjaW3Z
oisQ1n9JozhqdMwod7ipYPjdTz5jcMrNgJ1S2DClJfdA20pY/Mp4LwoQE1O8Y5Bwow6CG5pWFJti
hIx7Chdp29MkApLZnybNrkdm0+P+dsfaFQt3qoSmrgaBw3nsVMl9n/wQOa0oEPyUx5/sAyiv9K1e
BdVRsc7I5SabjGt9EIx81ytCvcIku+A4djb35LGE93fXjGSJGEWGVcMFHcfIh0lkku3zd3FFaxST
R6d8TBErsbhOy1vGi5dlHq1KHhcDTr5Nvw1eBNmV6e3L1R1ySQ1tw5zcmhzE4yaGBbUOWMsVUvUT
J1YwX3PSm1lDCAKQ0UL8diWCMPIl5WQuI2yYO5cyAa5q+GngjdjqDkSUDYpqBjwtS6g7x/sbe/rV
NKxiXI4yOYWcwo2uw+Kr7f8PSVk3HqwZyeRnQcwH/yusZ4zZqaDfeDH/qSjuuVqA5ilfoUIBysnb
5ulcXbqTdmzy/kQ95ljbMPr2lnOboRozUpG9ZS3uLAKVISuvPuZY9fFtZmGFS5+90mPnkBx396Lb
CKUZcommgph/ep/nF2oOhD9baZ3rZR9Bo1TkMNusvAwNjjFV3o6ThrpuBaIpaFNtoZlVZqQMVwNn
jxCGyW/wd/X6W7LtSDij2fkxNcYfGoyhdMxaZJ1DyZPwWDdfjRbaOlXHBK9r/ikcR01HTWrRUDBa
cDCYkTDFvgOAUJWJ58PetyeTEqiahm9GO4i6lkARODsNsI9Z6mZANUBrzMBB56P//cRhz7NtZJHq
1HJQNdt7NwrB7p9zlbnAISOJlJQHHbTJszaZgWt3ThaTyJG/A6iXL4lVJZjXMeLblv5wfegA+60h
2AwHYl4moR328EjZCy83pWvyu6lSR88ANfGPu3X8f2bDcyT2U+gTQuInjVFVh0ePvyxU/4KAozFf
/t3VrZOMExjNn92L4YFILnT+oJO4FK4lREFY7Hj3AOsHP1j0K+d+Y/L82B32lvZDTeQU3aKNESNl
PrJ0QRY6eiNjh59Ixf39ahEUkq4FrrDhd4bPFLJwgDR+vhHPX4P+UK97KVEullyKx+GvZvS2x9Ip
eEnBE7HRfS20DUCvpdnSe3clO+mzM1U4+M5VVieqaaTBxSskwyCtJFdR79ASgAk9roAemtWCMOSU
+u2tcWeXMUOHODncMKyMP23iR3IZvlbGlxFdv3+C3dL68tzCw1eBBXpBYDY9CO7n+WYlJ1Dy6zHZ
h2uHYdLLfRSStQFx41hsI05jntf44z8NmoJfK/tnU+gtU5O5qU23uAriSkhWkFRglo0zLy4toV7u
1qwRqUvJK6l88VvF4juSWMXgQeIKLJ94eBq0vprvEpYqCzb/zotQEkkM4p00hUtdGTWx95kGTkJA
/c1QQQrVWtJFNpFuSnnBpOgzdJSeDAyIAVg8jGtvKdF9q7Ae1wBWUwf7XFIIgrF2vqnS4jvFI2yM
9dAhNvOoJVsYNJ9ebKBcNbgvSdYqiA4TqqfmbgsbEUJ1AlHJ5SuPe+UschYn+EOt1RWYQAtr5eP3
bSRyWsM/bl5duV2Kzm1KE++RLJFDDk0gxCtr6pLg6cIgqmtGxlppngOqKMP5trn4NOd6rwO3QUKJ
KlA6/AJmYjOGHCDCiNhbCqy9xyECA9peVln7bol89nBXNLIR53GtF6LU82sa2DMnNuiWaIsIVH3S
IX7r6hjMK+L+YAf9FvVwqvYHW1pKtdkQaNREynENL4bTU62tO5kExUHauxzsuiUKR5XkFEY9wG8a
xfB7Z4798wBg6LtX2UgrADBtxCXIn56TOzeKlCQxXB/vHziepew8nC/oxxv1dTWrpVDYf1HKi8nt
N60dyNH2VUbjlmGIt/yPNVyDi1E83JHZtVCtbAYIwFm2rks6cdCMjsyKgwPSo7PD77TuzddiSqJR
h0rXlYyxDqyUS7ncJCCXuwLqm6qAZvV5vcMJI9dytPs+HlDOhEx6Ld8T6Fs+GF5agdSvSEyVrGT3
++9IQaARtsAZzTA4HeHRE7gVW1KZVlPN8DiRHLvF1kqgd5dpn49ONpffPQrpDCd9Q+sBhBRRg4RO
XgOj6MfLgtfxg0fijj7xhjjFgNdLV56HJoijMSUDGG/iiYX6d6cmBAZ/RbmiLowRHNo38wwl9Thx
ckK3FQ+pGGxrBLcJ1ENOV8Dge1ebGN0GlFhTeml6J6hiKyK+luQAlpb/psY7xskbVCFEhxijs6S7
PYR3BxPTLBvNHTwkb8S6N3/MbVfGtqFUKuuBIO+JoYJG0sHKDtoqZMAoVpsyHTl0ndydXzBRdr6h
ZRVA5xgE29GkpdKnNxja6g07tOl7b6fo6B5VRWdTWViX0GR2JJTdp9sGayqoxT+Uzux7kw4ZKgWP
Ya0kOpfheUUiT8hPpmgobjcWLLIJQsrjuDboLi+43uVnWXKcpLEOxvcJ6T4rk90Aquta4Znm1mOD
U/yt9CoBA5uOnuBA75UUOJV1A8aEfbadrWmJvY35EGKZ3vxxq2BNIp7V8PNMqkas3bbdwcGCk0ik
6c3xgV8GBxV8o+AfeyITeTKLUnUSowGerdmBItzLXNz900nxDkgl7rWOoT0K+BnJ20KKExwfKD6C
2NokZuehGI6pRRNLDq1r4eSfMvoB1nkpZhVrNCC+9vnHGzW7AUt7G6xlLJF9++k/jbRLv3OYTX4I
Odb2dWWoU/RBPVZ48cYMG83XkAEwZJHQ1earulpg6twqDlH55tyKhgTFoeHVyIO8WvSev648fQqJ
s9quHDLWb0KK1YnVhR0taLPPvpQOR6/M8NBz43zlNPxv0Co82U6R+w0drUOMkrbEnsLtFVJwtTYp
NQksZ5g91GOcBwqUuNpjOmnhRLqC4UzVAcGg3j7k2ACt9DhE+gNSJXfDaBanU2xAF1KvefwFlJow
3oAlGNgEb7zqSHtpRkU2Rlt7wJkMfH/F8WYE6m6ss3Y0J0Mc8VhLabvDZYLWZ5uiY1H1mU6ShZgj
tT7bu6r+iBFXWmaInWb59CJ+LYkcbbyO6+tW/aSosgPhxc4OUgqdtnnpWHynJef86bmfY1txkJhG
XFHO1AW5fddMGZeBPzxVKgn5uMx9+0xDP8b8co7q7rXHmVMMAfDxPq3YcFKVgMLXExEghu4HbImV
YKGDIPq9S01TtcKJwjQs52LIYyY2046gwy8sSPZFxjNFD2Ri5a99U6+aLAwkMSTqGtfWgtv6zqWM
2s61cSK0W01Kkr1P3eJrk3K0YxLFF9uzmsXsRF8wuaTqrY3et2+4PQ++HCIIRehDuDEzkikaiqtS
kBqzA1k41O37nUfF04iOmUxWxONACpqU7hFja0Neihsu7z2Nh+s6khxID9FNDNEmb3wtOVHrov7S
FdQmU2E50HrPTj5SWdMXQX8oWj4x7hbPTQ9FxXBWZwJn9O2N2ENCepqasgKO/f7gQX6YbwFM6PZp
XfIV+aYTQhfefC1DC8aXpPs6eFdWmDehQeD8SC72x48fq0F4D9yk41b0UmQksvwt2AKCnHfMGqtk
7ADwPWfnJEetUBdVN3yJt+3RDbPj3T2LIPe10Z5+FqXfcQwttq+YaqchEeYfw4jNYKp39YTp/yZm
5vKkE0tqAkGhy+jLc2SROgyEeuMqqT5B5AwSZc+bF1h3W5wFZAKDrnE6KpX5HdGixuZIJg9Mf30+
ifMy/CRLE3ZxKy0lrPJZn48Uw8m5vt4iccphS8X+AB0K18ZP0vJG+XLREZCR2zmVGciMjNmYGRts
YR/pCqZdG1+oisXtNrYbj6Pvjx31c82urTXA8/ZeBCZ9AFZoAw1bduvJWpPR/bUcHG/NFtgwgdUH
Tf43OnzyGt4ZfWsq1u75KKEbXDCx9+gC1MXDZGN+c3AR1+sVksJRq4FT6lKkBioZWSUyGSdf9xKg
j9mnWpeGLgNUVfk2GGQzSSYS9/uhxQtIdUBTWdp7KtSVgorJ4tPDvhf018+UQbwkiq5gjf9VP0/0
8mmoj0wDAIyyRrMBqZTxEGPnzdPhaZbG7o4PwvHvl+wwNxXfcQciWZIO/KZ08OnYl1H1SmBurxl9
v4YZ9Az4LTLQjNGp53or125U4U6OmLg4h3fPuh0JYzxHVCSJoHv+JUAVKrdewPGZSXBPd5mEjtql
ojJ4QUUFnKHKWoF01POIps8UsSMQjN+swaTLLVRqqUDxFGMTxy/8cTBZFZBjIWsCi7YDKkBGbSGQ
KntsOGhWom1sfYN2skAUKXXRwSoQal4479kcKwjhCicjqLF8duu4FmEoqDpADm76mE07di+ApLRl
9E2zIRhznJsUT+WfAX0wRwWPIklQjNonOvN/VhYyt+xbI+J9Ja6t7m/ZUZfbC91N0IqIH50ygznO
a8wY3DMC/wVvIJIRm6w1g4q8UhLW0vozot6F64xztmuk9TDzMOqpN6/wu6XpAvJZNx/hq6h6vwZD
fqbhpBh/rdcTHa65fjnfB91B9fE6oOD/ZTp+V65rdUymabWWyQ08PA9QKMWWkq/Im5dCqvcBsiGW
qSsJEPGtH8v70CmNQs8AtHABHxtsT4Vk9v82TvS1AQLQfnxcOAfmwu66kJFKpiscDqtRSH699kKC
V+aye11nlZuwmVxZCnQ5Usmkn2heGdVv1qx2f0J1DJtdv3ld9e8S0Zcripb3feBPEBwg/lvpxTC4
Aag+wdSMV0lzIjXL5+vfhwztdnlPBXWQECcTe7lAX+VfyvdwzVUeLBeEs6KQdEZWr5mK0qBBexX4
lpMtWXBCvl2OL1/VjEka0kP5XerwQH6lYa0fxbY5HmbPn36TlkbO/gVkCPYj+RFZe0/PHsr4OO1q
jfO7rrLpc5xFnf9cP9vDrxfev0eGu1cA8Jmzw3e2zgWZxGz+8CwEMXkXUyeQ2R5MklVxJvf6xL4/
cVVDkEHudtNpudcaRy/4uRYewV8qA2Ufc7VC7FvSK+1SJ5+mqL/4N+tK3Bd75hD9YFF6s3ythVzM
rlxBusjYQWXbNF4LuO79WlNTlcY36CvAU8g2+oXliL2BKMTDl8qqxpeEXVjpLlRchXz5Z8EXim+l
Ss73gh4AzSkfcinB+KpCZB9OWiW6/6xjA1xZ5tRtqNTtGcyrEGvszFTnSFHRiZPqD9bHNEzIlEYm
DNTctDTDhDeHUvjnCgGjioQLoZISVDfv7VJx8syyfLkIMbGFOAjvo/sgVf2EzyrNblAlEwxM7tPl
opspZL72/TCfRePaezt7u2uiErX6UNmmKpVQOj8Cdiw2rdvQvozVfEKSGgR68VvT/VMcC3ji89/n
Om5Z8eEHntyf6hgSWQVxKyzfG/uiFi7+TOhem70H6bR2G+/iwLlU4vaXR6gAFUwz2cHUQ+ZLt8eH
JzEfw2pajcp1TsT7Uvi49XzQVxt6mzehOOM3BBdt1DwYbpfbaxW1m4ev8T3auZ7XkgPixNCeJP+Z
v+9IFsKp2jg8F3uEP5Hzn3P6N5x1SLi/s/mhV4ETcOLIhJLMTX8mrLqAqvKamuPnK2pUUdRoRJP7
98QflWMGcSlASFY/mDHMHwmKPDMJzhlgvBBHqMMzE3dV/CvIejJ8y0MSi5NOaKOsjc1Kxnm1V+1N
YH/WsHSu5N2G8hPZhR84TpDy/1am1UA6nvco7LvHQUuDB/9eQYlddbRqwcX5iWCL1zJN+/jiRnNB
PmlI/4MkRl5qdI8reHTDEScuX+/7U9ZpTX28BBP4hAOUDt+oDGoq4wHoTJBopVmrEYCKG4c1RUg5
XIG7mTvz8EkkQpbkoi5LAEbC5Wrl6X6+lcmg0A/6nz5UmnGnaEvDKVjMiK4INq+A/2rJijvKOaJl
LtM7qX2lvfeFE2+2HLEy0hysBEGpf8HWdcRMS5EtmQEgNQj7HSC/XYY1sJYFm/1wcqriMIe/5ow5
SFQkLpDDcrwWa1DhxQkwDCKkXfgxgriPyFmo10EOGsUK7M+CBK7ilN/QFbqXhUIWmKp6nv/at2R1
7bmnGzq0LNw7g3OjUiJl+ZdPkQHlSsut9IMayvbKCdoDey128LTSt2t3j1VoxsoGOg/3YfrI4Uoh
/8pyk0UPbZ/D5MHLog/LuBPSnA2Pucjea05fBFxdb4lXYJ30zrYnTpP/Qre0Q/g5HeiubS3yulXN
QZ/uFYikGzyNmeMZLIgZmhUthClXnTGQ8ri/mww2FHYGZJOCK8WdF5URwzTc5l+DzNbXRcCLghe9
Bh9FovOlKHndN1ydp5EYGxC7lWdDOssE5xGCxIZrpVXOlFbtsS1y71ruobsEdl8h+AUiNfQLJT9w
eMf8y62LzoufIKETtQmnibmZLAX4vBnyFJgSYUr1xiAMk9FKh00pZ5z20tJuRtV9cvuX4gxhOBKI
mKKbxqHBARIW6nA4lwRLVCefrzMdKOHbrCF+FsX29GaBxCZQ9JfjY3tlC6tsQzj2aE349ouwHumF
FEFM6JkB0bb2AVyQIZP5ODhXPK/8N7EBcZLQH+6Zb1/C+giEfRWTthK9BhvShJ7SZq49kHBgf9Jd
FzmMg2eFziuOOWlaSn24KsUtwPK7iZfhKIyisQeN740d5ilDqFVAVE2dT0Wk57y6H1H6vuB8Fmvn
/dxwiiKCmp1Ot3trS0U+UZ2xuMu+DL2NZGTA478uDLEcuAmyPQvoWhNJ/EEjmGfcYO4jeD3eBDqF
yl8NRUYejKMdl3SU54HSN+xpvi0MEO1LDPN5NRFwQIx7DgpUYYCW3akhg/0R2M0HO2em9Xb+OBy5
NYLorSqve2e/9He3mdNx19VYE8lqh7eW3bLmsEKMsxCZQPO34rbNwKOup+JbWFoxdiyJ6yw1SOiJ
HXTglN6i++Pj3Y7u1+1gDKBMJQW8DzLBnRUREoQrEFpcaJviHADC/6OrVgZGtKp+z75h4Xap2b9F
qvnx0tttrOG/jWJFwgDT/kqJazDpfqxiWsZidkv+cIBQV02u5NdlhaRO97gYfAaQPgt/dZWEf1WZ
2MiLRPV+eKzSn2RXO8v5Y2KxrpBCUF/aLfPfMyh1LRUfrf8NS2CNQNQDNf6F3BI6QJ04AVCqZLGR
pkYDfYL13C4JAAUDUjiB0ZRMBFs04zflh8BCYwp/+E2GjJ0SwUnJx6DoLjnXHJgJ2sCKlO4baGYf
Cas8/a9TKb8goChaUPksJ4Yeibqz+p5+N9NdJcaPSgvVBZNbp/X5sG6HuYMqJVppLT2Uj78TC1zK
Z3laUSwjjDgshgBJ85KtdIQI56iU81FYnjNL2F+SSNs9vt1DjlCOWzuleThlzwZ4L6AxVh6M8clY
eE7hc4M5x8mkA8UC3TI/EVlQf6dBlmEdPYeIeaByyfPd5a6GBSLejnJ9y773zaGhuf9pc4H7aKpC
bgB8VUBQQeeRgZv196JoYyJOpJdZv5kPopMuavz9g8ib2d46K3zzNxDNP9ncWvUfttPL6Th6ugmE
8aFTfodS6RPg2T1ErPTWK1NvFWlURMHOOC1mqLPGdfHeWnSymTnrrth2Jhb+7byZPNwfSBUC2Dcr
trDflS7OggPIUprUMZ790ad1ByzydrVfRQKkKoW2AoeDIAgaV7JYQSBMIk3utq7OwpJJ2QxtbD+H
HJD98whmd3W43TXCvq+gUIODkGp8QGxhFIZlsU6aZi88ocHhCOMAVSp8PA72kzDDO/D7HRpsFG9x
bDYgT9EnR4iOwRtJH26z15nVcWZErTjgzmnTf+OoJzmmYyIhtS1Yylg/vPRtX1Q3ddp8e2+WNhXC
PrLs4Z5BnPNWn+2PQoYBakMXeZenteLlViH326+BSXLettWd0VrpGgGW3IDC6rEJN50G8g0sYOmf
haDhSi36/3pOJb75tTYwuCsnvCeUDLe8ujut5d1NUP+3Ay1PEP3r9R0FGQOECwfUFFGKUSDGcMiL
8F/W2WujBUQEyv/jxm+OvhWi7FAB0VoakIbg/2/86St2R6rMFoPzUvBFzB5wFQJ+dTPozU21UduL
50Bl8hvbK7yvf9iSCRddd0KstdMZkxD9pd3jsDq7ZjtpKRblyd6QqN+GxSL4a3YTIDY/htavhFb7
yVJQdv+AToUPRX9ZqguGYaHSHa0QqRjkZn9bK4JDd3b5brvRxpExgEjzXV2ipMKeKFiDxUwHb1CY
Z+UwnAKR23RH/nU9NO6p0/nmt/HxgqS+ecUFW3NMKni911k3vshemj1xqPWB1GKkps6lzwS8bOLb
gAO2AfhJNqNdF+YzjH+wfbzflxg6/EleIkxJpUPWwYMtxcjeUGamHe3OsJ8nYV/cehPNITKZn4kn
uyKowLAs7LlNq+Nk/w+NIZ80K9NRVI/0npZaVN4uGmBUVDFWNRTkXz+bDJaT55R2igjGalqDJH6Z
NTdsxJrhI2rnUoxIHoxo8BLO6GaQuT07WrjEOLyzUzRxMdyfZXHmceVeTsTrYl2ZwK7mZCT44RpC
uspuxtXfR2EFx8tgUoeIW5nbxD3oW7uP648SegLredAEAYROTPnrLNKdVpxrIGyg6dBv9n4VWbEf
i0Q4bt0yZYI9A39kYDCmmlQYDk+pfUqZcbLU7C4IAg0iFvNa5xLEocJHZKK1swt/OYvrofWjTOD6
Mco155Xaq8pO1oFJP0SVp5Ws2LI3SvshKVg5MlZ/mpVJbS2Rl59inw11OLf8dkWVLDWHb5d+OpAe
T1sRmNFqVDAT9Bsd5wzmQRO0eTC7qwPhfkSAxxilnxb41RoPlqV7okczSLi/H06R96zF7/maEKDa
D/k552d8LfrsSwIeDVA9QXXuacMTTMxWjlqwzOgvllbSnWN5A9I5TcqNKYsEGiL0MFTP97s4+yzK
un4SipxsB6B1wOBgEdF7QOzRcvkix1FNgwYZRAadWIieOS8MHJxgrd0cbA/jEbxOUJ5FnFVXwCiw
ecicAjIBcLyNmRGfzj0FhzOc8SO5WFXEIclE2jK0mQS75T3TL6A5sbKa6R5VAHR6INpRRKNGQYOA
CbbJqq2SOpiJEnUqjkmnyoW2Q/Ms0s90ZCWGLXN9ZI/LCKQiY73Grt8cl22jKQRrP6RkCoAG1PY3
GatAmQmFrp4qfhI6VOYTsinswu2ol1oLiDjYEQoODmaJhVeMUypVsjNuM/dqBn9ZM3Ije00dKW1A
XD12j4si0O+4Cp9HFPZkHioJsgB5oDrdg88vJOcJPfMc+zrWvqPWPEWH36b1pXtfwhuknpiKILW6
l+hjWx5zbCmPkzIzH+vP74JMMxxJytwsPSrsA0CU9wZfMey8HxpRfNhr/fEYFqagzyfDON4sjafU
WfE3HCOVZKQJm+qdWZr7caEdXTE3HXWLqKm1F3vTkhPXU23ZueajmZeHdm9L1EfcYLE7qT7iDAZW
3uuGpUkoSMinTV6iJ/54FUyTou+9/7ib2yPxaaWCjI1sdCKNV3wfzp5/CR7/bc+xwHN8CEXWpAnX
vC2rZMOueOronMBQWke4TQvgg2ZDw+rOrGFi5j3GJMx//R256hC9IgTDWNpbq/HM/yM2Z0hir/hN
37k9nMZ0NzO8YUfh+07Kn9js8qLYIeCne28/C/sDwq0qoCUMF+kr2FKCIXpdwehnCuUUydS5hu+G
K4f8H5IOIA+oK9S7udwswYr/Nuz8voyXaQVt881GcqUPyPcwcwgGKEKYbh+khUP0mPRb9DlGOs/w
nDBCEclNzrDmpqtBvOiCfRxeFwBDLDUI2nGViDMsOnEzcQjvt3HE40lNAv4GQJoo2v06uoQAj4s0
u2eRKKl5irD/1D4gIbRSorqi49zV8Te4vmcpLt2iXNpqpD1uMbg+aPuk2mQhb1aR4Yb2J7QXppVl
IAvmLd9HBHWjkc0sNafWXpyfXsyZmTRrza8HbXBvHUMQ2HblXB2VtgJcQIceCoMTpOSXXjjuJEtJ
UqD/VzbgEXI1O2eSGBic0Dnzljm33tDkgpYfjefLyBti+Q2xVx7yw0XInSleofkazU4V6uGKdRqN
gGBAXFZR0QBhsFf7peMFDoDgi5k87wDuosU5SGfuFGUginS0pxn9kbqI8uwhc1EdOKKbon576tp+
VXNHeiEeiQuw8974WDN+rwLfc4nYfg9hGItBtF2eX8Wc2X5fPZtxO85mIplBFzlZ91bQS4sGLrIu
3ihVhH0Rf/5MztR4VA7o1IBmS5JCkTELvUWLBoZBpEDgCz/Ek78hKX/f+E3+YLhCz9E1c3C5aCi/
Rbd1Q0ipXG2X+uUB77DgCRD5isXfFGc07pLpu/Ylcv5dQDXNCTVz3LG16INChF2RiBQFXThUid/9
KnicnzmFUGeXMhA7sMnGLfxMmqSwwgkOq1RAVx5JjgKx/dvK2O3PZBb7BjbqBuu7E4F7i9N2fSe1
pEtz62vwsu+0aS05H8bJaxN2y+zfEXXOkw0nAmahnf6qs9Z4JBmAW0qvinmJ8iRDpzZlkQ4tpTFe
oLIaEMTPU3oUoTjnbSKEkFUCwN036Jvu5v65bnVH0WxXbM6hmPnMWB5AXTpP2iKoBOSPJZm1+Rlw
ydG5b2Ap9UKszHZ5GCm+61NmeStdr47s2q/gZGJ4ABxGuSVGPJ10LMgdc1LxamJks6cVkmOYc46+
+0N9BX7oGjDRurVEeCzL2eXowjs19MaIvpjQ1gc7vV6MOEIKSzFfNdJBcdnAmLVLayQvn7WwSTZY
sw36AHtQrQ2+RLhUr+uV5gkznU7UoQLcHUy6kc68aEigRYE+j1FhOhestwKkyTqLFEfPrXcIIJM2
eVkLcm98sQzXcSLagImPzVHd3F2VOTzxQcYMpV9IjDPAl8CMc/eA7R8/pr0WtxRhZfnmrkALHQKT
tCIy1sS4+zPFzOEXzXv48WRvfs3iHQQ7BSXEu+EN2vLeIMbtvmRbFQHoTWl2N9NVEw82WlmzXWsc
/ukvfoITIOw/Zo3G/Xthu79tmpcXDPSD+ox1vATwIziI7XfqgRfnv7j63FIAqSfezDVcsGaPip3y
5PD9RBnLljASwZgEjlDLt5sxjXYIDqF2XA8mY7GBE6FSP7tBxEyDn0zfqOr9MhFRAEZPwLg7r/rF
m05lkfizqMTwFHAaENu9XrAuoa7seyDJYiwqQ0EKZE30nq1yXZrytWf1bRhMyoIsJRaQawEeG0Gn
TRsgNX3F+GqTiXmU2Vf5XJszuIyyMmpOzxKU4xMrQrnHpEYc2TyPpoFKORXYAKNrJ2nN9/qXZRBK
ne7Wndtu9pF0FMa3foFbebcHdeAQyVQvdWmWxrMM64fpvlKumIMtFKn8HMFt+8Yg8IRThoqy9EMv
rdz/JNYFgYb7THbSWowc2Rt619O/BnqC5d6LisoJaWY4JM4ss96dPXkuGvJ3t3BrewKgpGKozTdR
89dXGjwqLUomYt0sKWt9CgSVSKzJ7NMj2wo23TActv6IyuYr4DElqzWH+PbHhIVQxexWEF0tVzn/
iimntv5Vm3N8+iYl46t4lSQJ7dz1ABeFyOQEmOkOAWdOR1ynUoeEvUrvIBa9cJXD+owGGhDDqgw5
TUeds0e3Fa2aBD1T57GfOPHqcyq0Gjp/ynhIX3AP7lmz3GeB6vE3UNLyq6Um0h65+mIzqc6b4TkH
bXpJQ67gOOv8Awsb87UEbnIQVryK4iT5cW7mLCjr9o/y/dBaYWDbT5CIarR9DQOGBacKwfDkIi9T
0WICnihKq+XovM0NgGrvtLccP9I/gGI4Fi6M6/J5x+XvLkk7zbfSrMgqwRzxNQ/YeYYZG3COimrz
R9p8zSikQzTTL8DFzsVriSBdm7F164VvUd4NTUzIJY3BMJ2UyrEWYtsh58KiaSjwr3k7A7t5eoXW
wXQnOvdDDCqLSz1884ysvPsCgasvugnUxB0KE1N/fXMk8EWJA95sFlFCft2crURtzgcZPuuhvFIJ
4gDG5npj1mnsdSWuoh8HLJ/xXpSxepOS6W9ZOwJT0bN8N4V/+f0fbheiApQurGOIUXwyCnlQMcxN
p873flQ0eYjt/um7oupNzttFiy/hlGVcom+nSuGFvikK6NA/YbFyMwYX4JdgQaVu8CZSro0AWg8A
gukS4qS279lZbbNOtsyQkUAB5QP3+kzZsS4xeYJAAc3opeCIIrzZ8nvsCSSQp222Wsp+POm0GYAX
tr7G224B+hte0Ex7QzZjSkEnWFn6MaBbk6E8bfrF1oS21rZa26CIirwaryBBQXAJkrbmPeMyZgPn
RB3VqMT/YyPMDD4Qiet6hN4s+mZ+wdKFOdD0eO/mMxQnulQmVxh8tIYFocSJvovLElPjllHsPOjP
BCrGjOUnGTxLYeyZFw6qsbEqL1ioiuFruD/rN820JkRFvV1Hm/WSEDxssmx+TPsBaI8KwzLcVVOd
w872uf8IcgMbr+CHAt3qdjNhzTEjMOAf5vc3b4ibBO3TiYGiVjVrYg7GZe7nzUA5cHSsAryxrM98
hZC5pTSRsjfoDxthq0sJdIZa7iuf+/9zJoJGilzm/dqw3nQDKKBZaJOoR/I8yROD+1dg9jtegcKv
ZAsC9A4IuUvo1lPsxB2lJ/y+5rcLKwZDlTL7cRnxkMejeQI9vqIXylo9oNwdsGa6zMjVRoYiFz+v
LieDg+2OTi8HpbW1p8zEj9zDiIP/D6qd7adDpO1AcuXDM6KZcg0R3VgLe7+P0W8ZEzTttTEgpdgg
OO109C9mtMlj2Gc1PytGc26YJPrPGiV3DkekaSBnudZWy+7kb96wvh/OK5R5sqgNpFMnwwDJh+bu
8h8vkDmW0Jcp5BtxCK50K+yfDFA9Tp9bGEG+2JiqjYsAyjTj6Hb/lFHfxAdBbWBnG28hKweOJm02
JdjHsd1QC7zKgrINtW6CdSw34U0ExMYDgm4VejStgLnWi4AGi1kDa98A5ONWlvdT5ceo3/Ep/Q3g
qsPFUcGqHE0qGMuSyANpsZeS8fR/GY3Tg8XanzuW8Vr+6Kmm22WPQdV2/0hEV9q3/4U1nEpxW5CX
VXg1mfQ9VMZoaf8OJ1JT1XqeR3XLzCRYzVUkEuErTn9h1sfPzX5laAmL7cAg3Pg+6zZs5r0yXHnv
zyOGIJKP+Bldl9qxKziSQNJe1BM6QISyGjSITsIchj7K4T0fpYo5Oc7s6mPYSN800KW/L8uwAnLa
Cdr04HdsDEkIkf9Prq3YbhhjprgVtsdS6KFgWoHrPFxZ1XOBLKopBelhXx7XgtJq+6AoU9v/CLOz
X7002LzGXoT5UApKkk9m1MR8l4R3aZWyxs71yZqI7nDy78AddtSBh5dLyy8QTqxzephogK6GjfDr
kqUfWgnY8OnhNwjMQqlziPl1YRI8EF1xWWQP/GydHwTHURupog+cRUSATw3ENAR2n8erOxsOFPRk
Ya0BZgCSWNQLrpR5SyA4gPy+AGWfD40pcPg0YPohvXwk5Xj0XUnfFiXC/2rHri2Fh5SBNJ5//Q0/
8CW+3tk5++jbTf4rH29mwl8WFlQ8I7G/dwOWoub6cOHPuCa5JKyPVC/9OMjFamo0YjUWhyw5bkP/
qCcSTfzIUWe2vBGUprlNc5svgYuha+cyyikw5YGbqRjHpcj8nzw4aWs6ekpbW43GWBfYOYF/A4nD
9O3XHn4kH27I7C6ztDQfJlt52voR4pCK3pXLM4HyIlhwiTta2MM4xxEw+bzCH/srysw9BD7L5BSt
48TMmxQMvBgcDb+pZTG8o8p1yS+amKl5y3w8K6lpQNo5DQcIYDlSyfHfwJ8YDrCm8mSCbjkIkStg
GLuhdm99oj6ZmRxI9duAe9fJgNy1yKzfMf7F72TtSCW6HgCE1qoJqgSeepg63LlcwziMKRVI4ikU
FV4gT6RhOb0PY2uzsl0fAddZ6di/1O5Lt1sLzbJbD1/pOMyGeyKwOoOMyXg5J7PED4booVez1KTs
7BEoFTu0pdb/qjKQPt0Y6v3cGN3nKssMMPPT03qdjbmeVi0lUqlIXCbxhW0a1l6ffN2jYFyeIJSo
GpCWzD8k5nFE4xTFQ8XPEpaH385hY5SRcaN9Xlnm+kVKERuNiQRPuKmx6Zs0KN3YypYA3HOsWb3Z
/9GgrDtJ3/Ci9jVSuOk+GxLmvLK5rBbgOG4SsU+/BadPvaVd/RuWyXFkR+y9QiDnp51nwxEp43u/
5xi5IK0MOJCI9+b7BPmshfqMqWhxmeQbXm9Ts/ZLazNCZqueEhbCB11AUPsckYE1Enhv+GTL938i
+zr+7lSAmXeN5mcJjqbnEVPIf96F8FgaU4kxfNu/Ol+YoQYfgrna5WpPHRESfYXVmy+ik0ma8BQP
ZpetzwLidsVRBiUWmlqDP0/Lzqu3AHCKtX/VMieLuWun0cfx5eNyTTr9CG/vyOtxIIJIddGKfMac
JHlrODV6CJjmfyC23jgHuQTef4oRH3FhWM39Y8M+Wl0N9MQIsly7FHXoLucuWNGxWdXhJdKW8jRF
bk1wBkizE9U+jKtf4SwO5V+XS5GC0pjA6zP7HwQqLpUh4H1d8V3DT+SsRNhBtpt7F6kt3yQ1564H
nxzoUQTPkgOU9TWBoIo/yD4ag+7IPQGofx66nKP26glml/eLpOEUlcHIexZ7e7uvKKBGb5kRmu/8
+1KFB6GaRimk97U5P6kyEVHW4C2eGn9UTq/Xf3OJLsfYSOME7tQ1h2LKu8t2n0el+1ANAjtYwMuN
nq/VssqBuAGvpRPn2mRCQcDQy0wX4zgU8GEl9gg5hijVFnG/0nXjouaTsApktmhGvvm4HJkdcA9n
MZFISFpO0WdD0aVKD8+rGxM7WPs+7W9lMT3ib7SXOomreTGpjR3IFOWvCwd0cdXb87ZnOaQm1cKH
zYNl4yHIo1r/As+d/7jIyGQxt9NTV9ydWRlruhQ3LO6Nh3iPQa3YlLwLpGPtDIe7wfFYS1jGuo2i
S3z+3U6nHf2/ROHKW8YPHA0B7POYNTf7rjUzQIu+xf2nH8QTUvss+J+DbZsPDmWXGOts8XovxC4W
trMq4q+kra0BL4HebkWzM8bB+RWbJUktSK9S7+eqFK4Gk+D7uH4T2IzY0tb9XspfxKSui4OctSa2
ZVSY+k6UdYAUL0nunZDxJBoJqjmWjc3km8YgSv1xR0iY90BNJswD4QBRUPClIMjRA/KOdA/69wrA
Wno3hH8uk0IOaYDqJz6sETZygA1TC+3U/+PCVo1x+NgCKDuNBrp6CNW57N5rtW/Hhf2AR/CK8o6q
GTNkhGApDi+gdFBU4djW0fGgmZf/iQyNt5sk0m5MhnwNduplmFo2u+Lfr0511NfWWTBBU6kYq+2l
dInxYHWHz4z/IOxrFZQuFAoYp1318V00LWcwz1OfNQLT7GBpcrtxQKZ5zF5DFZCs6gGhnr5zEAsk
5qv1eocB8lMzyyaC3rWXUclP+jmX+1Zd7Wip6nlmtAwU8YbVixKxai+GAHBKqRTNNFUvK0rdYVJV
Pq92qIYFwT1T0SD8zA5SrHdWch6LM10DibfrBhzcyDL0ODSeEl+mhsK1si8BKuwWifANp21S+g4D
5Akf0tMlycU7SDdREuZtzvKNvJb03Hi9F/0fJ/yJSRCLtR3BZmiQisnRZjlXhtH+U4T6lSFC0IuK
d6zMrEzcZjXCvF9SixftIm7SxTuTf0hNhlSW5v20P4oFxJFHv8kNjOHtajjytHAIdmnD5Y2pkIBx
GdOymIndJJ1b+JGOa/PtpBc0v35dJVHZi73KtUdgk36Zt2Tlr8BCxevtLd8tSnOSbfqWmgWB46qo
UJO7t93+B7Jyt1K5qhzYbhEVRkBF2cYqHP7FS6+xFEXR6OMpJNbELHeIZPS0RQOTnTdwxhHQ/hPJ
3HkCXlClt+ym5otuqjfIe7hQZ0x1czaaGQTiDHP72xdPnM5170yNIuQOmFHp6gzGMU545U4MNqRV
kFn9K+BggRihVbi4qCfTs0bD3N2fZw5vm0gqt/OfbVGqH0xVBfjpLOXfJp7eW+NAQaMCvDlA5Ao9
4cxsesiFDQZtqVnnDQwT+bXd8VOC6ItkYeOORM/RWurO7HAi0c4G2+BBaTVD5KjqQwl/91yxoKXu
W6aSYe9Goqb6v+srSFQFImbnlA7ZhFfU0QKzXTJSDwrkm3T4ktHW7uXdDgf4TQuH/RqiK5FdseTM
ygc3qWVEV95vdzm8eYAIunaohWYxlEI9+6+GEKumGldh2dr+SYzaDPtxWLoj172ZNDyIq1mh0+QZ
6QGGIDGcoBAtZQVBw+mkf6C50eHjgCjDLBnnVHQSqPHvCtK4DPC4TwJX/ZWDSop4h75xl92KIeRT
XX4H1ZK7BXpyeX2eYymRBqJ6j3ic1LkdNvDR6i9euD61kVA3ccWXG8RKsSwf1Y0ZxYIsFvhW3O7n
aTkU81OfxtCubCGzOY/Fu0gCrmSl2L38BGM9SnHNZC9uTv/grE/PkfLJ3Ea8dpPQJ6+6zolmNb6n
bt4Zqn9YddjTE7YuCYofSYfiVUmMRZZrI+urT+nVh5sLoryCROkPOgorWZz8BnG3vPbXwoUgojCw
0Z5kutL5kZuSXIgqJbd9jL7bDmjHlDODqS81R7K1adfNPYjeq/srDcW6/6JXodOuHgvKB8ub6kj1
DIuZ4RsWVyQNfr6lN89G87GUXTO3NlO/iIWukl6rwlWZQSdgPLOCMC73ynV+5/7Re474wiFWmhv4
Vtuh12wHKHsS3jn9rgNZMVn6uykpmx3hHQvhw4rmSxMjJJuAacNfe2jQopT6ps67V0tejspzdZle
C0AKtwO9nHFfTuk0OvzTmgIDKs0ut/SdClqAkVwlgif43cZ2N77RRDGcRlJBYWgiAr9kwytZzdP/
4/dBwHzTTs4MEyaFJS7WvzcTkQhyDxcKM22UJMSO+ClHwE0dzHtTXW4rx4HartxtGgZThB1cXylh
/AA4wnYSxT++QV7/0fu+K+O0cevGeO+UIMTL3wGkw8UMwwW07cRYcJGU7evViuYSN27+sTmpqnAz
DQnkPFq/mB1JTZN1rag0jc9a0G+v++ad1xPmQlRO7WHYjLeNpBdBNFa8TI1JhcOF1aFhIVFJvGDZ
AN7yMHfrgTXLxudAhmjFJ824VWVHNWFj1bkvzccV3gLr6sTgAoUyxRRpZND1SkPUQgWXZYhctZj9
TD1cPyWqjwZvZjfrBrIOORir8GJ6JF0dgLhucMv+WGPDkmmbgFDWLadBFQOsEl39jbnj90Uy2J2p
qotsAokuKGTX/oxNc9UwmZgK3iwes+U5mEyUfZw9Ar4YgdyjlUThiHJsmDe3+2Tx3HhtuYH4lrM/
fyhrgZRYx2T1cG93vjRzDALhT7Ay69WfxvI6XqTKovynBMc/Jr5QRUnHccQaQ8z6PzOuQ9GKmuJX
git1sAs1knm3e80UnT93ialWics8lwma3LH9IHJZD4ZO6lUpmFpcC+4FKM6jxrwBmcP3YPgMmfbf
AxhUpz8rfzyMZFVBNGBiCpEeCE+YHVcOYbtq0yTyWS8sDnYH73XHFkssNCjkk+GpQhpiRSy/Zl8V
+8PGAzSWM32f/F1ifwAqfZ4WaaLqHw+YI6e/4Bh6Qc8Voaja9RcZQrLyLnLdKFqXfcG0DA0rgmd6
80zmzL3e9xA1KqdGJFLy0RwSiL7KBNtp28ttBzLLXD5/Cbr0dZGl+EzB0wIBqOrloI95WvLapnB/
xzEYilM723hYNbAUT69PHe8jyeYdDhDXeCoiKbRtXWw/7dF185mxar5YnaB58ipfhJpIj3vKi0m7
IeNSQBl/ZGx+dbB/EqqcLFae2ymMvEJt5xz28d2VCc+guwDjxWn5cmAmQsGRKUHFH/F4LCpUi4q4
/H1M7zNJKnhsq+r3DDr4XgB8aghv6m9OuaaiqgP4TZFni4HgG8peFZ3HnKvRFPJRDIxH0wteb7WW
Y2AXk8qfzMoSr0iWtY6veuWi19SNHAXO4JnJN2gBKH1NUBuBtk5eSJH4W4AiK37efxy3kBczUibb
fxxSJ8F063y+j8ghXlVyszr3lBFj/pUD1Yt4paefhQdxNewqoE4cSY9Wekc+JQrFyeNbeQmwM5f2
SDd+Huyc+B1JkahVXcmevcbSAERZVu+tTTsHqrLHAI/7An3OaM3ttuAHt3cvtz/B+JtoJh97tG9l
fYztzQqHgnOWLVlCv0QTH8RJKl0qzL4UGWUIvVH1sTCCK9IXN4DcHYb0PyqF3qf9YRc4jUfD41wM
5Xf2X3EMlooPmz+NxBrkbCgdXwjBSAgnlbmiBCpBNx3Otd3rZZu3lnaJqAgMo8L5csOVwh3eE61U
Zy8Bts7gvA3ijkjWxVtTEdNQ9TiNJy0i5x3sKeVr5iUXKJAj4hZLhGooRlCvk3kUexS4i1I+m1av
XIJmflc+FxI21ThFvVdhX33bD1Epyky1jgpbrh5m7lA/T2bk1IvMiEuRA576so341Q2KKz9qbd8N
DvyJwseOIciv6Cq1Wstmv6Rl6i9XEt/3mkw9IMpRHU5OxS1FfT5efH+aliS+XInGH9WnsVWGNUlP
yrFQF/nPvJQt+xHltu/CZZ+t3S7Wq5uBWxVF+17XYSQOCWPB83zeGxQdWQ/atPMbf/++c3U1ZyQ+
ZZF8m/eTxdhODpmkaUB67tTOGZ1gbo9z6fHK8aMhd4p0QIlDMvp4DOPRzuSxT9fprG1PHS+pvLjN
K7F3feFUWhYzlsu+Tc6Z4HP0UuopUDRlXrj1owdQAH7af+APmaEMsieOaBVS/BJmAOyIWQCjFfD2
jQs8f32MOoTDvTB41yKdoY3OjTF3MB35+lc3ZCuz97l/mF6z++qjMjB+QV7vGEvWNvDkOVe8HDnE
8vuvqno8xXV0to75M5LUAKMhndMznv0QARUibwAHn3KZb89E3gA2n70u6UZcIRZSoVThdm2jK8uq
gJyWt74DKL9IkWRGd3lT4B3wZskaheJKeZZ3xgnd//fxFmuRmdW18W0RIMmBKlQtCY6qYTX/V7hr
PGs4iYX++HY6kRCTbPHDoJPL7w4gvDkGwwrxNN3F7iQx+gn0sWKuKpzIO5fJJcKmN5sS1n5hr/Nw
SHfYVLMl6+UJqPt6I9j1Iszd7oS5v63yCAB97ndU/eMbQwmRKiuZDE6JzTEM0b+NbDufS4AQKk3X
gX+/O1kZMelwMH8w0YfUERLxOE53jQhS3cY+ksPQ4XHcVZsnMOO9tmcXmFLFe5h9IDqZ4FAvS/cw
DnxLV3VM2tIoQT/W6qqG7KKEP4Cnz+WipaSFc7o2nEdfhz6r5fqCyym+3wRtvGNcmdxamFaZmcBi
qd0VzaoCBPTZ007xXacyKgleaJzt9uWHXuduUpg9eTViab0d3HNTfD0XKWPUC00cIWeZqWFEo47w
pZ3ARKpzdrY1PKf/v82HAol9fq5M6B4ZofwEKDAWL+i6yM581gNV2ngVM7OB7t1jIr36lPmeF6A/
VUy7A18ODM3C2E2Y9ehmSdWD4nr+dk/tK5ewM0whuvEUjmFQPg7x/uKnQ7WRnbTxz8Gs8qP7Mois
ENBu4coe6wtqgtkNT+S6vwu/tbrUcPsW2nxOT39CBKh++qPl6qp20jzKSNMGzAYVmWxbE+7vUUNQ
hFLQNN1WXSXUD2WkRd1Lva/REvnFNIQ1cIJNnOUQoqy567EX9BJoDAE+Rv2grvEFpUuv25WyUiQC
rppIX/tbFl5aT56dRLaPKaPN0Ok4TYurfFytNhW/UDOpTxgSPRCX2OAOl/OJ9j/o5Pb//XBbh6Lh
fMdYvsqpxxQNjK9chGHeP03txkZHZ4gFaocUF5MdmwG/f/+O8yvEmzCi+KT90Rwd6B4RKN21ZL+a
pZ5GxGKDcK8T5tNM9XiyHKDUV+0Br2q4tbX7g97eJMxSh26HauqbY1LS1k/bQWCjkuObSKxpT3OI
98iO+bcIIbvl0p0IcDXZ4UPLzqxpRrxaxSANZHOH6L0s+VC4sUlWbUIxed/tMKG0AEsJ7S1Nbm7E
z8fBlFlV1DUB1DaUdLA6urlrhMHRXTn6wHNqDBwJ4sbgPeM6ugH0XdxmR0tUJc0JzaUWT6Q9d/Wl
Jg4H58MqwrdgPq5MVkjYlbSUC3k08mN+rODbP7rb+ttobfw2dQe1hpjtR2pMHuUVrZq5guShWQMD
p2JFasVKPRgcSKHupvT1l6K3cuVlychAabnrsppt0NCCQTbJxn8qv1Qry+fNvfmr8NBstE3A4VQy
rKGguiNa2LoRMcCpYPtbGM3KV8i+mATCZdGQj8tOEgX4skW8zj4l2G95Q5b393p1dHAv7XdQrIJL
AMDMSf+FZiwRx0hhbHursern3LwHsLZ9f8AA1WQh8N1TMWWLpS/HPuPETvwIsIz5/XEsn+pzzBM4
x90Fag+X/eHEWZD3s6y+m+paPiuWH/vMf01hUPajH8HEP3V2T+k0Wb54wGqiix5eSQNCNzDgUGDj
zgh9RUzgQiNIY7TGRZyqC0w1dYA1d4pJ+d4/a9p+YbefFtQMoy5jm6SOgrByALRQqwKJA2Mie9ZC
LUpvd02cXNwPZAFfJJtbia6nhqWjjKOBW9aFO2/9luDbFqcHDT4REyEjX3axNBYYhYmToH3+HNFK
mnplJAYw7v/aM+/4lIaSKHHmwbeAaK/xPLyalfe7NyCNx9xm0yE/3AWJNZ5NRx+TPfQ7D1MWK9L/
KRJKnMDTg079PNuOaR5xY8lkPObJhsvpKiNsswyPJsqei2AOxgNZJke5I1GWRlrJRxI5udvPnFpP
KeJIsCyzI7nzZIwYj4kS1xAaLxE0KeVDA07KUgXRbnj+yeWmLTHdrMWZXW4sjywAHY5f2thY6KvF
ir7SfEqoawrgkUXAIinHJXUozU06HO11S2oU6TPU4+KGBeAyeeJMF9qRHXshoFZBM/XddGjH+BoP
Dax7U5U3KECDNcBO+eUF/dMRfuSE8b4HjX5Ku3EQbagvzAKj0HvPsoewqdeN2WWtDwmxHFBSGK+w
Q1oFq7q5ciWcHnuR12MXjpdQAhMr6CpuGYe++edfGycPQMyRxJSwts/YhVrtQq91L3N3KzpzEBcr
V2f2AEdVAac6W4dGpZVH5g8+Qw8lbXj/OCIFUWkMpGIP+YNGcVDk0sDE9nTfikeMuf7y7j80x+f5
2C34u+xmv519eEhQSU37cbH22PAJd+CsE/z0qI+bJmJtlNPVnlcJ0TkrYml1C68RC4L2CuidVH4f
6Jmri0UsTfiGywvJbQxU0wgcjQ6ZQLL+UV4g0TxEVtjaANcKAavUpUGhetWrYhe6qLVea+34EXUg
gRt5ACSrjv1U+Qkor6EIkpDZU5+/HV84OGbZGDeX5ecYyvWFYTvKdey+NL7gtho33Pk66MRzV6me
mNjG73nTbe9UJuWGibaHQJcViuRb7Y1N9Vzv3Rm33gPOM9mToZNpay83/bU8UfyRumCQJzFfIwrM
23CYvcJYK9BY3Vn8/kwJFFSs5mjPXncUNjxZqQh19y3eQWuK/Y9njEUVT/5y+ivoBRpZTL+lF4OD
ZlVWklFEe7JgQDHHtBmQ0Xi9wsvu6hlQheVCvcHq95GSgO70hZ4jniya1d5Ni69NXnV4pSnz3EAL
vLIhxmJfLdBveBKQTrf/lPi7Ws4UnyLx+W3rzlOplyCX5Jhd1w4nYmhjfF0s03KhBLGgi0Bg8Kcp
3ZbqHBoiJ2rtJriTNhC9XATnipKAOpa7qtKv++Bu/MfRXFihr86a7xpQec3HM3s4ZpDrFhBCeKMm
g1G1ND24DqdhBF3VHWhY3U82JQ3Dg5Z6IWy3oZK0sxl/yqR/qyjf6iiS0391hERnBPrxipH8vZRC
t1K6RhoWHhkSERpKfQupOZ5ySp9DR1BCYRowQONdmNdf/4gq32iYoTah2MbBPHtquw1m2b/zFQyV
HjL5yl+BV5epmPmwwD4Iqi142HWa+/292ulJg5eQb/U0SZk41sjMuxthf00Tbn/uuArWcvs28AQO
ipfqFQUnKX4d14jos4n92VjzITVnbQJAzvBrepxG+5UuC31CmfGv0VPN1DlyQZX1flqgqEjNtcZ8
tbynPEKBMRHIb4iKdJg2mz5dmc6sOIIEeCH5n8NOvAWK1rwZ7+ijyUNYCdioXNTS5p1TJcV5Ap9w
SeWwDOXZAcl1BADuE0PEH4ebxvgNMEYkOBtDzQkZEdJqXpKEOMkwYp9iT2bzkShjCs7FeUQhDbaC
QAFkQJXT8nR0zZ9RxpRFWvFhUCsqRxXHIuMIOFEL2LvnXWZtusu3FIp5d9yTckPU9zGvyaQJSiD0
jOVSV0fm4RyFfzvZDvNKuXD1ifUjYnAmhIhEdJparna/9lSUDPNww8gv8qpIBXfVBvg4vUHu23xB
//HSkCoyIuO2/vAijsxIEdsi1ouqMCBCjBmZv9GG43dPJ73laeDoPxZde5+Y74hmVe+zpjFl7myW
bM96Rdhu5j42R465DEU70MgaCjAgr1FbrV146fOKAbK5rsZZlVFws7qZicMX0065x9R39P62Ic7J
NgoAO+ulA/kEaQmzW+aous+rCF3Jg7qVI2wW85CPyqfKodltFcvqLdhRfkwnxtHoGF/YdqL9b+Og
P305ywVY8R8N+l5GT0HdfnpmuF3yxLKRVolyeSZqqy2HRPupCT7btASJMD9cKQtb+Xpll3km8w1O
OlA2cgaoEPGvuhLMiHNV3CTFtTOM+txQYc2La2gtgCOSYnwXnilQyx8seUJPd9W0rDRcVE5HliJJ
6UsOhWkTk60rZC2tVcrsby2fPFytusz08KqpRV96F33fkTQf1vmufYPnSfsdKylEoIHMp0TnUyOJ
hyBIwhV2iro8y3qxt7Amhw9znczFbJ5kzpIH1T/0zrnPdHcJkroCitMhL/MnW6sx7i9oekeSoTBO
yUU9ddeqgKI3HGq4tSEWvqroAIQ+mPxGBqxpW//UMlLiQQJi3bUqM7u2alS1x0MPVjRintIyGPPv
MPTv/H9eRKc0VqBbrZyehRiLUy26tT/rygvbGPJfOuuZNLn3iYP/3jMP8GTnzzqRYKeY/4lQLoWv
0aMeGu2PY64Q1MhaZdrqVhW7h3x54pPQHwTQKL52P72Xtoqj7H0sSsseLxI5CiD5VcfrLuNs/r6c
enrClN30ZkjLrFAyJqXY1P8mkZ2DUSVz8WFs5f+y//AKwunGZ0xmZj26/50b4jYmyeH+YwoyzMx4
QMBgMpcujO/UEDIw2d0PoZ/E7hOK0Cxi/W+vgWdaf5MGkEjQag/MXXqkejVPv+sDgUadDVq+WJ/j
Yy+bgw7lDvOwyJYQXErliUgyMvIPoV/FDO92q/uesgfXCE7o0Yw3i/U1Jre7LU2jAFueeUXLZt/G
HLAoAyO6n6wxk0u4HNkIBKDjV3VjYHehKoAt368SQJAsH99EuOFtthrx9vvyBkTdfcF94raL11zp
gU60v6M70X0CkQg6RUxyBjuDQIe3JJ7OI/j5RT3rcgH9ZKaME0A31OuzUE4s4jxqMrooYsIrmo2L
sSDIcUJdQtqNrQHNp1++sjzeVoXWqvmVE4DE7Xv1tYH21MQNgxNrenY427EsMNR0d25FAgso+XC7
c/MB3qVWNjbHkJjYAQEf0xeD/3MuLF/PnIc/fYVPDZfOz4F6K6fn+TGAPAJzlfFasi4MaCyTiEia
BwiaBOMJJDqCZD1KRyac3Bnj4r31Fn1/y45UeIDZMZWsM+IjK+HWtvUpJKJ5erPHifAs5smt5A2F
xdFRXk9csX/oNNuCtnyaMsYWqcfRyNWZW+ayUky4Tl+qZOlz8cry9ASpbIn5vll7pZgudulP4iPZ
heruaoboMjgqgLEs7e+kMp/AJKJKqCq97y+oZ5lNAlt7v9L70Cqat93LxjLQK1ENU3L1kZ2523ku
HrRy7RG8u8efybEDfJOFusR1tzkRc64qhfMieyMJ5YZSm2RzCB3kz0+mJk34fGKpWyqZkaG0uRUi
4EzTSk4tpyZR3gG2QUFXDd5cJWdZ5MCXjrW1LnEreTLAPN18aWfND+ruaJJb/SFwc8bL7i30L0UO
x1aLRIAkrUAwkH7SYfL6DETZsxN0jw9d/3gSYYBcWJPxNGIDJUyAkyH9y3y52idLCfsrsgNYHJ85
mnBUd1HUSVBnw+Fdk/ajw2dwlgP32xD3+w4FmbIoMpZSP8ngEcG/vP5brGGqNo6XVz/GI1jd+PDX
VvdGM3BhR4AL+EAHbLEgIYuVu0FDw1podzxX5IerB5QCrM6zzxSDzmwieSxqqRW9N7APnsf6qgU5
lJhA85PaN1VJsQF6SmDTCDLUxlvVeoGTndaH3g88qDl0ZTJd1pUb7t3MDmtlz/vQIhYhFUUTjBdD
XuYUsjnwaVU9PJc8hXwyGCCp2ukUca3RXxzjBSLtH/7ONDwaiS80wbg0Gw06fflLrBAWruP0I7d/
UpC80LOZxiB5q2frITEdL7KjdnzjbAIVn5hwhx17AyF2yLdz+5AGhTbjCejTDW8vdOxXqjAHgxc1
gHleCHPISeFWWq88VIjrpOeO1apyssMycKgdz6sOIFXzJdND7Q9g6e1vOgKeF9ozhmt4PKRuYXfd
jO6y5PnN4hw/aKy40kK+pmgE55QMBB0SZCBDp4fvbG5uOtJ/yiABa00AvxAECmRtRWodS5JNRYrr
1VuTz6zQGj32QuSoInokge/BV3SiEWRW6XQlAlBChKW2a0Q2u0lA2VUF7Z02SVJvX0KLGLtbEsxI
XHzG2mtO2rIjwph6WTMF+LQ/e4uxyWYVSrjq4ZU5nHwxOfq6RU/VuXwuYGfTFOxjmZr5X9bGPOa4
NmvEO1lpZUxwavTVyvLApd51CFnVhA3mRbiBvZqltUz2CuSpL+asrGkzg0/WaianxY5fLr2Na4Rb
eJslyhG4LWmVIKJMDpCTWWMg8WEuaDapWPMCrquth9TkaCD/YtBsV5ujoJf8p731JxC4TbmpKtkq
/WnZGwYpMMTQbfs1gJa6Ip4XXeclhR5RUDBj87I5pvV65zA4kBGJcXFxIhp2dTYDmua47pFxNN+N
sUnPHMX6TwyP8b8YxqUmHDPhGJecp49mywFci/qBSBt8xbXtjoCEKdsduufIt53t50SwBBsLriOn
kHPZrlx4HK+lic3/IO8NKDR3G1FS0ip3AJh9WztYbD5gjq3Ov4BPM/Poi7L11wDLlD7c0PDrKL7d
bun49beI0VrfTTV4qyn7WWwrE7ENw+UpRWYeCYJq4V2ZeBoXzeRxETIhKgoOckHFYeQnP6EKVHNj
3Ahg5GJ8njXrcAxUof2ko7x+hcdtdQ7p8G9bLFmZhjYAM+JZjvLNqlLW8CEO0nnsr2VJ74YDdqRQ
e6V1kNGab0dP8+jRe7HnU9ik+NkQGBcOV9dTKl52XFQQIB3AlEeYKcWb/Zhv9NpgGFWps+t4aVpU
3CguM5y+awUlJc+RCwLoPe08BNA7uQrv7meaRZGbm3gIdTZpKQjl6go6dLTFwwswGiigzXZ+lYQW
L3JQzdqfe523kWVFQ25/ikgqxaw2HsEyGqcPg5pxTi2I6fGgIg0k2CtnDdYl7ofxTTm1JScisAqo
xj5h/gwCq1QG1jLjfJYQI0dB8Py5/6deggfhsj8Bq7HWiAlir/3UnDF36Y4HHzYbdkm5Z3u0eWuv
GErgoesX21XgsXUAZGzRQot/Mk3dE9v+hsVgRk+lKwbdxZ38JoTCZFkkcBBKU4Ko57a5sXXxo6O/
bzS0+7p0p71wj+1tzXSyYOnH8Cdj9Q3QJMbIuBduRL2BV8oXl1T2bSwoZRnp+EqXMCvdxfh3iVkb
qHscjq+2B3f2T52aXIFSVLQgNKNh2zFUCHqO1g1ro9TaBuQA1Ce7S/pv5O+xfAr2lr2Z3jqaox+f
9Q6/vVMUPfsVBEL66kXYd6QNA3kDQC227argalEDHVnXVOTZOEU6666UDkW8iB0W3T9d+jfBV4aZ
kSleWaPdhaAF+gddBKQzQaZDKR/5oi8/ppW+wdMUELRIVNd6AO+VtV+Hc20LrhMb7TGhaLT3fvkd
+FPxOr4FRTVm3EDEL+qzGsiiafG/FNWDaIEWPusJ8gRh/loIPH4fa2WMrogPPIzzXmA5mEp1mu+Q
zyOCtQP9GXTydjgtnUaf4L9BDnMTUVMjc/RYlIg2HuzlDoGYIr0N0KEsUbEQFkRWqLyAah/rPQmg
ASq+KpJ+Rekhfg9m3YCN8f9XPPPToGezTgJdzINrpWUBOBqu90WP+fz7/hrA12HgZJD1xC2LbqBX
4DvZMx3Wy97t+pVAF4zqxjGOWQEhA2aV1kPStilfyz9XZMfmAVPaQWaMaobFG+nLYGvjH/gnOg76
vfoszrhG3tfUuDPiR1MlwFhaXvi89IfGAXQsAIxlKZgh8NEeJbx5lnkeRcYQLi3t9KurL7KQCqaw
VD1d6m0NoPkHdyFqa+kTLHt/TqXkI9Pcil+mQtyRfQ07YTf04eRSBs8AenGtqgIqhDQUChJsT7DK
QtTYOOcFxHx1P5GrsN08AX5RcY1aOK+PV3YRTc30pIYUxSbQlql57GFYD2XyfFCK8r201lgq+xl/
anoXVkNBjF94M4a5in4EUfL+yJnys9Ur7p86qScreYFgc1qdEbU3ahM5Dgpd6Im3oouvx3JU7CKD
TPaPkGK3nI+SekUPJTYTzNa8fSDJNky8XK8m+ET1YEIEg50SRWOjzICGv3ivDqAqhSGidYWjH1yA
OWMWEn1jelqEDvaghWBNMbthT8UvYqneYdfFkty9J0Gyzu9aFENGQrg6Y+DT6//nhrPSL1XQLfQS
w1Md3whSG5is4sGOm640pjCaQEeHp8VASPgzeGO6FyJIdZabcKPtj5/OcGpbCYI95XYANBgEPgzm
Vo5ndnb0r+xFAAjSgEr02Dq0pkWJyiYRBh3xzXvJebUXukwPmpWlonRGX0tAWuKgDo7SdC95jpU8
eaYWwYb3drdhgntunrsBvJq3AmMnaY5ClEnUs2ud8l2m6Bp4Jgx5On6lbQj+0L4q0SMOSuIs3z83
9wAG77LvU/Ch0S7NSvdPQFGcxLhDz0ZWtPRH6TC4lJqKIH+R4zehf/Qjfyulhhw+5FzqqMUS+lru
J2FgDG6CRwdTcqB6Bdh3SdgNgKru9LjsYa6UWEjHkREsf5QYRF9gdfj8GhKUsGkzZMKAp/eo6/IH
TDlZvvhNV9zgaQSEuqMNc9UJSHx49JnUO7C4LRgG6AUV2812SYwKThP4zkHuycCmcY6ed8rIDhh5
JGhe76C1Ge/IsWi0bh8AY94WEYH5Li1UN6tawuyMQeGgdKw0ihxAcaJlzeRBk9uAipV79VJvCf0g
ADExBcUhE+47w4kt1gBlO9BrdTv9coisGefEbj+MboT8gxs1u6Yf1WAAtRdpShMhd1bumrZVEbSJ
vSBln2En3aOynj6m/DnSQZ4g+38ur2HMgy5FKWe3qZcZ+jQaPLEibp24vg87/HimHWel4xup7SIy
UvYSrug/86Qbl2WaYO8QVijG7Pt5mZw8i6zUSDKTClPMfcy2LMdBA2owswuVDKr68hMGQlU+4s9e
BEFapYFJ23e2y9fVscYKeWM51A4onNPTBRrni/S45AJ+rmGWdPMAGSKq8QfHeGrqyd069/4FYBDT
fa7RTWUkmJWTJ1dOfgAdn2wBgCtd6tDxo+jngOZlHfnvynN4nw4bcUZ+FJUK3u/gJheyJ+ENUXQ6
pXBXlGk4i03qukfKw4Nbk6SYuWeMtCDDfSSm9dKQs2b6fA0/n7nJQ3LklbCpdbjpXA1r4oAzc8RQ
p922QWZfr1CscHTv7YWd9gpVaLy6iDDE4wDvo9DJbVl0a94IEOsvlSoUOI5zyHkXSigbFMi4vHWB
hVz+m+NOtLSBCr1Twxw2zcVT0CiVoFUWSxMcQUWYCEjc3DREoq8oswbUIGbm7obcFV46pGhY7rFV
oGl3cj8M4p5NngShJ/cvhM913rrj/sqt1x/vXsMZwTId4t5ZyjuRZDB4HtfUAHMbL4Eqi3PBxgWp
O2XIyyg/rdXKq+Y1TPhR22tA6Nut0SImMPlqQ2tLohz+W0nv+hhdiIo5+B0iQnLb3k6I2pm7QcNa
Mk390Tqh4wN0A6+EAmVDllapxPiuC1dDK2sdL9K39mblhxBzu8WM78UHe5rNVna17zbkKo8KO+jZ
AnG42P0ys8WbFudkbK7ijQhj2Y/yqi85cuNiLIj6IjBmSpXRinP4Nu//Azgjm6OfNkQPzMeV/YGc
z/SuGane39/D2JUPFEpaBm1FVcBFxJFqix6isIIbfgUW0GRqwTuRulycMJaa8doYdEjssckXVT4j
3w7/Cf9rIBHXDe1tl7IMCWwaFczIxMDX9LehVAloebNSQwluLm/P5SyVLpQMKkAZkP7gxHImlMMx
18T65Gj1yuh34AY1YDTPdZYfRcuEyPxH844p/cLOqu9UeJekgcfqNoKPT+B0P6iVDwJJsWFvn0SB
mJ4FigDnqUZauyQEiIkiZinFJsiZqBbXxvJq1q9RoEb+q5KQTyDUGkEBbClQgD9m2NJJz5wv2I31
phLwJBvrihgy5/vajGIvKaV/95K6aRPtjJjHhmsrSKKXyyKZIO2e7kGTYwIHLWXTGIeU8iV/p0FB
1t+HTC5nUZmk2XH/N/NcKWOKCwBcMwDKje6EanUzzI+YhFLyEPgeG76DEyyDaVUXFjJjxksmUI7a
JrfRMuUw+0ZH1Wp7172CcFpxv2VaEpHKiy9erVuJagHlPVkGTLAW2Vw45CbyMaIDAmjZLyYPNxtg
aF3cJAJ+hRKzroLQTnpS0VEx4XTG9NjPsOoJSj3vC1rxULQlj13x2Ntzx4rON4ubB3yxwKmw3aQC
vYya8uFlpvherWIcQRXQgzR2J34fDUVp7KPfLAjvcjdw5uSVZMRZTnuTr98Vpp4qzBeHAKw/kgbK
782m2T+FV+/88InlkAevz6LPdQCr1qUDDP95ra3DtOWPPEU9C8eHB328nL4uZGcYGNie8V9aTTW7
zghHpA6HJbMNqnxZtG3wu0jTcOT92AhjTTCTR/lsuXhQAeaSBbMh/g3I+HyexSe9Z2pmS7IQI88s
1uc1Pfb+LlUzDLDH968rj4F7v5PwYsi+zF5OM6DPZBTA95DNByImlI8+zqAxjoINlg50obmFBgBB
XWGZ2kXBidyKeJynmkDoFe5aiAARgwqHxf/0L+MNRC/xiMqS0zc+h/R4zlzXzXqmOke+MAqk+0BN
h1XUcuOAl3zzQ+YQc2LyGKBCknnO/WacNwppcK3MjDiroMBeUkdPL+TL/nnZ5ds/iujk2aA9tHr3
zjH8GGc+waCYXHEI1iqgQes0Ui/O8HjJb4q3JvTznW5enh36LmQPoQLfqVdc9JS53iftZ1QLWGmU
tIqvUWn0R5NGZ6+Ud76X485VRFl0mmCue2XQlyRRTxOvirm5ld9hqm4aIIPeOeDf/jPAxg3qqO8J
l9MWTTnQblvvbMO0gZ2ABqP+2V8ZnSCegItOjfjqdTZpzoyd2YHP4sDDkt6djwaInuaW157pIQIQ
VN7dEwYXczcZXaavmmOvqD/Uxkl7E7AMvpxU35xltiD6OZQCe+ThQpBVzesRZL8I8XSr5ihZKLoY
5uDm60eaIFdbhCHSsv2FzBT4p9gHVsFLh6f6+pNlqfsOXB6zKRt9qAyTU4qypuJh3NvgihsDtotR
FDQvurRzWDb7WlD52crQe0l2TsVgIytO683SCs+MNLHraV4v12akQj02XHLVXwMSub99O4zBaX2P
dc7VBTDv2PRHR12QXML9F0sbCUmd46+V02PCy+qYQpNSusdnvt1tA0M3yGHxbf0ptJvT7x5AXf5d
FuYdFHg9Jm9AcbMCyDLOTqYJ4XQ64KhDsOzlWAU4qvxDK3Nkuv+RVeWxnh2drJugAFjAksZKAG0v
7hhW/R3gd7C/BcXikChKsElW3IjtLnoCmnz097xHU5V7oXAnDOk4FOMLA1Hr8YqvzmXKktO6jfT5
n9KTTcfxfS5BbVItkOwAi7p7tiJm9fugm38ljel6K8sl6ZQvbw2hqj0ViSN2BQxgluarb9jhw7Ff
mNAcsobc86e1/z1bMMuKcgJ9kLxgoSYTBPws6BOUkr3+dzLlkIozdmEl82zUgFPHwPWKTM/JDw3a
OItW/8Y8ib0kOZsWYz9WTilUWJZp8Xd9F9GPPMQ1RsplZvg3ETKalkrOBne0bLnwYZ+PEMwt0M+J
pxau4l60JzDSnu9blHSRtVl2RpiYlnoffSnsO7Ml49RSBVem4m3ECgclNtlDmQDB4A3v2H9XbMk8
AJxBl7+l/TNm6dUvhWdy6w+kn1guUO23d6/Z6YBP5rXrxsIfzbsqnBRYZjLDNAXu/Hgt22eKYLUO
FO7hZDSQled0Aql+ekDhIq7kv22MFzuDysNyEH6wh7bH20bUzPcBZqqRdZbajaXM1jsL3tUHz1IM
vowSZdgI3iX09/MGSHDCEgyeAgXWnV/bRMa+WlQV5DwKmas5gxz8LwDGYAkn5pyta4lWKCojqhxJ
MiobT1iEOjcKvQvG6SIkO8zEGNHqXTmYad/lyIiZmXNVeIlSIND3rJbuPyF2OkRZtnWuYaf9WFHP
tlJtzI2nx0thQlhSpLEg3i/4WzTuAo3x9oKBevqDBxxy0Z0JSw5SRLcq8NR+OE2G73GpEh7BHfkk
kGpSp6xsuw4+OScbcnt8LOlyEkOlbFc+fOJ7qmPTGtjOtZgFJxnpPtT/+Xx32tdj7Sdl/+fb8JcQ
u0VEc9KgcVjXgoHN4cogTV0X5ZGdI2eXjpyUZ7jOdLpjR4cwtkTaZW8Y2N3CkeylepzbwfWRxmve
bwjZLhlTIvX38GCZRdsICDZ+fFnr8czKqwdUWEvCnHRgtbJzHBmWKxacqLETpvcT86vgZgZsQwQU
PMHyqC2XkP9O6ChcLJwmS2b6wUJUI1HXYaJxMr98n0wLzeoedq5rTMN/txV6mptBrAgfPNur/mJg
YtDCUfRCxc2AjVkEtyFh5/vc7g+xZqGioYxEUyUj/dU/sqw9me2xvzQAdczMuOMzM7Jb6bHlulMS
rivTqVJMC5YuFFIcT9Ax8L+8mrkecCdmGt33Ya0Z5K899PEW6iq/zFcgD9GUFUKnvGoZutUalkcO
QyW7JJDrnRFgYstjdmUoKYMi91jzk/vVRfwo6mGfBciI9LpMCkTHolD2xFT+kiQphHiWzP0E5js3
yGRT2LW8yKzvDrSlJqZYMf6x6Vzq8WVYQV/ZEUjZCT5+bBm16b3AUlchoQ0C3e+lsaKFwGIvLYxP
gFlF1/iBWrIfHiYJjDFHPtopaNDjulVDcZMHWc6IEIh+1S6Vv/eZY3ZSwJiTUjDOd5J4jrjwcq/u
ogXdstqfaSLETOvMYoB1i9FS36TE1Y3V+a6r3aJ7x5Fu7yKzBBze/YzEhSxIX1cufGGTeKCPdp11
4/4XxxcNvYoOIPwN/jNA8cpMqfYGROSE1Mw0l5Dgo5FlapBYC7L7sdLUPvn3x6yLyrkXrYfspzia
nOFlpcRtDmCz24F+t32iHiRAF4f6NOAxIpWSHF3x58qgKUfrTaWGzcHESd4Xtpe31wlkdETLqZZ6
dTW7qxD7eyAwA/erqjnITpILFPICfxl0gvemD0ilrxjae+DGNhbLRVaNPGJVdUBnS5QvtOW4KLBS
dW9bvvtpvfBvX7wxNQeE+DDvNtaiOcHBUTWB+ykOAwgWd9m+4i2zuaLj9xfjcQUV4XHql26KmTmH
/QXwdValhuc2n+20Kvh8/yolbJRMPdad5IU0B+E6CH9uImL+DhiT1XK6XK81Fqntquim/QULw/DH
3rwPK9dDSb3952KfvDZJ5DusyxCJcHMw0awVM4S7Y799K/I13W2i5LRRNoVQfZMp+dNItiqWhBsN
kMGu2ejiwACqGPDmWywM+uYI7ahcS9p01KufPBMK2CBog7pildyvohaxwQEHZcwepAzB08V4aMCP
yB8seW1BeRVp4zDluE1b4NjxPn5qPqxmssYViOgbFRh3wJxwUiXpR4aCMFj05Fvhbaps5D9Ffsh+
3BfM68sAAjo0/0Q5AOybEbjKMCtrESljpJPBs1Rd7zy5CZKHOoNzscn14Dl/5LmihIK7IB/g2VHj
AvKTvbo1R4HtqmVyZ/Mu/FOVqJ9WMevHmufhUrrhWsBUwEYL/tB3RTVWMdbJA1IOtjULsYQuFyP9
ONTgm9Y2ObWS8HZQZGLfexDBJuu+FY01kD7pPqbXpupyvSzbQ3vo/j6egti2YBhqgs3XrhNtl7W/
jQCaysbcR3hykchb06gOwrYolMyBWY1t6yQlzsWkf2sHdbv+jm/nWnNS2bbI4YkaofvjC8/DLrqx
/WkqmI6ztDkOgcSxMP3Wpa8bah/y5r/szQpArXz+yNVTYc2yIxjUZBLbnx35+x9rPyEq+QZq5Q/F
PH7vWD25ubTvErYxFWc62LSLuvZuXF1Y0tWv2z9GWB5Yx8TXVQtg5UW0arlAhWiVTQN4VmxRXXNV
LFG+00ud+ipDUTOplI5q4NqQDAJ37k3SfHc87mx19twiaVn5o9u1mNsNWch7UwrTIi+sUYmhEiEm
8Pc9H4QW3SClI1L/QCQPiqhmcjJnRaeMQXrjs6Qi44HdHv+1HaNB5BzCzeJVGIxt0J/qhd6FgULe
kTkcfSFo3tHu6A6jfnXsie+jFKuF/Z6LnxwcAU7qsC0qcvSiRqUSN2GrLdNpJqhgshTpT7VKN6Ry
RT/jxmewe4R+A7Q2xYlr/K9KbF/FxefUbD2RCFrETedsOpmAVAMVs1qvvAyoblRBRqwGtHHKautj
u6k1K8tMsbyxgyrtZbSgjkhqi7iHsY44GQQdDSJaqeI7xWp4nV7DOaYzDKJUm4udMcz/4wrZilhP
cAE4w+Dqpr1Y9VFQ5jUDi+wmUKSd3lsfEoD7sfFNYcQgVIJSm2NT8nqoilYO6tiSqH6w7WEHutk6
TwwwNaVisLno7CPmAmFC4enhnpVZY1/ZHZCLXp7Fm9NXQrSlXH7SC56KGqH+o6dkscyB49THk3LX
S2q7s/KkSHVI/fKeJZ0OxHi4G3d6+NxZHjRu0QGM9jZEEAweI6npYkFgDAKDGDL/5ylkPchCz7DT
D7+TLk13DRRS6eNmtjBmSSuzD/oF4Pct3cSb6okHW4LlLxSj0/ZRh+r72kbPsPz9YI6CVurQZsZF
M+Dxr3c1+SdyHfXRSZBNstMwIczTYG/HOBX6fv5IAIsAPeDzFnRl/frgM8yvrBnD5KMtbWn0Z3N5
8mqruSmlpc0299bHImlfA5gLiGshVf6owSpuJ0nqNNGi65rUH8osrKHHeG7PoyHjZ9HOjf5vbS9b
kWFV1FGqeCr7zqozKK4Iu7okyPNhc0m5BcfIrBba1f+BhCXDB9ci8qFxRjAqbcPDuiuod98ynE/Y
VFEzuawt/DToi4eRZHnEd1f8ShpE3pDP+RrcmkCIuChHwpamqN8nQ0Q1zOuqUNi1XkdQ0d6uLEtr
ZR1SqL92w4wjNnqtRTKuBRDfTQbkafybNa5dy4DsVnj/ELCN3k5Q0mu/RPvSC4mvUoNxmrJ+umuW
lcu2Xl3PUWial6QPg4pv0jZ1Bf21xG8vvSL3X0mmpV9pc0onbsxRARlPHfbI6Qhw1MGyBux/TSuH
oujw7R0qwUv4PPDOxRQmCgXFnkg+MMkkSYGyZLk5X38CdCfRjWWQLi8N1maABvURoofAobvBPkzk
1E1L13NX4Z7gA9VQd8qvIYECwT7QgXvWedR9Df/CMPlWWUxiSaxkuvojQvUPLvdH02Z7JP9LLnyj
oZFYP+aFEnCJMqLlziWTHdaus75CmL1qeKaHOHKvW9AtXPtMIrFa1ugD4H31kUnw9HeW8fW7VMJG
R3ewlr8BOWwroBmwo9I1omSXiu2+lwtm4NW8ioE3RnC9mVlZaHUM8FC9xxxtfQjZzQJnoOO9ijbk
KOHgi8VK38kWjcwFGTyuxS3vmvx/zRiIsEAMAeSZW5aUM6ikeP6Cj821cXtMRzRbWcKDiQkyTsAB
kdygfj38jpEpEp4VJEasocfWiQavI/PsXmrxUwaXlXzoP6vwWy8PhAzcbJQpy1FNDnh8H8gbD6VD
TxhN7rWYsHlb+4T65ymUplZplG4vRwU26d9Qz6WOu3yigiM1xUII78cqCV1jA1ODAItmg1Uq3dpL
l6Cmz/bstGFwc5WQlXbVQGxZTIhuQ1VWeDhp4tKTTloUNoEOdLcptCpstJWmE4v96sQm90LHDpMD
Myx8iWmwx4rRa3sXmymzT6Ll0VMWdMt5+aVpQBOEQFpJoe4OZZ5P5yWftBD9aTx0GbQKLFFT/I51
2GDi/cJviAO4uVJtmVRB2Gszt7jRCnsM3kQYVPtHpg+n35TgU+vtpX/3zlFn7U3f0Q5FjXwrtnrK
A/DWsvDAuzs2PvUTz3inQ6cpSJakgLMLdoKKpj5vhzq0Nx8LUjLFMn1MVCQPNEqzz8nOqUpP8Wda
aMbNCmMc6n0T8+y+gbKk2wI1BwBRec8mPKGFUA0B+2x65a0AdW6PhjpHPu3ucs/hACDfLxHNOGUx
gLp7abUbF/DV3SL1HtKXVMzB2mEKlcXLyWBZ88bqUVM/FIzFeEho5eohcTzHV5MALwxKVpwTcCRy
wGCh5OqaoRUxFzSfEhR2XPi/sGDMbz+ZoVHWldyHF4i9zfqp/ZFi8Tr+lVk/z8+F7vKgZ7CmpJV1
/QfIWcEjE8URMROJqwh1b8xMw2fOGLUxSS8mf9XY1XqtzAkH4yu0Eq3YWvOuJ16Vg1jROklilSLJ
C+lB/5cP6bBphAUGKoWaLr17CK2+5quwW2HQz5xaBdbq+XmJBWVmMJzICSNGIsg4os7VSCbjVYHv
n2RseOWlpcQSfw7rV/wS12DrFz5E4yV2MwvJ3qdxoAHAys1EEE6CAq43c+kf/u2ApqRq7ACqzSaC
4Yg1Rz/e1KXfmFQQYb2FY0KFJfy5ThJH3C93pVxKG9DOfAZdx2H6dFtD8YCm/ON6mYL/P0b/yUoG
1q5MvXRJLlr42JQVftiuT4LyvX4a8Mk9t5XhFxfvcfFN/dmvkO/ywMsLZJ5Znd11vyAcmI4jzi3U
tb375xc5rdrCVlIo0Sr7HjdsofMbZFVtF8/juv/O3WzNf6J5wTt8wIfCtAwp/4ZGIYf/Qyiirbgq
x/KT6iViVrBB0NhJiyxEAF4Ud6xlIVmcqdNStEkClNmX7l0iUoAMgTZPxKsjOCbBHozPmmIox/Of
o77xEQJX2YPpVOP78d6fjKvrTbY8+gdgW+Hrlitz/vU65A8Unw5boDTtNLbPkZqGeU6ZXCL2b8Db
noY4SQvOSWZ/Mu+f2usyPH0DhyxQsbCS3wikM3BkARZV73+PTh84/WISD2sNf2iYu5KYxyhkV8IF
saAGFM7LQfgEaz7qtavYGRk1k8TooVOHiT9kNokJvamZw9hqMKVGBIi6DdNMXo4crFeNhVAxWhB6
8Kd2bZxS9XykpTQrVQTa0Y4MJava4H0zhLvGCmcBMX3WREZS0tIgwfwDnsm6NFgMJgpUdng76nkY
vrijjCv6y0SCbjjZmrWGj6URMdMUbfQl442FYPTFzuNxe/7qibTUZyeRoG+ZeteLxBXLoL6cw/wH
NfjWWIvFvrUMAuqaVnMkUwPU7SSa4Pc2WKtQaCYRZJmVMnOSy58SF9r63Ry8OY+Aixj7n0c80vOE
CK7Z8bUeH9fAeqaNKsVL/L8mwqdMcmsh2Os4usjJjTkKVt7SlQf9k+etGWIxOpJBLuYUlj8/kUfy
ShzQv7UMWxn8x/g5WAoDAn6CoSshnZyPRh616AFvxmnZq7nbu1p+7vm+W7vouFBW+m9UpCAfgU20
2uuksyZsR46Yi97ccqPtWpFgNsnQjFD4OWRX6UNekNLDPxFOQY7eNeno5Wb/h/L5RBU/r/GVBCOI
VyXlpaDcCkmDyYNjCt2Un3OZtei2oDPl3MaVHO4M+F5nS2piu6cplpzYsoZRNujl2k9cIz+75Q9O
2oWuG/DUGi0oL6NlZ2Z7B4OnMUNj653IigpdyHXLJAzawvfEK7H6zj/nf3WIJnFWtxqXMl8yYwuU
Vcnj92RRID3em8CIcqd9do9Qlv3OJExBeZSF8HgQAxBzX6ewTaQ+cne3WcAMR7HR/KzbB+gAgDMn
GGAoaMj1sWLj6as4b/NU5vGLK9A9Yw/FI8SXEVPldTR4/UaFjHjMul4X7sgw1GYKw8wGYVIO5+D4
51fp8GL7FFCddcobTfv5GX5Rn3vuLSD6PjRSU7TcqSVNNCaWQg2UYN1O+LNulHr78SrKXXb+8mG6
5qvosWu1TVOFmmUjC7rqyycL3RkvUpIvEIxsJcI/50ddasoNHjlGleypDqsURe1BnwC36h9LVCb8
OAU8eui811Ah8EQ9NQGy9gaKM7oItmHqac87h0HgUlkWWR0bcCfqu54R+hLhWRmVsdVpTwzIcsOh
WciDNnFEiC9z+kgNWaOtUAozQXX0+Y6roNqA9KFZUEs8xWYXy2taeQuJ0yQScpDs8yI/45kuNoE7
6shZta0toHYQOvcRjKzb52+uJDZg4NgQw/g9Eji/GtSXtWsBfJ9hMfLg9P/+PYy3AoLdVOaFvxPR
w9CkGIInhXjBT3Wn9EBNNFEgkXr3UeofIOztzUY8bSwn0QKf7utmMN+r6XmiY2BgMm3os8Us4kSi
UDo/ZLQdB6Jim3qJGd/8Xy+uykYSvDu60GcTTzINi8vw1vzQck8OMv8Ja8fXnOMeS0q0PbyzBW2Z
K018yvqEa6F0Z4ytAt36LujHqAE3VhRXO/vNjVZ0Ij1eLMdgyri2vDUVktMOERkh4kzwSOvJ8vG0
vp6X5J6LYyKYelt0t68rMD3AiNiO70SUJsdZBgNIYnripdX/DtgLrEoyMTQWbqpQk1KbGBDqWxMd
uCNCiF6D0HJ4VPGO83zs+lhH9+rJ/WkI/YCXgqVpUNPLBPVDt/Mkr77CeRH1LHjHIVD5wwhwaegx
RaaaiOhygrZqUfHHHWtfgwkMgyLGfRBfmfyFaUox8d6mdyCf4b6IFRaAxgkzkPLd1Hb1ueV3I3sZ
AuFos5TCLtC1eMAwqPP19sSuz5s2YjC3il2GnNzApe7BlsNacRentcuYutSBoeEzJMfN9OMQGBy1
byzdERgukYbxxoq9OBjlwDuoOe/saugf6Lgn0yAnYO58VnduNGjZWK9lkNngEKfZl52L+ERbZTm4
4YrCNbUaiJVvlReteIQlsyXwfaJscHHJSf7nncSvsDNnee0H2WlKy1rf5h+CKr0ypJh7rujpvPKX
Jit+PdyE9jQXsAPAifaOaKV/oUd/fpUNxuQ3qAXsULGqY4kysBKRHQmNlqB9lkxZvZJsfvbILZde
tHZBPozs8mQo7WWKVklxntwDYvJfwTae88ykebp0lIsBLE+6AeaE5PGTZxAWrCn6Wqbg2jfIgpC1
boSxw8DyEtmAb8IZdcu8IvC2kT+inkl5yNMWQ/uHNqIysPUY5GrwvarvFqoxACK2okRlE1rxGdoy
wz7pXGEvWvGvJu5X5WWoXoEQxPaPzd+6vYsgXrIxthq2MxsvfXnaegXVY+KZUS7sHR+ir8eV2q0a
cLsq6fO3rs4fYhE7q1kcVK0wVlnmmUrweigrlECUmuP2gqTnrFPTF2A3YV6tMcyiZWCvdqmXDLyL
VrpGj0WDUA0snTaocHepk/NJmtJVpzGaogtG95524DmWZ3eWEXlljh0W2YHVvQop7FQcpKgOFSL4
0K4cAKxl2OTxo5/+nV5FlBik/VvzlNT0FNntwpRk5koDe/B3sG6pnFxDX/66R5b2LCigEYgDE6CA
I0wFbMAYeVZ+wYnDAxC5rQXEOaHHdIE+D4myvD3XMdlAX0qw890rl80ShvCFfFkO3v0lyjIGxaJ/
3PGJCWZHr1fMDBfymu3w3zykeMrFBadtqcPmz9UNm34w0MbRZvYZi+6A7tV4AIAKsT2U5ZCbr8lS
UfHRY9bBsvajIRMSUfJ+5leIJY3tSboqWPuOnRV2HHENfYywggUuQWvEfKtX3DXAUyTzE0ZP1SHV
6Xn17XDPn8CsMtcSvTjey1FZQfJCXoZLAa5XqPGoq5imuqNDDf0SQsApxbLJX2NaHgcF2LF/odrK
dJ7fk/gLnPYOiONFdDhJTy1yDuwxMykqGj2jpxJx3phv7WgqeFuPeEtAZh2FSHXUG/8wtjcbBzza
hK2ocBsc1xWz/IAv584L8Y2r+dERylh1udi8TtN5RwyOeS42kIGdgPD+s0/8EIioKSUFL6SKWy/j
OdDZBTAlX+Go/BGjjMCY+Fc9nIgEcxtOZj/owvn1XY8f0eGDWMEjAOnpXvoNu0KiGoxlwn22+4AW
+zN/knI+Uzp8OiYDzSV6zD/Wn+YIlQwEUgu0wPwN18/HvLjkLRXlzy/i8k+ivoDA0S9xYD5T8CdG
HipWB4Z5xdXzR7n5o4pELO2NlCyKQLoi8vDbPwEKmH8phqTfAA8XX+cgxTqM/ZhxtfJguFSa9ltG
FpP5M+mF6W6LozvVjQR88qp7QWogPNRKMCVB8Xe2CVQ/uDF6Z2ZVDLizlfPpoHug8e7FGUwA8IzK
d+ZjHjf7cnmr1IZOezzRBRl+PkhN9KZ5DVz/X9yHU3uYHHi3dhxjSS4Tg09p/nTjh4ic+txz7CWJ
Br4HnrX0ajtLZ+92bZK95POvxQNEOWLTMjLQPcZvu3p03y02SFkKOSLDMIki/GVHmB774kFN5IK6
dvnvfngK4ViH+KS+Dk+/Kb5wbSaTg3ZHsqOqYi9h3XGxssKGHWA/UNoBpySCgKxHsw1C66DehuaJ
LDEfXHp5GJo+1VLd54O+RP2T6sUb6uDVrrR7fqXLL9kQTsIPo1GOmw7fai/tvh+DY7SLYh3vBxmE
LfVCJ93InoawrBCyA83LbKtRsdOzy4m5K/BRGBxqgZKL9elYNfP2ogbWkOFh1F0dYxAbfYMlpsya
JabdCLhEMNJpTiFFksqJg6kBFRn6S8u/HtyHEwMAPKwvbiodZF2HfFo9TXcaRh+3mZzYlA9lRQD2
Gdem/8aZO6ftK12uDEXcCWXlF8WpdYotei7O4TxuW1tGo+J1zk5nR5QuCQx0oPsNO/jbMOjZuEqR
MYqn/AC8wupsNnW9n3aB0CEvGJ9f6Xl6eFimLxyXLGpjpOwBBxm54AgRAYcj4URZOlGvAxkCfIPa
Xq9jpF152uY+iX5jWRcJkQAARV2IPgvuziuUslcRdZQkiHOiCS8ORtQEbD/5OkXyo87QGz+NYvPZ
sMWmlBIyIuvOaXsjE2PSMqXGIKXtT8P+nKL4hfc9baunQPXaB8bzCdLmOHq1HthCEUlv/24sv4sh
2BBFqV+8Q4lqjotbfo7e+XT1D7OUFSIzg5C/g+xd10hgsd8/AL7PG9juqFLNmwVT26yE32vg+OOk
yA+FoCkzWfqKxebWEJcHdjzV/WQzcnjE7AFvfk3CV4U/c5xBjLe5HPJolCP3sXEN9q7i65Nucz2e
f3rQJtnCA00TA42bsHO6KLGTjAuW8fqa2CnPZyJ1hIAGfFgoA7vVJQ9WMRru1xLFj1zGn+0OymzE
0pjfLY6cCqW0FQFe8b6PwfqFkvGZDTBuF1twtZbPrX1sPOqJ7rV+33UryYBYVVerngR52KZhWaUk
tXq2Z6XjJNRXWav4M85pFt0xMy5XLUTCDvyZJydbOEbKAEJjiATLhvW4dUVHLDsQeIqYxtiaDT2R
V9v7kCXsrAyW1XQY+aJlotk1uuxevOU1BwReplUvWK/A4nTeuS+BJ/qNlPuzLMVur76xPT92lonB
UeV4ITULZR1XwAD89H4NNQV9fN8IULyHG20fo0UO22XwUFo2NKwdO55kEWTY2dK9zWUbll2hvodN
ZB6rOHNKqYSO9H0RlDld3Ph3y3Bm0/IwPt6IetOn3O5135Jtnv0aYNDHdHYo6+9uVBwDyFRnojiY
NT0TwmEN2XkgZzjKSmHnoKMcLKGCI1GvVlrFmkWJpb7gVn+jv+37vnDL3lo9ho5H7l23oBvc2TUe
tXRbBTHtkGzgbtz3/7r85TiahGovluFo3dE+hU6+w0KqSbU3vi3niX1KZx4K/vfHWeFrBuzz2Anf
hoPTEL46At51Z/7GyI6mjP4oF83VDSOJ5MpMUA55GlF5F5VGkD4Y9RAn8NUJUiTvY9UYI1Zxp7cO
ANJfOoZuPffm/KBN13RgYqNsD57c3XNDY/UmGGsbR5fZTxwj93jc4FILuNqyN+OV0tVtpUKwClcP
AHk2/Mm2E9NmW45MWUdiQjcHfaMHnyb5etFSNuQc2/LBJ1/DIrN2BJ3hDxkucA0hOkm8mqwozv+8
oGLQ3fLZm5cIO3cRiyzqQhMOUIT1+y0kdbhHAk9+SoPg/HSpgC3lrZSj8yotXaryHL1aAtgN9qRk
atOiZQecAkKZ0eY/r5jNsq3bMYQpMlKuOUCliXxOitNWFWJdoxhPBBpojRrAz7ouWtcfaWklyIDP
pqEPeFPSpOSraTZfMr5IFRzy2HdR2DCeJnAge0aUs5NvIOawVSb9e94/Qus7W6FfNDn5+Z4MUQ/S
z8Xvxi9QlsNC7WqtVyL4QILsQlY9AKAQ1lpgLkC2yg6mmO5uncHP6TYBY4LXrXGuKIcVH+v2a+Bo
7K9g5w0RfaREkAtmTNbEO0WtmiqjfsMcxP//2ppysTJQKfYxF/0ly9JamMm25NPE3xQxvuGdzfFt
TzYDYsSrkM6V6q9M1sivEok+HR4BVfF9BSUlbY7rkdnVKT/f1Io3MlLS2OImWgYOWGntpswkJr0k
WhaA87KZWhyhULoZA4eKHEc3DPiUNp+S+RLxyyt6kdKJbZI6Pz6q8afSqvK6Hbcx4pQ9geE3ROK/
WNCOJv8zWk9Qv3q4pXBThwu/xkLp55lLQDQeZAeyJrzgUYY0NXcJ0J/KjQSEipZVFdPqzBvv6DNn
xxOxJNODG3wggb6c5moKVdtivsne/tQknaPFJarK75KTNuZTeoiTOWVLI/3MQRT8pyzFzt3svD3e
PDLKlM/tUIzgFF0v4QWjXSQZaCIZuuk3BxURwmknZIqrzaTWJkNQBim62K2lQA9qlRBMvlggId90
DCJrDBS4foDHVlhaSsHzgBNAXURlF/Bj8Va7Eunznx3ev5aZvReJ9MCCzfZ6L23OqLxrUI3Wh4de
wZ+NHMVlJgl0DVv812e1+1uZCE1QreSiSvzASc8nW6jMF0358jN7wkMuxFtNkV0x4r0E24GYmr5u
NcvO9LIkjCB5PGu3anSYIfqe4l5Yhj2iKZRycyzmpCYNPfOxRbVAqFTTje2+8AHXEMoRX1AZNMXc
rH2o0Fm64kzR0+DCCApUms8zD/XOZu6KgSsqoRRl1mJ2x31GYCObfOuSNsQpUHSmN5fGAqM4a6XJ
AHWJ0y5gRBKdLVghkqMYtgXBnyP+4vRBf3fcxvMst+kkAPuFnpP6lLkbgg4CaWIBu1OZk3Pd7/wh
ER73EdzNTFVr5SpuGBZ3Km2wcNDYdf6rGA8Yx5KR2s5+F1cEQzqr+U3Kb6BA3Gq7P47GjnJrGMZ0
FrLvy4D1PMQPxSW1WebFXBHy5qXYP/ppf3hpEXcnd6ol/EPuJ3FFDdw6ecOOBUmUc/v2sFNK8p6v
/if642VVBEDP3bbTAVeK3/C9v7384L+Bb2GAiOGSR3xmnNY+2pgb+CqKTzkOarhogWQBjgap2asY
DIhIYbcZ0+5i7PGyEcJqvq0KT2EIz27P+fjA9HNHv2S2pnne1l4CfYe2jVfQvC8tjE15KfrwIu5l
VnT0UyWc5nVDP3I3PWcwE67zAJxozy9b9ZlaVFRJ+1b6Z2HEgW57k6veTJSG2IoZWrgrgTzaxhzv
vg7n72GUjT37o6Ni7/1jE2Xo5klbCWe8DI8EqwZBXWa+htPGiOHWDMUV7A5XYvoOkDyJsKg9Tn6g
Uax+AlGSNVH6HYNIaGA87/Qowx5tOJAe2lgFcYHYkUtlvHNTcb/kcj7TUNXr5ZPIBK3Mz7q2up/H
MNhlXm8ZgV5IThSSvDnBlLkyn+qThh/HUjKLs17nUnaYgDnXc64YY4F6teW+Ox2N2ULa6/1Y0VLg
Wb0NM0CMPiJFBb4BEpy4/8so7r5N9VJnHPbf4q+FsJnomvlDjxeXEip7g/NVxMycBqoCIEzxX30T
z7fYwBmVRBb6SNOKHDiy7UCqIKFEFPRJ5HZxswNBXJk5IHMPxIUhF/WFlmW8HlWMTUjONCcNbEBm
c1HHGgu0u+hZ8RXOHDEESHHc+E5MZQ98fEts9lHEr/DVuynTR4F6lpJEWCILTJYoeceXr0cgqR14
M2cjcnELaakriB5LnD0YGVQZZd91HhYQA0YMy9Mc1a1PwFu35pTN1zYwexMF0XYnpQLlKEJuXOrV
BRF19Bd+2yPvV0NGCzOGCGN5J0PkEpF/BduzfEf8qFjhdBmOJWLq2DZoW7NE8o5YZYb0DhqQvCQY
xVUsrvf49KJ+EgQHjp30kyOEYI7d+FMO9dQXtO3wGl0DdCptrtAqhhr8gOaIY/IoYyS3aidt1bwx
GdfcrvkbEi5B/aQRCcRM5eI4A+GvOC/DuSQafv5L4hVCzpwjBfhFsGLf9DjWF6nmoeWjTeVl4rOw
osKuPLMUKYzjQ+TcG4R5kwdyqwYkIsqAS0ig31vVSusu0PhEuRCSOMKRkaieYt2jVwCldfWkuD/k
NH12R5qwp3+Tnj+c0q5icm9r8wKKIuo4T9wmYieF6qPDEQa5OIig2B6PrU0keIs/4KcoHmyEZo4+
d8RMWIz5F5o/NfL6Tfpy3mSSduurwTwRYlvcAR1LAV76f7LN/Mnk4VRQfRSCSmDndbEiVnGH+q8Z
YkqA4XSAdAetWEFQdS1XutaeAAW4gb3lL0UwIT5x/F0ylUdpD3wSBmhKSfmH+EJWV7/nksl/nf6c
fVJyuNakAtbZuR+ps+28iknEcyAhcp0tzAQgPkD4wBeOO68vRJNEcfc4fW6cLwAbL7d0b5Oh//e4
yn7ZXdbJ0LtNDq36Z6rdwk4tXAJ2luTZvzkwzUVWVTPSxoM+E5DY2shglz/gKaBpJEodHoO8UmBk
lJhx3dRQme4P8KvhU3B38+eEpcJx6uyPv49JrhPWsFghmudsgH1WHJ1vnI6TIf9NiyyVebvRZwGq
Nniq50yMi697cuUijFahH4VLau9sjLJN5m+yPMVJ+q9uXBOuvbXtOe/cTJABnReKizEQT9PJKoD3
LwC94l0nLniLnxrc37b3OHTYvv93QglYE+yF9n0TzvSCEkGbXl6wWuKjHhXygH9hG7rPQ/+67mFC
vCtMfWU5rHH3BskjW+G/tvkG43pxMKGpDeYW4CJw8dHyAYl+HaXcyx8xeInrr4vkJ4ZK4sDI7RiW
a4wgtcQRk9keX/8D7sIOyI+N4O5x9FZX5yUmQP4yvQNhyPq1dMHK4wjs8bB5sgLkoW3iJ3539daZ
ROlZrVs+XWEEkJvQOPhPw9jaHgXiuRHhko/RdzCqmmNZFyONS7kQ9jjHBhAlvFF1oAmTKiwzPLtM
ETkR81AP4YSRFYPHfLg/I2Lw/PlfFeyR/cRf79Z1tbIiUbv0NvG6Sc3xYY4WVBKmX7JwejYHA0Lv
n054xRRkxUOH8SqyHiOC+DIvHEYgCt9trmp+FLg3VWYw5UAx9iOu5eLUSbblSBqX1KaHUYybhna0
txsDXmq8w9Pi8HGElfuAh0fMYqkf+B//1EmZGWcTLQ6ERXh+c2bjrd77092dRbT7YfjWPwPanFj5
vKsBPRCzIVBBGGTTxi0bJffvXUe82iryraotckNzAyM9cG6XI93vX2H9ZDk4qX+Ky3ItQ1jkfakH
U3VSiovBcxp0iSCGC9TwhBYP7zGtuA98PcFJPSkcny1lwt9Pwot70uUb/rBjQ+/1Y1lvw2IJn6dJ
TX4Sgb+mwbsvZSIj45cr7h4kUhAJa36RoiwWyHfhT87CAc1PGUVS+di+4/FW1hhwVgW+at1DuqfD
5ZsEf964Rv2CZ9iDVk2/+Ld/8g5RccwI229xu6i6YORW/5RsUlqJSDI4Hzj+rOQh/k6RoM/4bVDP
kg39Z17zmcPufDf1w7L7vhjwW40bKHI9zySVaH7ATB2Eo+7weGA2HznEJ0fX28+prOL3Cb4XMMJV
cjfJ6yr3XJ8Aytinv0MfbP5cvZ1gcWTEhRCNEDK8YFPDQh83KVM+RPWvYQn+yJAfghb2Sy95E+RV
bKhwOl/owS72+Ncz9c9AJh6ZgCrsvoeJsDP7NVQuS2mAsa0b+Ki41ylDMEZFsPxK5BWwX/TU2AQQ
j3OTgb5/paJhR+4SZ+d3zeli57dSLzSvIEnTOTPmEEwIo++qRuwIkxaCbu+EmPGmoQmeBylFj4zK
5oA7fcsLDH2hJgTr6MqCTzHWQYfw0kREC+v2s54Hvvq3PfmujdlW7sRS3Gtv5JhAwNpi/MMHNKiJ
NTCvGJD1ZRoyummX+/gp2kf79sH/TCHFRgbi6mnCIHOATdM36LMwDUO75n6zYRiJ4IvWsUo3f7rd
WEnqAuONiN+gwFiwpFDufTD71Ds7wmcM3zNgPndjtsG27R3uj6rWo9Jy9wLGa1eJ5HtaVrIsrkeG
T4jWPhxFlGDjmPhBiG0olV9/aDcyg4ALnBcn1E5GuAWr0jBZ4DLDM09PrcITvUAgHgZnByfvgVVM
VYOgHQdosWtVtb8IEEBhxETx3zS4m/pkCubTmyn3fFJW2VfDslSzrWWhx72jCpOPYdAQxwI7i0AS
GG23hgZhfAqp/7df6NmO90uEB4bJWyNT0UZVB1HaSKXdHd5F8xNOL6nVUDVJCVWtdnYZEETrDe4o
mq7/EvoqVk2qXCo0Di10wLOjDTjHsmCczwlxJEuzLxSRFIc6ufsnIb6O6DazfYOnjaClHm/gbbFR
qzBoGPQHl0vxi8xuasd7mj9uf30jZ7Us23DLOOit5XsTQl0yxQY+QnP80xg0fYpq+jLn3k25fUkB
5jllFQYJAWPija9vt025/E3Ev+Sh1kKBSg+w2hsoasIOjA/2OcGCgtJt4QBDF37vk8/WLEkTfl7W
TIZZRJEIwH3tpuyXwS943RJltuTZEJ3V7lrGI9P29R6smCKdZT+RZ6ENWlPWMoCUZgM4NU3Hre1j
TUiH6xIQ6f6EQvnKNBTxOILUpOZJpcAKTS7hfy7tEjRLo0c+KpeKlPm7m1cCmWWzJuvCk4LlsIDL
jkFce8WA65Qt+w/V+tONChDms54gA6IgoBNtIinPVaoljU+j/OXMsVKNCT7nh2iSlbHg8rAS4lcA
+9gdLudpPEImW8Xk6zvjQUj1GnQ2iPgOhsMVCMAxQ51jKuCVyb4gjaRkbmv5J7HZBq99fEDIwrBG
+aROgValtF7Zp+z1Ul8t9Mw2awJa1xsrE2YNxZLPlsQCDThN8FAaZiZl2EUKNYGxp9sINmhB8hby
3nU42pogL0pT9LpLfIurxY+czBM98jONpdXzcxeXQpyHEDd1eqpaLqPt+Ev5N9Md5ges68ZsOdyZ
zNSB+LsduSBeytxRzw7idfZHnyaMcIW0KCr7FnwTsu6oL0pS2aouC+UjZA4xA85+hNS50w1TK5oe
PcrxpotsABFaioVGc+098YGyaN9JE3+v9RR2Oo1+kfTHe5ahY6IEE1B0M3IIXQ/6SZCePtwZOFpZ
guiBy/3eY/nUS/lGIbsfbsutbupazyMdHJceyEQMFYerq9STjYX5IonrNFvFeLNn8SxuBlPBTWV5
rlSK1ivwIhhl5Pj31rMfH/fkrQ2imX9y6p+YPRfiLCFIJb1Qu6G0jfW/TH53AAA6UThJFhJJJSDQ
cXy+o8iQshYO0ENARSEq42bEVNqqe+SOVk/Gj9Wt+xCcBp6NIQiFFu+ln9Z+hQiXmNwAeVWEwjQC
F40pbNUSO7sJ5f2r/MB4xFveO+pDg5oFgn6P1CtXEPNZKPFKdI3QIsQFdfGR8jY5ARGkQoqXTSdb
Z7IdnEMd4t0VFrtF8ITzpJier+sVxs0pjH8Ig8n1bPZL9NcOMM950UhsDkqjVx0MB1z/5otp2bwv
0xD7mf2wwMhHOGcqblvcFubelM/QRUeOLwzfNvooELwfNuP5RXV55/d/fpsruRJGQ2QGPotQ0Y2R
pIdCOVfP+h/IK+ogDqtT9qIXvOGJjtfEcdX16GgD3Etn/FiMRjdp5vzjM4ADIF59MYyH4qSl2GNN
h+Hyf1m1KkxqvHQFLQMpgxt0tA6g8ogSVsNpCAZRBJDXr1ZHEVm7QA3v6MO2jDZa9Vuc9E7NzIlP
cGWw4/r19Bh9OAXlCXq/ki2jORg8nPG6IrXFWMyDgAr7Npk+oKrpGEdFX+ZxqnWWRfdI0a+WmRy2
/cf2JL6//avd+4C+F69JmIun25IY0BqzEcM6duM4f66atIrTctREiDWDtkK+BNSKyswu4fK+xzYQ
9IKfAjS2YaIR0/8H9pptX2TRT++Kakw39ysZWWWTHeknOkH6xxISz6X4NINenM5Pbr4oRLmQ7uIb
Nx27yjAAfuaADgwhcQAD5270Cz+3QS29Q8n2837cfHcdrRJffiAFrPRNY3MK+3CxmRnZa3sR7N0C
3HU8nue6UqTlRZHSXCyotZK5dh/4hrVe4gpEX4iegTUjjl1KxMoEDnwotHFJoUh/EOSl8yoaVwRY
40Ta+q//gEyeaNGHszKGQNKDpaIocoukRgsrM6ahC9wj5h2ypOEDRFzzptTQ3h4zMTv2CwR6YEc9
uHfWfiDntlP8z+lZbv478TzIvtkizOxOh1WyxlLqvldrhHJjT1G1+wWMsBhpryYI8Y5hLeW5tk2y
2h1YdTrlOsgEH6EW7qR91yP2IX3STUBb3KkVVNmFJlhhggmxJEOhVN54UPGJgXaQtzNfTd4rTquz
qfHizveSzKRFRTHCpScLNv0dYW0Gh8EGXgzkcnpo6dEk9Bf0kKd1hdkuzNMiXZinGKMVDhGYAjq1
aAxRyZ0d+XV5q6w3Lr7Cify1oldwrWGqBZOnIqXvmKsrHVDU6ZPXMJgkduq9f/8lQe1OelZ/beIE
ola3dRRuGxhJZymXoVH1SDD/Ug+dWQLFc7uOBGsqP0xQ6oLCMNfseDDMJwJy2Ckd5LpGs6w6xOuS
bX3I1Ja8gW8/jKsCHnBffjd8mV6mTlzyYaYflQw/7n5fXA+vZejAZHghJ4wvJLSFmdjx5cbftPgx
1J4Aa+XwT6YRwTtxmYrD21FHgNCz//828o3++77NppRQeSfFfyrW2zb4jM6vYH31mcvzOnSpnBcc
s/IhJTFZJzAoRnktrtouqhdNfAjN/muBP5Wk5KWQQSKMSqiiuJ5vxhGctnpPbWykIci+J5zPZI52
OF56jeWVfl7ecNBOb+ozgoc/xYbbTB4TMxkritSDjMfjA4/Lshb131GCTuK2KRSGs7WhR3J+U+r1
6Qodgh+y/RjECvtvIEJ83ptbfnvSuFHQFekzLws0F5ta0pTkrZbgknSJXEPLXDw2LXwR7XY4yjQj
dNNNdNEIAo8ZKmOrP0T3iBirYlM5f07GKZAfs+HTufjDRo4NJ32jODa24AFcnjQM9uKTAkfaIG2M
GdYAuYJyXxMk4kzKFZFOOU1Mjf334vJNL5Sc036ClxF8ZhVLtCvuJPZfKoNMhaYfK5JqQilVK6/2
tcPZP8zb8qdiQc5g+PZy04hMYrvojNljSmjmD5QhG7UpPJy4ekNozJyKM9ALeroGlVZ8nUWJmurd
5qWYDMZiq/fD/UViErONzezhkiOCQudr0h+TCOzJei9NazgFvpmx0AyYtaZhKI62ryA5DT4OrwD5
FSpnr2ALgHZ/VjQsaDflO6vejeFNNG+fUB7xinBYefIP0Zfk7/4VdAWsTcPv+m56xvH3WBdgnoYv
K6qRYXERZGil32aLkBpNnky5zfnCt2KJVJhBdtHuNncBlJlEptQU1OHpjtAXJIK35H5O+Ub6Hpwb
zulHo0GO/hdboO2lUHDK5Y+DxA6b6ZrrWPP5FITi3QKcu68+K9hWduO0i/Wlsw4ybsU+fd4s1zBx
EUxKryiHhEbpnfUlMzri8VojaWGZYiPKvnLbnXGVFUjbcwZ/SpE/bHHyGmZ5bX8FrcxRHKQrQML8
c/HepP3m7fJNXS2CniytTJuDAwA5ALJtHRGNnOC69bAz2+La9IU3EhSLZl2oIzEG+C9LD1gqUS4r
Yf/UxJwifVh1sUMcs1+/OFXjdhbj4pwSkUznPxHRRC0xahEtVRPEiDiiPJg9TkbX63ZIsBJVDe2Y
sklu5uMkovhrNTbctsKJzZ7S5lOIzSyUmP8XqUuQLQw0JeOFd/qHTuojaydeZo1pLeLWKyp0V55L
BBL/5Oxthft37zekGAw4kWFQ3P2lTNibD0tdoJ+P1QQd+7gHWBL5flN94uzvDvRxUzKCokmEM/gP
6gVwGQvRp07xSJRkKHL/eT7ZIQORz3q7bq74SzEJB5M14DACtSH7qLr1BU/oir7PP2DkOjlNStOZ
KbeeM7A4tAetQVaqdYCSrN+Ol21rGqjQjHVhElb2pMSrrtZlxDy9oSn/FbrApfZgK17y3rUHeeeB
8M0QSZJdHO7f7vo5DdoVS80tqZofiZcWLQ8JtBDvlTAPuSxYcEB7py/nA6Xtx4AVPuLqJbiRQBf5
4yAX5Bknv51QQ1SpHXlSeWxJEdAaOqgcIGmWo03SBmOCexXlvGwAk3wqsIKuXAiDUw4s7Vk1d/w9
GHQwa68mxZQHwstYVgSa6B3sBVeMjj9/LVZfBLK+mXGIUJh+pKfGFGQfw1yKAjX1tim9waagjl1r
a8BO9WyCkaReTX8+4JhbwE2X7mNhydw8d5wGHteIJxsjlS3Ind0KceGwlPvV9PFUBwVvcoKTzL+Q
ngpmkxl/T1GyGr2MRI/zh86SIgX1HPVt+9Ia+fYCiLO9+9LUhVFfXdpcuLEovFZf9nyceZ8tKOt1
kPGNKEcGweXBUO6owiuc4spbyeCz7qYl3EjRYSIJvXkhKYU6BdG9OZxLGHLuFr31tQVxNQkRMzV2
RH3T/tEGwiutBGyjn8mZwzC9PbYjzl8DfaU7wcFpcmeIr+DJxBOmGTQTg+Ptv3tF45y01vIVjQFO
Rx4TcJuiTH+8Jn8FlUnw164WaSETzFlccJcuQFDtkiW4vpx7qBQHlVGDi3aLmUNOk9Cl4Jj7daMZ
jy0OCvOvdH83HSmC6TYIWwR9SY5MHSSSsQliXS+Eu+lKnFBKAAiGjyTO0MzDbTLIvI70SXQZANxS
2vTTnqjmrH4jfiqY7JCfFTJMUfnZUI1Ugk/5q7P7ZvO1gNQvSNx9Afv76TqXNp7tFBQ19doaGADW
qp8+UTj+5JebgWcJWZCn12bTUNADZ/sfUz3ej9yJOqQBMq2mXEMUvaeOrvWC0EDeMyYX3oZoYhCv
Vb9bnLPftelEuay+rOxpRF5CLN1SzRvAGMUxtsZHnNOi0aW5ApzmtWvYx3+D29wAPiBTao58yqNx
bDhRscU7abqow20dGTJY8z5b5YBcI6vC8nSrMaeexHsMDPdt9OZK85WgufZb6Z/8dElOeyO09Af+
HEYWKyAOhVLaM9S3f+ZGf1ulHY2XSLQ5nOZ+bG8f1jkAOaEjKCxXDtKX8suR58AinGboiFYO+0cb
QNVzkj+DQ6JTFpl2gyHPryPzfDsN3PBkqUiEC6lM9g6SpUnU7omyE6Ol5ORasAkh2OO4jO20WCTe
kUaXusREnAxoZvQZMjCFZXd5WgIlgQNj1S/kPLA3hzIVf/eEa18F2nQmf2jGOqUQUjpxAif2em0t
Z9gblxkVFboNeoXsbKNYa20xptDdXDna8+xB0llxP5BJ5/c3UlH4ckiMacavfudxefvab+fpU4Hm
sy23F1hkYAzaWRzOTEwaoQuOdK5iiI8LLZ4Xy5Mf1fz5AMJGrsyRqZNxFX9PMNwebQWLVLDVwkcN
eEqbl90PFgcjFkASJcJaPwpLfjFHx+LcYt02v69qt0J0jKn59xNpeytSJkm74A43Ocfmm6kWCqa4
NGwnOd6oMcHifX2FdQzFTGF3RP9JrRqdRSVK39HU129LTi6h5AogXldYNjXngpwyOQF2eeOejV70
Ui2aARJw13I83TtQpAq/LITpqrckOy4R3RaJO5+WjXlXgLnrUtIS2jq8v0wGajF9hRMhX7GsKbQe
GLiKPqrnJJQwnNH+DHlXs9a+E7OMaUJIAZhvmAMbPhT02zfvZt6qWom4q+KkZB/JnmA4nTz/IzIR
oXdjz+eug1CKa2I7D90Kxh6RkmcVElBqKWQz0VwuqRKUBGwNsayLovg/mXEun3RuAT2QLhAgQwEl
ElfxaMlTx5bG4pli6LVhJLMjfW6Zs0gbQcisB6xbMQPIFXcWZUvvLn6MsKsY8z9M//zamlVzBYNw
hMHNFGzmJTYGtVP29CuL7FYz5UZmPHZfCz+MUg0pgvFC90wZIshOF3Uo/38NrSBIHaESmgS/RnWg
Tkg/VNzFxubimfk7ss8op+rKHvmbphhrNL9Gnz7wRU0GVGRm3bRAOMjROHSfGNRDA+KQL53jowSg
1f1Lx/k7rD/0FzAdoq2AL0d/cjueUHgvQm11FCN0r12YtsJSodWbSJ9c+/5nVd7tl5Id60qOXY6W
WGBpOjX1UzwRWEmzwR5Je5UTeqd1trqiNEKgx2M5yGS/a1E8Hq/QLW90w4PzPIaVZF+hZdSkXTAb
i3gfMedGdUGvvz6GGfR5Hezu1hCuR3f5P4nBug/Vh0uyI2EkAQCoEeC0VydLtW4sIeB1l3v637Qj
7rzy1ZkngBou9cszml11Cb/SgCCSl+R0fwfnhR87qnFF2iYoDxZ4KKT7rgDNXTeiC7WKOIVpitWo
u+NZLEOQOBbvBdksphPx1Boi9D0AFsJO8FNo50fNULpp9zWcEAOnKpWXbRykDKaMTOSYeqshHG3K
Nq6Nb0M/2pGYJVlzkDmFQ2SriMeWMRc8ahdfuth2N5xGMLbLj9ybB1bTIvpy67S4ewOJFpqxRO1Z
LW15R/xYbm8BJ4VnCadBj964voySX4KnV1UiXl4hpdquFWahhPd3DoWUfKnF1MY4kdzk7Z2p2KKB
lXfvmwC/HOEKSO7PQLNVoKYPnpR9XaDeHvVixvjNJ3xL/infrcHs021kJyuyDz4CJVwidfm6p2cQ
TPnkMMn2ePpZZjH8W7byL1Nr/FYx7SXh4pIi4xO8F61Ul9RKY2xrN4paj+TAovY/TNRDiH5nFJ2O
lU3JGCXUWem2AZXHfMWTOZ5j7EqbX+zVq7NH1wXap3+ZoBehlL/eo2JNqMTUlS9AB4nVQ6Myqa0n
7uqDZTyT4KxCoYPs88L4UcwxIfojNmcHQ6wOF3XKSlZWofPjCRtnAeSYQ5t1ZG8Nh6otYuC3VfNA
1vKud0zPhA9GxnC5ZHzaRpTuKW6DVZQIPL5WECjKJTg/C18mdkRX53tfyRrntFdADidY8zRuYJcC
cZTX5lrd4lavCRUPzZqHv7OwlhWX/gXqDQpehaFnuAmHOXVOOX7zb7dP23y4/rgECeJhC3kxco6Q
nZryEYKhtQ69W1pmIbEpQXELjaNWo780YuOGyjB84Vsb8dZ9HS9rS10pXy3yB2FqSbDBtYTXsges
b4xyWP4Pr4NLQGRaR+WSKy51qqC/38d9WoyQ3ZfogVmhi6HoI0CkneEdrPAV4VAiPaFU84JwZo65
kh7WuJE3IHUw5y2GOa+mIJHCJYb+iFhOhjjGTm5/gmNE5z2XgVuV3gcb4wCN7YAIVDCL1/syXrFw
ddXTj4y1ArwBsyx5J4waSQFwkQQqsbYWNOJ8N7C7Zj/QXS3quJN0H98ttPzz3xXCvcDKlhtDOpI6
0kigLwqUXKWq1kliG4f+hRD7ZlaoGJ8V1+cKeQKwnsdO0FEnKJ8H3mlldQgh2wCL6dAfbyaGyN2n
yu1nDKWz0YKBqGcX6puzRReh98Db59H3PEAGOIM2142hqllCR9fYXFLi6B+XSi/yyKGrMhMBAnpp
QJrBmksH1uDQnmiGW3gX++Fia8p/LUth3OYmeHHQifvWBATdU2OLD8hilZCN+4wf2UH0nqHr0UPa
QdLmnbuqhjHiibLeInxVygdQ/wwjDytizwOMomIeQBxku2G+UiNWSIbNRTISk3hXCdvwdKeNMYbl
AD1RzOLl2Q5ThyQHf+r7OMjx1/8s4pIxzz3gKG4A3tp3ZeWc4PpLADj3rhCckIgzJwnkMbL/on0P
VIz2R/1SVXhh1JwNWk6PyCgdUQHLCqdgcWn8+pwpzgGZJ6kNcic2Iq/32SQ0AOIxv5bLUDep2rCE
d2L7FftzxNQ9edqFRdPL8/8oVX1yPvUGvcTr/BK4qKB73QSvRG9JXfVwVzjJKrKKUbWb2O72aa/D
TrZbfQpH/VdrtkuTwS8n2H40luqfgnQBXDAgYZewMWjYKU+riGwE0EliK99oAX6vpgWqhYmfJwK+
bNIv/gwN3O/IS4bTgx8T461zhg1lG54xxTIugX80BarQoz3YkAC4ZTtBuqz1peeZcB0hlDA1hPEV
i/qEwi8Uy4s0i5APeLNmFL/0pTaFb4AvxgOq4bX3dJIipyLhhT8nozPTG2UFEIg7dPkoahCBXaR1
vblLQD6ChxwgcZmzINvZXDl0iQ7ha+GvwVNPxpjzDUhR1lO3UbY0eO84aj7hhpvaPbmmZt+yQ0/5
yr95/uNivShzUGMUErC4T/Si+pHSZfjVIsdEMI3uS6w+MjdjmYVnqhV0td74cDA1ncA/nSqS38yO
H78tqObsuwvu65rbKI+k5gVJzrpAxWUql+ZRI9hQnkZTDJIfsCgHmDy94LnOmX5vR1q4n1VQSo2/
7ZSvA6twzSBpfi9BENEuxQxB/yY8LwjR8Bok4eopWfB2zQogn5S+ISAQW/dRsZuqgztffS81qOJa
/RO/X+rC4POx/Rl7LDBIVkhOcdFB4JuXLAwgomXhvytqR/HiG2YZXKwkepA5OeBjGcJfh7fypX4C
ZkMgXLzlddlq81TvMs5Gw3cf/DeGm2dPeQdVitDxRln9pHHgmvB1qV3+Dd4vADp2uSAWZZmthTLn
k1LOWl59D99GGvAgIn1jRnfYlgJPtsC290qk5vE+CvFfxA1YwoCqfyjglG/nyHaFJ4h+QrP1KT+X
1I+2Z5i/TTHVkQ4na2leQ3ezjV3DZIaoZzIaQptjBhiuG2ltJmNDHKdG3JCHyZxTPT8btbHAsPfG
9IIGnmqL7/u+VeGIbIHcrd263o8wE/7H+elQ/6ZZJAFEU+25V8whzcA79J9wJPbicdqu7hXig2Jx
WfnBnJOw5TMl4Ma2v251nKT0u+gkGFJoezNqevQ7/3bMgqEGUSrLeOZnwtvAFAIuVvqg1HJSd1aD
W5aOMSKn+UCZk+xqWktnSuTHrwOwXG+nrp8759i52fUrTVHfU5UnJBuESitKpjg5IK+Pc78c+i9b
DZhHzGxEy9C6n2OuYZbZcFj4dbyed/47pR+pzsMFNOU6NeGzklrAggaHThIOIWMlBsDFEkyJUhiO
z18ma0BEb+ieirAf2xx3VWttv8QQBUP7haRoKYN7Pumv3K1FU3wvapfORtMq1g2aOSax8oZJWT+P
O66JGNSAgaQTJV7jcm5AHwSPc3PAOheTm61kTfcT5f0+VMq8ig3wvz8d3B6uS38Yr8IQAh2luc7x
GwDtZ4HRQBA91aAUIOjsboc3MImzAb10lZ5hM/ajZFIH820Af2gvuuCoDcX0U4h/wyORpFzuXte0
Kfk9RWTC3EkNeNB2Y76jxkhaaaNIqPkdzSi8TLMb28TbDJ4GT6OU2MRZeEOG9QquNKRTqT3VT6Yf
1e9BWeSnzHnmOFIVP87z7LwiNQbXIiT0QX/qFwsi/OXRN1rlDKQvipVPbn4NFiakh9GTiOQ6APwm
4T7HiF84TTIF57CSfHLH+U0Q2XvYJHegsXU+Qw/bZKIXy/EEsHr8kItxg8ft+4VzH+To5PNIvgxi
lYRcGSGrum3GaC7XC5Q/OGmTAViS0jUcIZkGPcYPcungrkFDZiaiQlfbZdlIJInA4NYtXNMiEXW/
hqmlVzpeyLxDGMtkjQOkIIMpfkPb/k0gG/wlV2QnRzQuDzdhiUysDOI4FJ3Zfhihbbx1nP6evJs9
YMNTdetPUkoheFUace3LcOpBiLjk8BOs9bVp7ojgQUxhVcj7mkeMxbhbnTh2PMu42OAP7xXVDLZZ
4znoGomr4LlsTuwg2k7GOcX1QP0Q/cpIx8b4y4/DVc0OHg36+H0hDJcbmouAb/tMhzWNgbbVChrW
/7TKYozObSBppMhSNQbpnLiU6zFc4CalIoSxuJQilxvnJ8e2lTIl66SEG1uiR8RrVdfmPd0eL0Zz
oIHjCOWuUH65HRZVWxuL4ua34RprEz2hKrFVzEU/4Aew3+cOhJZ9SxT/ePrsNSuW9kGVNrmOBWnd
eAPMeUdqW4STaKpyKYeR4TaXgKF1Eq+/9GenA7m/MiAgvFWRRopM4TpUfvTJmQNoiKuujdtAk8Rv
DfIGFuMFwXNwWn328Rw2t+UEsUfs8HTsQlm5FVHKtRw1EJOQvjh2uYZDTerHps84soy6/K45baiZ
9vIQJ1GtrYojnscJtTYNPtTpTLqOo4yKJ2QaehYA6Wve8wlufNUEMTFSja40RsloQXOctxs7g3ou
k+oA/Vuip3r7kSvtKeUXs5vFqhnEWNLE+iqqNlvx+ZrbKOyu9825UsfAkxPpILpge0DAEOQ7JXkR
zG6G4geyJ/TRPKi0sFBMLBdmXOCKAOtl12NG+JCIA1XaHbPbhlLdqcAqnfhMeTOZ6+R6f8RZJvPq
bl3kGso4u2cNWgufp7fj/jtv+L3etX0Ui+rfE5R5cHedSvNBc4n3st3X7Dv0Mhfvl02zxttVhM/1
fZWt/FDRC7Lo8iEM2SG1n7wQRRraI0f+SlUJ82x9V/acTrKZE972qn8HttRlUX5EHzvNUmOZyAQ5
DUtnsB06ogfeeAybl52Wc8cwPjYoYa83FEABZYsENYT9pHnZ4EZPDQNYHj/oecJmL2GpkYDIIhxJ
bTnrUhH6fL/Mv7r03BQ0Qd5igSjlJZfZXQZ+g3XwZmzrgqpABh/ippSQa2yVOnbArKpYXvhPMB+I
/kXCtAqM3xBqyCpn75hnvGzSK6r7qYnTEb6kgczStq5LQ80wGaAJFh0UDX/O7QuZejpogQ2jldyl
o4IdnwNx/6uL5CbuD4nPkFgxWUglsZr7e95Jxa8H9u5g/3p/nyMWxC08+R7sESfpG5nuohUjY0FS
1H3Peanz5ayyMTgKQT1JfixQqT/AEYib1mbVJzMlgEtbk56M/m4iqluMlXpC9ohwo229XA+61EN6
CDNfKRAGcra73OT04uvHZPel2mxHW8bHf4cx7CQBK+voVNcZl8GzErPK2H3nLZE7PwFxBNH3fOpI
WwfGxHt4ZF/QsMEg9XaXl9cgMlUzMVJAEUTItrHTHeIetRALs8woOBVRj1OxU0q+bN1endeB5teU
hmtZSXBcfKXAPoI7MbZk71DUe3gdrCb0MSM+zjyv6z9fGW4fh6ObJcA67d4jPnBqiEGTTu+8Fl5k
hUsu2csstuDGk5/VWizskZr2Rw8nZ4HG0MoWQWBK120oatuzkaI8glUyhKYtaRwb25bXvgZcuvfn
YdossDf8omtY9kGztQ1fSJzt7HNNodqe0jBuRKze1Ix5v0s/6XzejkkKgv2PdTKzg3Psmgb3dscH
seWPjltHAuekfycV79PC2U2NLMEWl3RK9uTpYPijIefuBsvIZgoYYpa21g0CMF+SrpZW3DHpX1j9
jgapcymf3bfcooTnFY68t5v1q68w/q/sboYGLct0EVDyjtc3Co44DfdgvEDFYZcf+RIyEVxUozFx
Tbo5Kwp7SYL0sevYQRoiqa3M9ZsguzOFDLY9QnXjgQ+ftI4AiQIE2SZaODsxKbbRhCwj87BYErEj
/hMun/GYH0L8Me4gO0ylvfXpLhfKC9ZqXxLDCz1WlL0tESRAoxXLPc1kC82R+64sMoUV3o0F0OOt
w5jqKKFYC3xRWSzEsBGmI1MzQ3KjelF7xd+YNP1bfxv23VJb+UO+yfSWOScL80DuTY6YHsKIxOTT
fTx3C0slp3xJ+TZ5uOn/YJekfieI3QyOCJOIuxC3SnxbLmQeCJqij3FHa7lgOO2fm9S3ZO6jrnvp
pIscS2JdxdFyvVgHYmoY/8TOIeYo/fEmTj/SPHoXKvArgyIF28HK7w+cNSlkywhj9TYvPoZhVyyk
vqsQjmsAzOYywgYBUivds84qi5N2LALZhhPtrMbJyUcKGYqMdVB2s7FBhqqfOdPM1yAPyc1y8OvN
5j5ZXTovumOyBRcvXMgSlgaNU6ZuUiTfjltIppf3z8iyS056EaseZArgEaCVxTHzsQYyM5N9OqS0
pGDulWOKdgsSjcQBJb9dv6snq+x0cw6KYn6/fYzhTZ5M8EVZnmKKO0/b6T5EVdODIUmRetIjJnuC
C2sKwmOnjQPNNlTzQyqZDA9jZ+Fc5hepbyhnp+Bogdm3UpWNsEDxNJLaWJ9eKpcA7W+tkNoNcnXB
0C9KWdp2mhfuhY+F/tB+DBOQ5UXMu7UNTyUDJks7mqfAVg1hVBSg8myDbdofcg6uU7hlcXQAS/Mz
MfhsUM8bln0nSPduxYEPX9YwQ8CFeXaIMXAzOpobWUvpLezPb39HBmPJs7SGPy8xHpbjNP0btcpT
8iyffCS3W2CV3yvmbhrUhttdY3XgIsCIttiUm4mahKkGk7l7Bm+Qr/WcsvnO5kt6A/QyRjue7czR
gaiuxlLC3V4IA+r63JS5xti+CZ8COBF3ejnZT7g5aJbFlVQ9RnkeFclGi7Z0IjwA5AI5EwT7JRUe
5GAMynDWl55hUJZrAevKwIaNcyZLpSxkrUXYsPbl6UDrfvVRX2+Da0xJal0eiSFYgQtQsm+zsuKs
pdFfomLxA74TnvB11j2guYphZUjrPO+gnlqmrw/qZdqz5wm/tLO0h4O5EFXG66qeh+cKljN+WcSh
WGfQElyLt28mg9Rxxk6VmGN5GGZTJ1a2vRiLkK89RJT0tHVxfkg77x5QgcQDRx/4rkkpWJV6Z2Rp
3TufhBFQ79q3Kg4WBUjbm2eNZFQf9M6HqKMHY7DJiBgoa4Mw7gjD9InOUiqnFiUL6fvGVSL86Zsd
XPu3HfT88IhMX1K7fx5RM2986JYO9GEDKkYTzWk8006T9NbvE9PeUs80A8XM4ATXVeCyqXjwtf+6
WYgyvX2RtksGy3pME22nZG66gdxemnaaJawXMcEl4NzPFmk12xtZXe1DZN/QZpH/raZsJMvY+25/
IlUOEOuQrgVpXzmrub4tmT9A/HfJ8RHsbL2I8EI6cusGOKRbl11eKZjXrwpDKUgytC2HtIx4+pnE
E6kAPnQXmaklkWRfwC6AysQC4/vp3VJTC4oVEYHAOdypVMUCDZMCR7VYqeppyh4YDXrcMBt+5u6X
b8UmYXXYZBpGvqO7/+dKfpFu/+KCfRop3ZL3bTXOhPgufAdRF5BMIyvK/80qFONKlW2mmmroDkH4
y0NASQHCJ79Bq/E+Sct09TaT+qThP2KyWO61na4DalvQN0W5PSMBL7h8hqpZyMsOzrIzLXXGKlP0
0/U5zbUpIwmuPoLkEimPTtDwRoLLYYjVpQHk85xSD44BnC+25n6kaf/gWW2Dvr69c5ywbrjCjyW5
JxMrZN7/1YYGaujmBUQqSyEUs7PUbbwBQiLM8uc2O9vxWTyFWE0jQRJCeL6Wm4SlN/TVs/4cJEKl
wICeIOXfsXTFrcK7+QA0U5m+HQzVhMdQCP7NtQw1oOcAsoTZI5lJj4VQwOs6f1TM6LcK/3eFu7QM
xOA0EmyqIl9Uxrv7Ajr4LWL+zGdT4N1kvPQzEokjzNXoIdf1Ce6Rh4SR8xMo4zd9ZC9AV0IsceiC
ksCbIfhqACST13Ep/7BXiRIm8LXd+5S84lAivVAOynYF5WNatqIF6ILTt9oP8BmZr2Z0sFd+c5z1
+SQ0lE6jiIy5Ira9316XShxr06aIf/kWaJHQtXETPdsy5xfB6sGi3k/te4XGyaworrIGRGImv3ct
C1lneupf9P5DyWxM20G7+PYl508HBHetf8183Is4vv21KO3DWh5CsXbz9bMhBrWUc6MKZL4gZ/+K
KOUYSqyU9tVC9RIdHLA3Atm8TA88YdNT/qdXE0ANIlc6ZVQCB5d8fVTscId7SIHcZT2MRve43xHS
UvNpIihGIrUTqivP9Ovfwjqi1TsydeIbTNKlcVG2dATlt7iU8moxcA+GzvL0VUQQ0+wxI1Jl3Del
aAP2B/YWFuzi9GC/WXzp8lJepIlaLawpoahWQW/Xcc+Q0rGLTDi4OHyLotU60uOBCFMRd+qG0wmF
TawxZgAsMVRJgyziuEe9t4enC+W+1PYnRdaJUQ/1fQRVGqcARobCRmiLMKgLwMBDzabBzyIXVyFL
+qz28AkmuFyFoIBfKKKczpSawWaFvxKV4HmI1Fmr99OcUFTC+tU5PccCSvgebrBB4D3MgGOjv3uq
xB1N6Y4bMZY/9FdmO+CkRkHaDuFOUF6QUZ+aFkMl+yrSg78IOmBND9F5u37pfFdq0VDsMFlm8GHi
+BzFOVAjybIN0JpAi0Kmq0LIZfRLh2MW+Iwpkof3kJB8fLk6BeHw8CyuhTcxZSTlsW5Mp0adE8gA
toFdSKemNSi9u2kzjHUbt2+iw/XiyJFA2aHwxGrkfLS8YuZg3QfBdqveDCCpCESqOXSLdbNgSQGO
2l1YawV+7FIgLU2oZKvrnepxSDgsGSc5Acgr5+frYM5SFyO0u6DqDWoVJR8mAu95tBakedr23bvy
0FvBNiZrRLDnx42pv6St0htNaqWiiAynfQruJ3mXwnF7RnNktvW+KUWyS1Fkq81+S6cg4LEXkBZV
X3vYXYS402r9QK5CHXP4suF2aTKYHbitJ7ueOPgOC2zniUMGUZjrVWsuh7jmQMtcIzHQxGAd7oDA
OGOd1iF9VhjIf8fcF1PHY8KDC3yGmu4fNsXKhf5wBsKzGuQEj5xZwjuy04byXenrISJA/84sFkeR
XN4YruVmInpN6d4H491BlCCaZpDnZhylw/vm4O4uDMMrdDH592tWpbgXN1gVY1hrCK71mXenXWot
G1PIzFswWPwz9Rjsy2Ze+tuY75HwlIxC8vqSYLvMlsxcJgH2rIpkXcllh8n6vy6y4XndIa9HyNBH
8YOZYT/ir7zWUDgHqdgzUzdS9amWjf6KMTeMXkonwmkfVf+qHeyhfmnZzY+oi+f31G61eukXN85G
YKr5ZLkRBbVo5mmfT4XLcyD5KgawEbhoohN3xlJibsrUyCK7ryUAtQJup87+ge3pAwVBwqILttr5
tBgkvKQRw0KsvQtywqcEaiFhji03GwX7quFSTvtuccb/hDH6YKF0+QqFne13aw1KW8tbMXGKnUPu
+cE+9Ly/dFZcIBIHfd22Rb8adUJ4A/l54/VbxfwxSBvXwSovk8+KcQhE4lKZtyjInXANblKXFcto
VuWD3bhmV4baeZqVrMgiKu4f4E9UOfbBUaNMcocTgfbfPSU/P39zUw52E1zwWLFzzrClq3Qf87wi
ls+ICw3a8V7vVEVJ5VRiPSUvSg4iI6xULfqZwbs926IF5Nmz6ANOe+YM8aIw/973T64sQJneUzG2
xnDfCSWNdrjVraASf8qyBpUrGlQ3+pb9OfAQ7Zwvopn5cSQYibiR5InB8aVBxwisBRZt6LyoGtHO
AL5ttHjEpT9hO1t5yf/exup5OMowvIkEuuGJy4uT7qF1PFL7FEcIEIZ182If7gZ+2pOAF1KUtX0s
wTlpW0c/2lc16u1TmrABrrfWaGceDElNOKOj9V9iOVfhv9YIYCMmR+T0M0xedMeN1ZXqamaFaMKc
uf4ICjjyWu6TJL46v2WZ5e6urC15hGpmNRefcd/ZqkDB43eutxkMwUiKrFAuyDaN5lQgEafFWP1b
Mku/AOdKAJK1PYUY0/6z/S9YqRChWL3xB7Q39gYLRpGQKjunk/0LAJZjhtG9p3qHRDs0UFLNHWED
N8ra+IaGXxpplZS5UqwoXAW98aXysewxqkAepjlEumbZ0+TYbHBtkN45jq0d0Vb79lpTsVqoEQqP
DStbW91BYa7F+RKyDXdNbvzTsVbkEFSJR34D1sNBIdsK6mavlb0/A/gpQpQyoQGd0u3RvQmsOxW5
10YTOu/Np0L6tadA+BimnFdRHdOrexJwDoaCut9vUhlPDr8q2ZYpME4LYiWhDOcyHBDCluGqT7eP
8Ba86hmF6WI+7xOiYqdXJyoQjEqXqRAgse1mpycCQcDtV7On5+2StX3SRZBqhAqbLYZxIqPICs4+
To9LVUd41z+RZkwLojRj2xg/3O/1NZeaXjMrskYYzSVmUKQBsvQ/cNfPeCgQGx0zYDZiDTCX0roy
QxEjyjtzCBiP+6yMLI2cgK2Sza+5lXjWR5JXROMdwUypJ4tGfyj+gzPw7uxq1+w+WXnCmkY8CvWe
0BLDJpSUCGvvNi0V049UuFlkxjBFBVG0WoLUDk09sq1VEYG/74/xJ1VktetPCaKxGEPUcACQQIhH
C1q6ATf1Tp7dT0aXHvpoc19Xi9GeO+0W3wnLRP5ocRpCDg8OS303M6LQZxYPWtpNPfgtoxFd0h8M
Ov8J9me9O2UoOVu0kyENPApO/+l20dZQjaZ2Jvrj5Rgsbk9jNdcG8BW3U/0Gg0G0CikZEy0Ge1pu
odUmKkpLSYJ7bkOLrZMT2i5MEcRlF52NfcS1ytWFTpO0fOUInZjOzHUzPtlLy8GcTVFn9d6z1KnL
wH3XHpeklqTUCedLKx/iWPNOhTaDFqlvM2dnTyi4CwNRP6Aw4ehZSV/scR+F15wZM13vY0atM3+H
nUCFq4AiPf/EyWCgaenVeAt8o0j1wWV60YvyrET3dvM0tW7MBoD0ITQuyNtOVv6TdMjrj3m57u4X
H76FaE3DQNxNQ4WSg4+MhcGeHGnFp9DVrN6nKxf142AaSyz0xTMJbomf/7oG9H7lT3yq6UX1a0Vx
iwc3CocbfCLycOY7vOlA0iCDkOsi+ZIsh/uCfblbfwh4FMDkms02BJ2Ofyz6NNs2GL/vWjJxrUYZ
4LgxHiA2Kp8t1K9ykYAmvdUfgaoDA84+2Z/Qd/0bj8rsKev0Hg4QnKw/Tb+3YfcNwWl9fvTCFz62
pAmaWNapAgvZeHbcvj3bmCad9sajCSjMDbciXyRVpFxHvac5CqBOuhOYWsLTmIMXYjH7HXhFgYes
GIvJoqP4s1akplFmq8o9aVmO2CHp5pqAf+XiA536hXjC/Y10OPJ85Mbygyth6kxVPOPvHngA3Ww1
dnoTIOiaRCsyDU20B57pijg59023+aTZexXQqKzzS+HFfkbxf+HjJGfK4GPGjuays/HdeSUGpaQG
RCqEBxsy9RI03NCteOyk68y1QMRBBNWCG287wxe7LV2SeB9K2wZnD/d1vOGDvqWtNcYG9E5z3uMm
C12Fp4MGgfSC9vbn1ZgViSJ0NM3kbgK5rkUBXU8ALyunLouHS/GuLN5ZpnMoQDAAFaEZBymnre9R
bkqYUjirjUvIGqCHNc7NreI6yGnc+nyvPbhgUAljZy2ArBCMIGbcr9v2QeQF37eA4pLPXa72xt/h
YeLuzrYkHvKuRAyOCUI1F5B08QX7K12m1sySRH/WdprUznun0k+C80rqEUFwS8NUxO85GhxxWvh3
7oZqE/tAC0Y5MKdy04CPkxEp4xgJLsUmD44bPHqLmKWrZ5AIkzQYgOK657kVwTV8THptIj4vgJmA
vJsf1EsQB/miN6eBU4Qn1JV+fF/mcb9sYcAV6TK13p7Wgd2duUq07UBNQjyPE0YBjA8tk8pXXM7G
SzsyjXOXCGnjjIEl31QPhWAR34qZnORrLGXxCDUnyIAtVsZZlc8bTttGFglvBnyE6N+Ms6X5I587
FbudmORw6ujMl8by4SZPJPeN2/Hc8B+i9xVV4G6kSAIzsTiZF9p3HQwr5ktAdMCYFaOoBIAbi2v9
EhXe0N7fZJgH748kvWPcX22z4fG0AAwcYnnmyJnQlQKaE2ONJr/2/Rsdl7bRFzGddja1cdPOJhLQ
2llRybzYf/cnp2hkVVsGnXZsqmgpjQEGJAovPI2U0/lTMVv8Zf71VZx2jucqhBpAISUWBmWX+u/k
lk/uXoqXqvuqWiJB7o9bowlVEpY4HMa9sjRZ5Z2cQOQpgKDfpRTHAj6gDFdcY0/kuCaCrpKCs5F5
itRT8IBW/WWowWVZB13r0NpDwVdnn1xutEXdX5jL0dxHAu4BknvEIHFxZ3tz5km1qlDT6YEpaXkT
CnFYTfxbmjdAOk6UPuWgT2ddBxxM+uTw/6FsgitR3ZxzWQE8PB5Xc3P0zQPSfdDuWS4Sk4igPAHO
sTu/95o4QujuhlQVauW72l5Tg/o1kpzRAVfN2R4ExCqHii+XeOyGKip7lxFek8k05pAHscy8UfXE
1AnZ0Bgy8FO1l+Bx6RQajrR25GBtlJb5yiXY6I5E11N/sHaAWx/e61V+pqhDGwnmQQXexqA7k68i
H1PM2fKEhCgSn0dPsZ8CqkCGbSBaqAcKR/unnbMPaX3qnNRcku/MgPDxuVK+IbSGK63hTfmdP8ps
dA+KR+FeZwEmWRAk33nMednm7aVe53e3sTl2vORD70U6CdHyMiwzkeeUnl2+66xB4Ow1m5F0rvd7
coM7FfKEHOi4w7V8ma9uBmZ7WtB/Yukk7EV9uoHD557lJxTxX+G8pvurhFgNY9f0mZpAjw8oXq6E
H6Em7iiAf2Gq7TWQ1hQW6epNx9TroruUnE5tT5Ny98NouSqNC7ExvxKWicdAvLwhp4nV8Jb3YRru
nF1fe/Fd1CqTnb+7AekIOWisy6OqXMgnogNCcIDu0rgZEfFxPEIGt7mpWVmEaM/eqNFqq553lZ/+
gEHS914/DafKbm050jvCDICdWzfiDj/T2ZjIEzanr4Ug0yGj9uaXO5fx6QBr4yrZVn0xWNGVOMkt
G0bqfuj2zKSn1JLTbBK48texJxZOfsZTnNfPDCZd+RPxXnXM4xb8BZIeviVcd7H/QVVwK3wMx5Q9
8O7Ghm2ggcXbXppQP+K6/0WfwVardoUvnDvYEYfFCTJwdcIKo4zoz+mGs3bNR8v64MVPu2Dsnvkj
kJBlquAhPUBWIYu0BPOjeQ7/WAFHqY5Z8VV4VmJVKnKSBUMQQBtBbygJ8JOCUOMKZbubQ4HPG6jG
src8s/CXfbJxZi4gAPm8Vxdz4icnOoNC2Uttjy7oswx5CiYvSorZPasuEANE5HXSp0dXfsifVB2X
E3UwEyCIZtLe2zXkViH4GvPD413dGt17CYlB9cFW/zY6hChz8enivvsLMuLpktna8XbC5k6H5bNe
xNmu+a4l28ElkGcV6d0uJckBuzr92rLGHgjliTZBHJ5cFranPhABAswcWZ1xCKg5r8ZMmhqMCmPN
6juIzP04CkmLs/iP5YleotFB4ratAwpMKAbJ8LB4qC3L4gS8hncHwS8OErzJ/zxOdaLyaZjHVF/4
Y9CLF44jAhDs0SuhKu0Dc9DdXHjSr+5uxYTHVz2jZOfqeRu6+DgrNr4tPe8wXtgMDSdEFmFcxfUB
KnT1dT3dIr9WOPhbpHc915QvjwabUhCnTkgUJ6/KmaiKNGCNnbhE3nxX8I4e2IA985Bpl3Q0J4XF
VgQMTUUJP6qnIDvNenT1u0eqj7D+Pyu2bmoNmE5tE4pEUHwRv5T3xweFkz31NA5CuB+3kBDSB/o3
860ggUV8Ph7FkYwsDJWbaSJcQ2cpacBbdjV9D7svZPULO2hZ0tquGZ/uAA9tzuSR0uPpAYFL7FxP
E50Rz3ou/xEq4fQcKsAfVuwOKINlIV49/kx2R4ZIlGcx/tv5GVahw0KGBHdVVhtWAwcGZtdROmkx
KGO+pFskwdklh3KwyTGeSqlrpPTTC+MooFWgJprtQxGxqJ4dO8o4mnqFv2+Y/UfHDF3rddN5gM0O
BDdV4pZAEtyxeJFaefl+XAXRjUdR+926xWA0AUAdRM1HqQZSr6mAw+2dMXtdwdg5pYErO/CxJBGc
+kpP4iUDGD3lGyAp2vb4kPLjia1p7r37FtP7nE5CZluF29ae/Rz+lWUaSe/LsLBwn7onYIk5tmyI
N57ISjWuBLOT2vnIWq46Zu58EJuFwOt6PXWciw7eyEjkRQ7AVxnuRhLO4eQBHUDv5JYMVWbQ9VUI
FePCP27tnbMcsJoOH5MKMBWSWRshXsnOqqwmh9g0NgGytuWv0Iq0Ify6fY2GSZYPpTjudCSySR7A
7DT5IpLDSeIJAvuFDhbhXLH9t1f54Um4oUjtbDgaQApk6yHzurY7z9kRh70VzXezXXpptpftaVnq
syCdocDd2sW0RfUoCOdEf/Jo49jf4C+HRFPqMRHzT5n7AagQwm+S3eq3T+dUkmKTRw7PlPie003T
o2V2c+Qr/v3kddDpcnk191xXR37XMjhs9wy/vqr6jDAyVQRtljZebS1qUmFrVqbixTYEry+E7/46
jqhvTkNc1zuyYULbxCQAwn0C4OIM2qThICZpahRa+3EbS/IrPxpg7LTM6ZZfmD10UusPe759YPCC
AHzSn09NE/dT79oYm1p3ZXdWp0GGP1GpJHbcvhGm7qGlW+Eg7d3Tt3laCKiuXZDkB9PDEI37fw6S
ZqU0f40P38rwojG3cTEfgTQgy6vEXh6PTtCmfo4IGyFno05atxrhhOYE0HKVHB/7Txk13c3PGPlM
tyNDNlZmm2lvzbr/gf+Ja77ZjUftnhqlfan8dufOrNFmuz5rafH4Pep6FBusAJYA4ghmCv2z0lCc
V+Mjz0zyfFSXZvGvEYenTTPNITJqQ1t/EavWHXw1o44oPFb92UUqOXCFhwb/PCdB0so1KsrZ6TTT
d65HLeqwL8KnBgB/YkJOPUE2VRDB5WvVn4gxrpBMvp29qw9lrhETaX4HuKkd8F1kvE3Wul9N00uT
lm85V13eEg0y66Go0sLGmMdlDecO5/XnQk3nCExYaOfEkcF3zilp9L2j2BUpRs0p5qhzBfSyAnF4
fGKe2Qu2JG06Fl60cX+DqAjER+qC6lw+CwIEnkGc9qoMkrsYZL/trFQ1zRMuiCjjFwXACvYDRkOk
NyqZZPo3/y5jxtoqQaWwdKSfSZcv5YwudzXAux79yRzqnlQ+PS0CIOqt3v1evCNlLms4vj32dkZP
KKQ3qoKfo84Tmo1YwU65Vm2vB8mOrVPTWI03TQSjrT1Xo2gSHE4zJnaXp9cU/NkAPtC/FopqOd+f
cIJJspv3s2CzdQC+VPiNft+b7Cu2Us8K/MwwXzIDWlozSvHx1qdkSt0b40rJbl7R/gSfigP5In7u
7ilauI6GlmvCFn2tx1YEEINk2KbxNRF8hoRDPecyHv0xvPPM1AaW541J8viU7+wrth+TQridIAXb
d+Li24xN86YU5DIuk1o2neZVxgSV8yaObiRw8Dhs3msQ+cyeaGWOtqsa5KCNL/UpPcB85YwE+00l
IOi7fXLMci1hNyttNXgcj85D7sHScbIwo8bKDe2BL6QDwVT2R04c1xhUbG/iyYaqMYQgEhgJK38w
wT66fc3s+0kZCB4dzEWLldPZSRI6RBajNY1g5cFTUwuBth6cEK9YCOFSn0/rS7lKIUv4PcIDJa0/
UKl/9AFlbD6emQLWl6MHLeFEIU5NZzD24PakgByVlgTzKrcweOFFk5pazxxr65GN6j77/xQmPWC4
yZ/AiBWOUIbND3FTiM3PAVGCkL1eqejXbJrYMwVu2ke8MRB02rYCWhrmvndny+CnucfRiRBtWLhr
vkozrVvS+WgFubrq5um4i0PoXIf/USYg8bQKbNpOp4Bcm/jmQlaYQG9PcIUglKAMVvB5gbxGe4L3
z1xJ5IhR87P8HHrj1PtjPhdOLt0JTyNyKwwzcQkOlQdhlCJEZhY2zpJt4CVPzE3/3GQJannauV/C
NRgNAQ+4RfjdaguX89SNaNVTgvig4uM5ui5QVNnzHAY1rHUO2oDsvYlH34SJSXGJu3mJQfjZ/z43
0n68KoTUkupcYvyxX0/AWd0GP/V/4md4tgiePidArllufintSnFvyBjUKveeEu6ZhukaDOzL0tbI
2dIn1bLsdKPp3cKekBsIB8Jyetnq8dbVS99knLROKy567mlwoteSOmDjBNARWL506ifh9AdcVxue
TqJnO096ONWBQzX3DgZeC4Ulp5phDRs6vuHtly2QHkK6OT3pdVxE5XVX391fFgPGxuCgsdkgNu7k
sfP2evZg9s0QM9f3KQrJKLHYWQ1HRhWFT9skZ6HZ/2qJyvpIJtcP5emIdXMDH2qg96tbXLOztK29
DHYn0Gwa5TArvxIYXh6kijK7nd1UHpp3xUGvbrx+O6Js/V3KVaX1LaQEhivqT0/UpqfFTdHYpP3C
MntpE3zxduQ4sTyT6Y9Gmpanolpxv6del8brLzBqZY9Zy7Es5hbVS4fVWG1MLL4tVDoMji7uGAfz
aVaiGW5HlD6RU0uaQ2SVB0d4swlB4r+txVBRs/xZYldY+phcotYR1nyQ4wJF6R6NW0qEKm3jMaDh
Nmh53DKwCyouqVtqNm3efw+FmWYPi22aL1KSfoKMBZQ0nwDI2z9+iTpoVTXLJseHVMUZulc3oumy
zr7BnITcFnIOwSoQUp3m1VmhiwvTxj6kMnSnoi0YxT9s4f4BZHoFrdwNxUZjm2PeHjgYv3KaoNjn
hnPj5cp/5OKY9z915oatPw+l8aKWTvyjtIwenwKygX+hDU2OlCdwhrXnFD5k7y4MeE0Ci8Aq5UZt
iKkFKEE18O16uCU5WRPGfYratBR6BzdpBTRPopeCduWPh+qiZmimGerya6WzJ1ngCFdNfrmtKg+m
eNEtIWJWt68203ETCOJXhLNP9GfrA1t19SMTBfAZSmk9j13gV8lEPUsdoQ6Iv858q60MCeDG5yMt
4eOFNJbchoSWZZLmiiWivitSGs3GTYl7lF1ycthsGiUeFIAi6b43NIjuTwcnR/KTsJEI1UbBnIhk
sFd1CGxq6bym3K6SgaARm1BZ/fl22DjCtJkM4YYqGkLRWjOy4PdFUBiguPKj4NkAomagB2YYtKMp
chsr+eJlKDoETSHN9BwTNSlp8VrxGzOwBm011H2FCVbON3RKyiXPtjhw6cyjjChnVENc9oQWUslA
5iuYdmm5fSDW17CvETn069GJt6QbkKsYZ9OiOSJZO0KfhyXq7Y0YTFxQDX0u79vX+uwwOOfp2fWT
iKFfDA2Hq0+p21KhucS7ZpFlb13VDUsPnrXQXvg7wgYcrsV86A60DkricqbqJWRFgN9Xdzm4IPNY
PikJGFzsYYaUg6maXU5KJKyl7XMQNeyrfdd1mvAVln25YSExtajT9zsBa+N/xsWuPOlzrzIDL8Dz
zI9P8FjKsffcXylYz0Ylm1oi8n6u/GztAxilM48tcc7Wccu/NhhPJHrh7+IEwLHgYHUkvE73POku
vGKc1GmVIlLe0/MH70j0NCms196cLPzEf/6/xktzseY0oK9K2ci7dJuBhx4aIkFnYMN8NWWK/qqc
BWPEAxUr1Sc9XqKTfZ7GkVEPhtfYDe/hLXkiZ/9XM47GkW+eiEqKAlLw8UfIilvDgGpKoqOc04dc
a+NtKAprTMcZkvvetdsg37am2UBJ5NXwEhwO4mcA95Nszb3Mzm5i68OSgO+msY9LPgLgMUi84t+A
phU2adnwxRgH03S6ddEpEU08iQtvpF2II4UD+YuCRoKAFmDLAbBfcmMlPOTdfiWyEhjGDVAyBbcF
DGqOKljxV+buZMwDR/yk0wBbR4tfOOmizuKL7XMSDvYNjzGLCaxkzEPJO2UsYljNp3iitoa8L06b
k+wLGzqR8IRq6lTvRVORvxnQK8XJJQMlGECPAODWntM4Nry/mwyEWQYXq7z/y0N0qyJY8oABrnbb
R/FIRjD2k+NjkTbFmeqqRlUJCuXmLUZ2JFDVG3aQNzvcEuNCEabmDcZ50AAQ0wvQmamDuQFH0FgV
e8y9EI3yIQ+V69VElZfkpPneQn2P+RbwQyA50xxzseW1QkPq6wDsXYmTKWitBMdl3wRB2O/cbzJW
obmByH4ufgPE7Q5FIfmdHWQY1sp4JU262CerB8qo4CYHU+R4WscEVVM0X09r9Cy+LfqwLwQDIlVj
MdjqsgPBxsGPDfHB0E2segOXO1Je1WEHAAnmfGSVwNSPrXd3tPIq9EiidK3dEfa0jHkGV7Otn9/y
GMY2/NcNPTH2pSQ6ZkIAR5jkaaplcckerc9SIf1TkZ5VO6A+eHMzv/0Lki8yNr74SrI80rwZOFvS
dxRad5SI1v5Je6HZ/5M1wdqWZ8qFOb2Msxp7IwxCmgaTZq5zEEFSZFE74QfW6Tef+ptYfYCF5BXc
YJhZt5nxlukDws1O5v+Zo0sgYKxBuOQ4fZPYiqmuG3N2ozyo49kR82USkhsRz/5X68F+UCyhK7sf
O9wGyweDInS3pn3O/81mBPjRt6Pgl5JqcYQ3WWN03KBwsRLN9DB3UjLEY4+FfRP6g1Y7/tQEv6oQ
Bqnp2nQXRTf32MldJZ41mml+0ji2ciR2CtovdoCVfqjWdzVMpMU2CJJmsUKW5mYv/vQFhW5rAh61
y8423vEoBfrh4O7c/W4H+nJsry1/FLcgoxaSfNDRHoWPOIAXO2jPsmxI0tC6F0ePPe45jFfwcKUu
1UuMSUxKMM1jTUtK6NQ3CelZtlOIMBgCVmaOdISdchmpHQ1R5aNtYrdyK8/QV6m6peOrcsdmUU5o
HesKng+R7ehiTOEv1gx+sHLkVlTGyRtcC4jeEzmd2xqxtTJDHm8K5O+4wYVtmbXHDEvDw0HbbuTD
JWeYW1TLSKR7cuzgQ0oC7AL1Om66cVHS+MktKDat39Nh24w2nuN/ae/rI8PT4Db20HeZxRasqd7t
SX0Tbeh9eHqbkRV/u32Tb7mYZ04QrUA5B0077cAU3SmfNddlFTzlb2HaqqqlrZP6spzk8NQY6NdV
od1jPtq/pYYyA1UUwTd+b1WbWL5cdHEO6ZncGzY767+C+q4J7ObOpNi/0tEoeROb/q1gtSOSkFLm
MeB/rC6pavP29qwWD/SPxqVYqJqDeZx8ZebwYpy/vcvuI0L8NYleif086V/e0GRAAMOe9S1GcPV7
3vzDk1e/1w2jwaxqgWe937TQ5FUvh8lUQMI7vu2yxzjOSea6vN0qZAtZP0/T1F9EqYbisNFKBxru
FkShMx456PwaoHiF+c2TtRHSpqVsUBh9GEOWmOTcehdIPNs8wasb0bqNCldwKVxim0lXofJIGYUi
tPDvDGhow4UiitFuqYslryzwWNf/Gp9w3dCXgzRg8mlsSQJmig7thrp2wRpnQGeRvx4KWUWTkLBY
KmQxaZ/4YxHwKDsYy++JPwslOHlQ0QgVIcX35L4JFWTKYJl4PcdYWDSzx4ZN6/tjl3RI3jFfiM39
u+66sFgCfgUmkxKgT+4OHFNgOR2QhYUzpmmk1wWwYzk9O/ct+qxkm7uyNGF9GjmxgU2rtLxqjwWe
hdj3Ie/ABS/15vk3ronWER6rEyqs4y6hlLfLJutXbubDcGmOcpgjoQrACq4lvioK0AdKib1vWg34
OfVDNMp3VA6OFqnUo2ILaU+94mz++gvqUv4k0MonFav+ONRs1av+OdYUo3l4aPATtEBvjU1q2yAA
uexCZpIAobwzJ8JCwMz/y6jBiG7Qr9VtOWT8aJE5n12LGmvqfC3ZM2mWx8/0dekSKqCGFRV9k+i0
feKalMKUGS1PyfwVSd8QvugpwjJFc2lZ+R3oFCMPVbM39J6jJ0n3Rsk3qbOZjMydObb2p44BiJ0g
nDT5iSo34ya08SwIuNSES4dk+cn6cogsymLXQnvxLW3hrFNGUcf1lydv4Shj/c6/mbn35kFFE8Fk
6D66OHaQuDE3/q7aqUAIwmeatUDgKrjMi7nhh+9sTxuSmGuPAanQlC5NJaNTlPnVbyASy1bwRnUH
YV4M3PM56IFDO46g7TLYUJIscubxLEyxqyB6QnvWYlmi8vGTwqs76549pmspZ+jLq1dH397iFPH3
YKZ7jM5a7RSRC8iFSJQBDWuTRE9SDqB55a3MvMB52b4FPGT4+PyXmokvp136Sxt252PHiAOR7h2n
g+IAyAuB75B3DRtHSSWSeK4BpA6dMiqHFh/Aj98XOHSnL0uz/AL1F55t2Xwj1jt9tPQuXmVKCRaV
Z2oeHZz/j77T9lCweCy3/mVBaHHCsvfTu/1DQ0ptChPSGLW1xHw0jPLFItYI+VbibE5r9xDumO1N
bDf68cOHs17wGJOz/t5vaYaqHEoeECxNu6Gq3hqhXHGtQBLw4rB9EziqQ/PF8l6ZIrERB7D2Z9r8
xsFTJ+Ss5h8Ol0gSUA1R+sVoSPpTq5BIW135qGjrHxAE/rakMu44i+luvDX7LepeR3cB72jI4Lgk
AIku5kLIQSbTVePdEx48GLfQMa6UoirMacjVpb33sfOy8NelZz/yuZm6P2WeBd+pRxMEaMiIzeZl
G5Pkr/IIUBsXyTbTCwC+OjfgfuLuJWW6I902LliipkGQZqNskzwH0dFN+sw1umBBoLsCQlyBWSfv
Zaa6AyuGrYwBIgi8+4TWmBtzu+kOGIDaygLdvOtiP+SDYuFgJGvdYsjQRDjk2AN8hxNL0M2pUDcb
5fk2fsytNGNdxaVvc/qJVE3KLbxMtAfqZaJQXsW/EdzoLjr4g3JqRWzM38+6jYOlg5nsM7OToePG
985UTfcGvNQX8vpbBpnfw7XBIVCmsnxFodVDrqtchyCFFNN2KMqbk0gRmxu73LMiAl5SE1tP/7Lf
ihlwOez28vEgK0/M1Vqd0CXy9kkhjBej4GtXGdFOe1216uWbsRja5SFAQ5vcwaYVgq8xGYfbnFdq
oJfmXa70hJXwK5AYtS4z81G/g9UR8cbMmQ/6g48n56Mx3A9zB0ifUA42idwZXOlCAQfm/zkZouSJ
Qg0FE1hIaRGlzAX83FfDIEYuhE7xIEIgLxa6R92qHRQXHXKyfzkRx5oi1Q6BP3pI+KViDZ2UC7TF
AISUXN3B++f4yg8DD3NUOuvUayjctQSnDqgUnI6qo1xS5oursEbuVgCAhi3gIKQT2uazmUQ1fYHL
g4qVDovqMIZHmxVkAXz/mzmjVXY9P+EeW5QvokPxG/5ofgkvfVd0xDGBIvsNbNj4FFkurD2MYU0j
JSPCOgtwQuWMcy4O0ATgZostG+Vy+z32riND+RiXVOkdzKOberDczSXL5MtZW6jP+5gzL0DIG68m
VfvSTBAuLcrNuDwbWWSyg9LgzVwX/b1Ofg6lXYpPlO/fcjO3H/KnOYeJvV97SueTYtLHL9rvro5v
KL/+4fmkL1HStVZ9XSq2lytTt/ApDyC69FR6s1O++IdEVfwEg6kwhA8mkf20QhrUZrHeCjoVaWHx
MujLxglHZTCL/81GHR7JClwiCr4WW6XyfXhzXIQ4X/WL7i5w4gII4cbjlcDGnVXwz6DPlmLDnYOR
dv4sdmeAB96SsOxFaWCkp747PiHOkzBL4ok1AC4CHVI/L6A9ib6BGcVkOpP0sN5/qNmkUUGixBkY
IUKHPrqfBcxOgX8oXxwe/f1EIQN4REo5fVVnTbBRAchd39f9D8Cs4m+nYk0tv6o22qVpiQ81k5tr
VxdQ0N7YCLULt9AN7ymx3uyrixZtK8/l40nhrsETcivtjM05uqSIHkJ/wBQf9pfV9sv+FMKVsl7l
go6W6UlsOVJ10aZSDEa9PFcHNdpOdsH+FX/BAUceVHYvmfsm0tkTHYocr45sOu1MSeHSxO/+IuMo
HMYQbCZ8aVHysVZhPrvyTxHcHihSe8rfcw2eXrM0JIEEebQdq2kixetb0t+mOI0yrLqV5o6egXx+
QpHmaXHjZ5FXBooZf4Kw+gXGw9H7zCoiCaNASEXhXZI5YQWfi7fXSfawplitrHXA43o734TG+6Js
9RIm3+My9SIMJd2BR1iyAbw9N+0B6ShT0oMhzwQyJOdtfD/a2C2dnAFTRWpHqW3TwsPe++u6E2HS
UYf6ESA8xZhpcGC4VT7fL6PFL6cagTyDLcazsyMTRx8jcRbH9E1oR/+qcXY41RAaLIfoUmnh/U3e
A+LOU230f+L8SyR6X1SgiI7DRIRVaFh8HwVtiTsGGBekUxPYY/ZpmVNRu+J/Q/k6A3ZhsmWRtu2P
oOLBHtfx8vrZ66ZFHGdyihUQLjWkGJgj3CpHXkS9WMqXzCuBmIjf98Jq6yMt1ovChkREh/4Rfd86
yq61GSUZ2Xxo1c56GKOOwPqQib5sqq/09H5nk5c/Z73qP2fnZ4dZXqDhq197l79JnzlnB8JG3KQY
sa7BpO7cqKlVnp7qaj5LOJ6jKCNUMgtWz+UqQrYB78+8rqX43tHURecgfSqPPv44Ceq/oyg9lqtY
fhm4MOWu2KEOxKsxhvIDe2NLuOJtgCy3lGAyvA90xVWGBwwsx8a6Iawz8WqLD+z+UygU3SdT+pv1
QcMWoXya/3fO1c7tEs5ahlBnYA5UQAAmfRdyFHwPgYoPzXW8afq0Oao5giGi/4teFFXKtzfVdRrD
MSXEuwvtDGJgc2U4u0pb3A+HPH2H1n6KXrYQHlhLHilaATw2s7niz+jF2amLD/f9j+J0bUcttD09
hYD3+M83DpK1mmdsr25ddd0Hm4wALBsZ5D8p/7/L6DAmXCfyD9Sog46i5ODFVGnMEiPglKmxZq/y
wRV9m4VIaNaZb/MrXwYSke+j3WyJ2TJS5BfNRDtU6UCeg3adhASpVqP+v9A0yn7LJSCk38wKMIo5
j0X2aV27ZnITbSu7rnwE9PuMJ64Rbc3ap7tXnRUT5K3VjtwyIg1c7G1kTA9xOSyZZzeivPVC5SBv
YmTc4c7kASacaELGlGRN2I1pJOehTpa0N+kpDLhDp3UmITCdUfeKcG6whE5DXFv0RGjVA70vjCSV
ddEM6754eJNOONBvEJEe//8hey1UdTg+m4Si3xbJqEya2Juw52cTPXwf+ydaYJv27y5aUUHyLIvF
+6JhnjGmKT4tc/p7j8dWcRp/mAF/7CbSr3OqdSfEXU2Pn8wuCnfNyLtTDua5FvgaoXuZj7JZvypy
j9YuMv6mMntSB4s5FZZyI3WBhFleyzvhIZzusBbmSKK4jaWVe8CWnWo1sy7If0I7jrf8yw7tfgKQ
Io/mHEwXO4lTBrc1JTomB2jkXkHLeU4If3ISzurb4VbHR1qxZKPsdor3O0vltUK2Il6vdcRx35em
972uKZp7mm69/Sa9XtmSdMhPNQH0iF9UwiTO7/xhc79dvxZCIYdzimbwRuorV4/JfFO/r888EvKU
IXf90j1P0wGclfAFLg+rlOorvZdqTLlT+98XhhL0Sa964LID26dkNMS0IiLqb4J57J968j3YyHTt
unFM/WcdzSF7RNvMsnvTiaw4Thx9WqK8gcp/yIIckdXNh0a2InlJ9LhWfwei4QRM946jEptX+6Qx
Gw23z0v235wMdYQzoy9bdgabpoMy7Oqui6TCYq9wUFIkz2gq03NSEUd8U0qKUfAX13tweIXvwL6a
GawS6WQqs54fwoOLnVdMuv/PmfqjM2BzvdPbcO/m9Urc6Q3u7Ix1BNPZIAmv9mgulEJphjOLF7HY
BM6icW3xz/HOFOk4PJycnfcugDS3ii/ILRX2yNmbAVocc2F2gN5sMwB1oNC9bqw0Y0EQb740v6zN
ufNy1XxACdb+sUei0ufz0i1Cwtf2C8hiHPMh/Q4ihNYFTzl3OZiB2jl5/i69xYDElSGxAV9iEfN+
GjjaTCJb7FwVrmSvxS2L+fmcT7fKDS8iUiS4cPzng4Lvd+bmWKrC1jUsd5L9cmg+hEijNTcIJurt
16v5BdsWRQODjrRC4tHXp8jmFXn2hWGmbG//Ylo2jUYxNiVE2pL/7386P87fW6OHb0a8x5Wqb39o
qoT7A3DF/bkmlALJJJi29WCZ+cAkngyq3+jUg/chjIi4uFdaeP9ZzqxhmNRlxHf4b6RmofqAm6bd
Vkr9RKUmuiY9U1cXzL6dudTnZ0zrJVwaWv7O6ySlUk1uVLq50B1Y5ILsDt6XPLu4df2pFn2jBUCj
9cN2PiSM59uTMstjX59gEqW4aLv9hlCF/DKPtQ35tkNGU+0YMzzc1YERywMn6HKOk3Y5paB7WHaW
oq4cwXaYgS7DRVLQzPAN4OthzR5Sw2qfabxt2D0YDHporWcYL6IBHnZDh/FUEEcFg5LlL0m8PjHx
qzWYnYS8LJBoQwWCQJTm3BZpURgFmny+PFYkfdgDPIHOetHufEz83UKyl2At7NsBnKORiSKh2C+a
V95zhX80tvqULxOmrrpmVS/dFwAzBe9JsPPyIiGErvL6a2rXfSLjBrvL8Fee8dwIy1uVseeeBb3N
JIjo4k5Q5c8yr/gTWi7JoVoTvLF3im1hJEO1AI9YFcnx+UFeMGhbijaczuc0U+Wha0oBXif2HAPH
w21Ym1vR8cnTcvpthtjZC6RJiguIY1IWLxnodBn3qde/WrBAAlilV0M7uGOVM6qMV46Zreb7QKoY
1ZsuCuWj+tVKv6Yq02Dr+bBCmI2IIAdHrhXu6tQv4i/UQu1JiiNK0OXL9LdNMomESqyJKW/9iZYY
0Zn5DKwpgQwN2coweT4eNKrscuYwWNw3XPWlxw+6gnPCWQRo946gidIwjGaz0jmcZ2srhbboQfX3
BoV+MvbQ1vk8zA3hzzQqwLutW1/mxddqv7CHOu5uQPMdObRhjSWespTyB7WTE+uhsMqFUMuNsIoM
v2d19oxDlDNt3SQWixkZwTP+B/Eak28umJg8zcPHdKfp1nxPf8+xekenqpcjabQ+VnMIhwXz6ERi
uAtz5qiWsbLTyl29wsPrZZbGDRp2AzQ8w29HsI86zGmTj83pDBEQW+Z+L4tqT6HmXyfXhigTjYWz
pss89dprXqWkl44jMTLZDNWxwvlbx9iFxjG0cG8vRtg4y3H0v5uoJxYQ9rgzg2LD514KOnmKKUHc
k7Wb9JPUh+WqV3ZHynbbe6QhFBwchZIYmWVI1WjKvdYj0u4WvtBZ4/25b76jg7GKf71uNeX6Od0Y
oT7kLwoWVX7sCFvrPTxPN8Y7C1vfftUBEwYM/T6zK9AYuGr8CgQq3jDK8X23aW/05a9ZBKFkzNO3
iGkuYa3KBPFTYryz0Vv6AFOl9OvIRVBgJdKbwsIag2/iJIMurIrQftKHiNK9C2khWRQgAz0PGWG8
BWT590PRsAINpvTqT5Ht0jzpQ5NdCbZxVN6w11/eOHfOAOvwPcHv/NpdH89kwhScG/qeWbcEz22Y
GSqBY8/lZY00ObcSj3hpfdEdRsGngr2m3AA978PPKKXr5tbe1OeywVn8miwIVBMDul2PSsiCvjXZ
IaojsRjOJtUwsqUaRrs0cw/DlAEi7H7ZEvuANhcV6avUad8DTfIkJpK+ySdgkKadQyvraLHgmoRv
XqfCBMUb5c+QIZTFLBbs76/01oQ66B6Ms+wQ/4VCbZwna0hLzenMo6hQCEVSQ2u3J7zFJCeLFt26
awXSXD+4tAwfRg1SGiIsnmCIPxoC8ExOXBn61Jl8xkE+R718xfB3G6U1iQx18OQm1Enk2ZJwy5s8
OPsW99V9MjcsbsVGPcixjUtzTveMG5HQlfAYXFhWHwVCbZ8gzLh4dsBaqV9QFV8K7RUuycOMGLaw
+EFWbiM7QQ9VbHtN5DfBqwML2Qe2mU3sVPHLRRt+g67onsvNUYkbc+tElQnUEVMoegqpuuYAAczv
1F/TAo6L+ZAz+HtGARu2I+NmXfGFb9S7vUQaxs64tlKc7wya9lAm543eQQy2EptAZzAhY1b68751
ybbrFPGBi5zC2Q/cRpplbgMlRPoZIiH9uwYh5CDWiTo9xE3vaRWSczuf3R1Oa7KFe6jZ5dkZldh3
S2zeE5DH+kgS0Meo7H9e9icR0ULN0xkUbbySkghVNP6cNo+FbEwGlC/6sNQOHmAlC8S8lnvdR4Oo
CR8kPIcLhAaDph0XEOqsEgU9SMcSWU2f/yaEl0gqj6tffqbwCGVEIwX/XYRrblm2T3CgPmyD11oW
5UfATxbvAjFOtqh7t6h99nEIXVl+DUFV2tMF93q1f88hRoIjjRH3KJeqLPa7t/j2vQ0Fo0gyp2sn
G1G6c7E4eOT7JJ/lowJJ+9qfWi2iEVJUd2li9cwmC3QpKDM38+ujMSsgWgg0tblCjAjSSfRoeifd
g/4kNxkR7hLMhCs7wsWcnd8dtcUqyRJMDQ+Hj+eFotxBFoXkSVtJE98zWNEe6AtHcQzuWintcl9G
1AmRfWSOMke1ua2P3XWiAy7sZ9Xwld9PX1nyK+G3PXaynEY/sT2n+Un3NwI7c+iSAO56yBa6k/Zi
ThfvapPwFYZarFUw3Dqe2ymXVEm8LJIGxqdumG/fJMU8fJc1Trsil0P+lbKtNpmvULLTUtnuCcGH
22XZk6UhPxW2Pokcc6VQUXtvEEmzU/Y6aPR0MNjpDH2LTBUR4paEtHYhWBoj92g35urNG4AJJHd5
88qi96TM1ZZOnCs7XyXGj8vkI6QzGG284dU9ZAKPZxa+zhmlwi0p1LhkMa/Z7lWvj38eaB5ctHUA
M06dNlB+E342QKHrDJoIeYtvE9Po32sv3M9am/dVijCzU+kVOJ+CmHx3Cal2LU0oS3Kanf6EIxBW
5Mv+a10XIyhEoje9XyCOhUidwP/gT3p3w24/Le5I2Ge4C2OUaHTVkZOIoCzCEiKHGKBIqHImB8AP
RVy+PKcxmgzaF1EpivhPzS7Y5Usu5UgakxCCQdxnM95iQFJ2DDet2NTy6TNOdX+vZBdDtIVqFCDP
kg8d2QqYUNSiA7c83FMxE1ccWgl7C4MzHqaodo/DtEEJKpUC2l5jAUQWd9Koi01nt+a36kYRo+ZD
XBnmTTRypb7VzTat2O8zFEUnK++KwBI5b0a0YdNe1wAzyp2cZ6XBLELIm6nJJKnqF1REUjLWZzsZ
IRntgY3kRhyJMCb+1WToNSL1KOmbqLeOz6HxED2zGvMTYOPWRnVc3vEU0KoIgkLqIfZkslSwlJEI
Cl+iRZiLFItk24UqSYdHIrjAhOVByK52qbqENaCwb3DkMUINs26yXTQV5J5B+Hwe99jALNpeHzJ1
cyyufHMnpbROcMM084+q2tP/3MJ56gRtSxrrathJ9mS/zTPykgPxOnbVDkyUtT/zIASzZ4fYEYRw
/QhEAgGHZYQVWF/98InhHd0V3gJ9dyLrW1YIaHTUpqz+vShDosefwd69rsHUcewP+7bs4or2xt7I
D2uTzXDW0xbQnNuF3xTZTWPCPkcuo+8QUBAzsTWtpp2WrneEXliB4mwk0npj3ZEuimxocNp3OxeY
zyQvVZuZIODhlbOraku5PfrOAgNxveRZwX3HdFl0vSsDfZnb5ZRbu2vje/vvKWI4Y6OJOqvZyklg
W4XbkOIKnDjL9yQ8KYOIMyH41tvKkGhEM+dy5OdbQnR7/Tn8nz/sLjMhuU4d/oy6WT//P6aI4nYl
XGnYyghX3DWcemTPAFmd3zGUTpURWSGNgqzlxnyzsIKrjHiBDUpkldw7/X1jaTXaJW7DHtgXK87m
SEQ2PeM3yzqSdVHaq8dV5nfnXgaIv/87FmZgRQppquJPmTpr/Kv4aJe5RxvgPBSORVepX72WSg6I
u2q5Oey+svx81sR/2Qg1s0KSjASFefP+REXQdcji7ubc+yYcMcuCc5GNwNMfFiQRXsSMAU/TMla8
p3D8RvewZ0GpgVlrJk9Wo8FbHYXGsdLgcMdTAjlgwtxZHHgzS3eLIZUnReku5xDy5CfIYzUMyClh
QgBgj425g/F7WHrAeo9NrIIvCS7fM9KmlqOu+WYHhBbhvaTTB9PoWkXdPVisrhCusFNMBep/Su4Z
fII8oYc8dtCeMEm8sqrF2v0YkdbTDKR38xwiFK7pReJ8NE37Y1VPVkmT/nYFsBkAX1JhKbM4vYhw
naoGRPdecs3J+g7EVfY3WeVEnCJHRY9YyZfnN6b4An3kcFt5x4rJN/cVMrtVtN82eCl6aCkYt+DD
I0nQf5s5BXgX3mxpzILzxWttxZ6GBXnjSz7RicejWriSF/594pRsSxkb2a9loWU1Pv8HFTUHkiod
xjtKhXuYkqfRkwwmZtsa5O1MMkaM0flD3fNfmHpHhKY1v4FiV/tTw/IcG3+lHQ29ig/8wp8bM0OF
T46aykVEcRQwrhcZ61qgl3iwHXhxDOJVgR2TwICOfsr26kDXcLAqVBqk7kq6EPzXM0k9ElC4E728
diu5nyz69FRdJBr4CIfKlF/qSSHQvZnLKzp2nHvmjryH86n6+/u3xQp2jR0RLIJNm5r3tfVQ6HRz
ZDKXufp/CklS3AHNpVeJfBMw28O7qivwXDqWNuG55AtkroAFQNo3euw0XMX9+9FCJ9bFJVOQDV/D
CqHKeFvhkCBsX3zq+HUdp7CXDKYb4BU877ZCtVSXmsqdiqOf/SjUY9qhGQ7R4FlE0ivI/j9H53Iq
dD27R4IvYHpdUGKTtdQLKbWBfjpbh/fGGw8lMddiUYOQ16J9tg47KqlMaNcznXGHATry7nY5Kvx2
H6Hx+hoMiAC1yA4tDZtRy1rWpg6Vk/UKbsl5guBQBGQsOF6Xio8w5Ctq7B/Xp0BeRDVc80pmyHjn
zY+eN3SW+7nrrZ4swc3g3No9u5wJ3B7EC2XfmGLtPEdnfPNMDLDb3xv0oQ4dmkPbb1djo9olEZ0M
Ddg+GVh8S6BAXYIy+wTnkQFwjQzgCucXmxDONmhgkNPlbOTaGGuDRBDhmmH1qRfYwjeBwd+rlcLK
eT7Et4r3tJGyTn2mURgfMCbI7nyIXVshlMbyRUBf6QsVgR1QP1yvhb740cCQqZLXChlBovC3or5C
q/adQnW1GufTyut5yDDTs97OjGtGssuuvK808nNQGgTb7w/rve7Q59sLviCLY4/GGVEmrjJYubOP
MiAYcEoK8LP2AxHLZLOUmy+1hgBMIorvbNKY6i8PJfYqOXnEmjrZt6dkLCpUCnwD5hngq+e6cqik
lCiSAuiuncI8Iqmkk9gkeWN8sG59FP/x5H78eG8daFq2Rhw8f6o9/j2wqGNn8nsBPZLlrdSTjE2S
XYN1WPOCJm3TgJ5WnMU1F9InM8vz2pQbL902QRqN+I1tN9qkT7Y5yRXkfiCa6BqYv35lG0IncXUd
1iVqbCLjACwCjZF/IpjyCidmdJLobrIkVnk/lMICYg0NtLEe4eeVhkOhPyp2xhcRVN4Ku9Y3160N
fi9HVJGVwzzcPCgCoxNvcilghcwFhB575WypOu1iN+D1yFco2QeG/iMEaHvk1rhikV1wuJws3T+m
eN/sczjO6IYHk5yaG6lrU3eWeDffd6uwIm1OuUfmVvpM88cnzp8CH2VNIgtQwLYO22doqtOu5axI
YPXHRg8dxAjgJ4dGKGlgOn33PENCMi7ezRTlaFmEuNokPGY+WdsHvgwmxKI7iz87ZwaoT2jjNgO1
EpI8XMmfMPsDpxFwipuyHxlrhdYxXSxbwjzFGgycw5vls2GPOvphqbrU9qtWJkClxT7lr/UaX6Cb
mtgrosaVLuN/sHG0zlQ+wvIO9P6FbaFu+qlxnvWavEv4nzl/SmBPwYTSvTgaVrY1FxX1eZ+EaXKO
hoR1tKhyZzwrjD4PnZmEy386pYmbZXKdolse0Vxmflzp7CPYDojO20llfMNGRZoxX8JTFSE/ffMD
sc/YfMovKIa/Hg+OeaZ1KZ2GmP+b1gFea1REzIchPis49ppCP9nP8K3QFcHIz2JX3rbUuWaMIdK2
G2V3DWdbkW2vtG4/oodKG6i1QYSF7zrk4mfZvg5joe2hx33gybLTNsYmSFSHGOo4BV7EhVt7s3U1
YKoTmkikC9PPrcDsWSaR0PkU1mI6BYaetaFqlO1H+bthfUpyZWT17MO2wnkoC7Ec/XQdFr9IerHO
+9d2VdC21wLoWHRTfs0TldCIy6QUtHzIwUqc0pZc1DDnCLklv/pF3j6IGTK/zYvBdbs8Z6OIw7EB
jhJpYYG7edE76V5OR0xUsEo+5L2z2ueiAQpyhkj528yPVBjCke+mRj3IaN/dVlMTjFPABIvtsR3x
uO3e9Wao60yi+n+jTjlyTMlcZI9n016JV0J3usqT3X5D4W0Bs5TP9Opm/2KZVChrhpQjI9e9opNL
HOJhCl3LATHya/ktH7Bwl0OJnozWEi559doJ7mOK/iJubYx0gJesZsnAo2rtVGNYGS8upKP37SWa
2RCc/0TpWcsSQbD+so4h5AjRdcNeyTigGM6zC5+vWtLlbn/fRgQILA0Qr2GvVDhLXuQFgx6su5lz
NZuUVWfzaxoDwOfyj6Xjcq3aGXKkywyptgsm6baB1Euj3vOVZI3K1jBv1yOQbnfEOBiknpm78OeO
HG8BwuUdTZJOqz+rju05Z3uauFWINrZvDOGgye7/VNawninsmZDl+nvTWNKbBqPr/jxAzHhTd3Tn
mQdG3UF0/FmQSgwDFEnODp2Hp96ZzHSHriXfqwK9GxgSevW5nm8xEKYEfGggBaqaS7saJIsI4LSC
4tdCvGGaB+6ZzVKYEhzgNH7LvQ6ZLsXXAAaydoLlIve72ZRiWz0AxZkMEW3Lx5/EgswDSNc+rj+A
aYidimh6NHUfDoTQHq0SP73VuX8cYbY6o19GaQ3Jw+hHovn+/boVmXr0mhgjdP3LY+84ibpCJpwg
R6GOQVb4TZZLIHWxkoG8fz5wnxvnprhdsESgpCgsh+la+txoNtqZKvAM9aelrUYh3bxU0Lv6XFh2
2dkjCygS9pFKoMleO07Qja+SyV+8E2fqI8LYTL2C5bx6MzAQY61rlJC83ik3+rCr0n0n4eJpoht0
6q81/5Q5h9jJKoyL318W8UasTjDBRFkM2Bkq70u34IRVm6+bZgX+Eh7UZto2pq2Dp30mKJb10yvW
92ghJYbj1lfMiHDcjEv8m/kcJqTXli9l2RgzfuVy0Yipy/EXAlhNGKhWn3m/0H3O/t/YlOGDDAsc
MJgNv5yXN39epGilK62t4qpjB6Vk3YW3ALSAX9i4nkwDcGIgZT+bZ+qqt6pvOxgu3N6BiEDgEW/1
Dc2rSYz9t+Q+QMnaNfLadOuEK1avnHcKs1hnKGrcNu8mDtjiLCRi1p26GgGmFHX0ylaDQOL4LEGb
lPqnURDMt9HzC1l7LLvvfamM2Vjj3rSRFYq248+7Y1/yld41pMEKEmS3ntCmdNXGYwkoKbnw+x3r
9yLGzg2ImDEsCpd3CqvZW25sRxJHC0UvNt9/ZWBQ5VOb+ZNjFescNkOddSfvYLlw7TGJKiq6tgrI
fZRZViAcItyNLzM+3adtJSmYgNRzeu1g3Bq/DkMDCy20SUKc6uO9X96Tf9mZm/Q3jVNkrnOPyn8i
hiicdm/LEtGxAcANw8lbhO9hUmqSQDnPQnK3btpwBvHYlq42hh8Zxe4SLFfAX12ptZq7c4YRSikw
/nShhbgaMru5VnZo4yF3+o6LYs16CDTOoM3Mp7WkAqzmtoibyVTZ2oyatjhtYeYBWPV1t17Q5//h
gRCIky52oMUxvIOPQ0KB1ydJn7wrjnIj6GZTkjB7DKiK/XALY3ND1QfggyNp/nGX7ft3VE7EzeHd
5oYIonGUQ0c/4aMZP1Z0zyL+4pevpAFd64qBQETB+fJh7Lgvlm4Em4iaMTC80aDpgrQlK6T+TZwo
JhMshA0hV2rLvM4lz78g4yDhQXXtYGHiyWjptpz/IO1zIVdwiOBAHKkPa6msoiucZA2oHR8qCN1W
HlwrvuiYMrVvzV4dFh8oM0XqWGWo6s5i5udHn6gcLoasKG0vSpcUgi5W1kVU8RC39fBzdLkvxfzP
CT86jSyujEIjFQXzW0u54PoUxP6qtWQ6msJKh7TDX7PwzuJ05GTWOmoMmmBFfiqkCXOGMvbwSKXZ
5f0Ec82Cw9B/5YSlq+5U8yv5iL3KcomlA9vG6FBU2WbyGzOjcyRkWOUXYCfeAj+CJxLpUxZxT7Sf
OvvyQwOZAM39dm3kqUtZ1zPpisxCW5VbFQEbAXR+LFYfmuu/DYFqzwHbwZk5vhAu6cJSXfKNPEG7
8sXuhzc+LZfSPiUMjC82DB3S0MyIECrg/L4ES50ftLt3rGZAn2JRna4C6Sp4XsY89NTBss0hyU0h
SffsSJSHklUyGL/s54Rksm2eRaXr/fFuanF99t0vSvhO+49HvSJR2gAvN8zPWeynpG4jl2u3Sm0B
bR+qL2Ivx1fDOd4QQ+J+ROQm+dGs939xi7A3G7Pwi1Yz3N/f39P6vjuj1goWS+92GhJXxxTgligq
GE5de871ASMCSiWQcffFe3LBLYSr+j+ajueNhkUdbquhnn+xHrpkIkqFEQhXQYFJweP1QLLCvme9
xMSvgJ9iwS4BwTsdX2Hel1Bw974Zng+L8yW4ItfA/X1EPFqweoLovtn3oEk+EPi2hRymedln+alr
6QBu5q1SA53aCIVg35s62GdrYctRvvkJCwtZQpTnr2ekrVfWHvWIzUxxTqL4qbXGTARbrwK6ZKJu
n8hwE4epvNojAq987dzdPAHpaJD0Zq68s6DL2DxKYE/aro7jUYgIDYfntm1iqfscvm02+h5kN9Nk
0ZR/+tgA1x+z+XPfEas78+pCXeqH9+hJSa3oOgbloVMUiHyWCsvEE1nHY0TFc3JXkkMDWbY0Gdqx
gHeIHqu7drOMRBQTCF6Nzx5gauOAaqd7oDSvVi7kAh0cYM9symrI7fjuks8O6GUQrHyQVGsH5Xqr
J2zyTvK8patbdPxNkGK7ifHXP2ClyBtzTCVsOSj90D/8KE4SlbbYld8WOxWyTwAqpXGh6X0VeR5v
Mt+muNenb+9MHxw8OR/X5bR9vR7XI8qrxCFQL9ncwJ3KArD81bShhTi1QgXPrMSace9XgS0C8jGE
55swvjsrGxMbX4nBjZqsLUoKPE6gsQHMowzjOl50ffN8mE98otvO4gS+aAaHGUO0hkIxOo0SlldP
uuolNKLdeVORtvoRYYAXADfOnV9btV73JrpLNaBCp9vtouxFU+n7NIJbCrg+DjWiNhxKMderL/V+
Lt8nIghR6Cd1YRasl4FeAqCA65vJ7w6m6POiGlJPNQAWxj6t8+Vjayg//irNGN8u5/HxSCCLrTCX
RJpaF6LqJi0MLzya/e8+gICOljEXiap7cFuSEScP4ol/lJ1ll/3xmsZjt3AbeK0AFDzgHhrSp5zd
Da0YhYUnMLk4kOXBDT+05IK+hZrmqBOEiuoTDWeFHE5oz3fBK0OkGmOiA9ru7IHvopBghhs42SoD
ZIAzbftBQUpXSsGB72y5sYvTRGUXKdZQuMJ+ORBQmNtvnzAkQb9GgN71AgmMN/czsFxUw0chlcoz
RHV5xc7U4nVZ4IfZI+aHL8U+Afs9IgOe8ItIvRDE0yG8yVCkoRhOrfuKwmwuDpzJMGYTWIH44/iU
BpiS6EkgiC1nW69VOdx9iCLQrvyZ/OKQrzwnLrjfERri9Gra1LwnpNKx0m+VUY7m9PTy4NJK5Ukd
Nl490qYP6KdstnmrqYYckBeGfHwLVaOG+cAe6IWlB8iE8xXjqICWNhKnOTTg2VLL11/8fT5gxsnu
ZDbR+uVvH3GxuGDmhEdGGAoD0W/B6gySnIk+1t5o6a62mk/TJky3fi9bWwvWiEBniFtJLaumpbfe
ar17gyJi+PJWz8+RMA/StxxTybYt+jJK/Ye5zt+Xupe7FWTrrNbBrOwcg30xZ+tb8Akq0aV+i1Sg
LOzgmf3znB5uPArJqexTRvnmXkUFKpuanRZN7+msx6W33X2WkKfMoo77dVQpeWklQzGSCTah4DbX
O8E+8j5W8HaYY0GdYoYpFyYFXyv87W27a43cqgolMhBK7R8UA/Fx/Bhpwsirq8WtZackJyR3iCuH
kZfYqNLZzFNenE/RUpw4oTQpHSecEJX/pltOY0UhAnTy3nKnyPL+JOMBFpMywChB2gk+uSVvGHEu
BP53DeTzZ0zZOYvhvWDrSG9UmSNF48n+siLP+bHwg1Wd9NPrmsPmqkYrdZ9bmoTqI7jG6iKgEGtP
qBzNXHiRpJ+YcEwG0hoZCE8xIQKUL5sMAsZNADA8rUshXJeeta4pyQce51uEmMYfRQ1QvyVibjOE
Chqn5/MnTl8MFpm0gJLYxc8WD/R3U5Gg9m1/OahRLbdM2ZwL6y1X7PZt09ek6WoXH3zdcAQoRvsR
mZwa0F/2iKbKkpzMDmnXLf5zebfCPeS78aLymVR4qKZCuIP1TCvboPo7Jint35XwRQ6umKL4154g
6HD8vkjUxc0H9KOD+r121QTiUTFQWK78cNFHcB3Rsg/xw+hg7kW0PWrn09FjL8ywPwdpbF/NBqtp
JsVJAC8b6pezC+5wNc1I8dm/3hRugPak2SLiAuW/dHA5ibE/C6m9D7q8rKmjsmp2s3ftIUz6W1gk
NM7GDo2USrHbPNmu5DBrxGCwhElOTQPBZYFtVbLxPtA4WOWrCRwRgaXsoMm1mNS0ECJE/YzvfeqU
hAaAdXtBsSr1dEMa3c+v3ocj+EgASXpA7svEDRjJWoj2+cGQTkmf9i3OUuYPwijGkvZoYa6lutUp
VI2eMvKYrq6KqtaC4GnTy1J5QJGniVWDzssI92WK/eXbeX1jB9DIJ/9k6Z4/4XoLwHuEtMqhmL/c
D21/95B+QcRqoqhq2MD0aJCvjnvHzVYI9Gl4Y7jMSEexK4ucBqGGdgwuJOOm6nWnLZ+MWG1gVLZC
fVxY4Zr5CFC6z0wjwjmT2rujL50yqoV6FS1at1tJt+m/WKMlVjT3xC6acjMAo/VTAzNRW5hNl+K7
nCCfK79WtzHxOzTXt9HI9v+O5HzunUV0RUV5rQKPdT4XecxeSpaHmEnfpPn8uqzdnDwfjLIjlA6H
+C2Mn0azGmEBi2FluipGDOi9lJ1cSHaUnlMQKR0hlwj/FMxmowO7Wjh75stbG89kChDL7btmM/SK
wTFe25AdCu6dDrAPeRg1E+1yFwYJ9vQSy33g8n4X7hEjq9WT7oOWjLij1k+XALeEUZoV6yjpK5ks
JRugfwu5mK+E3yIQnJdqLCNk6y1TZGvDUIwIZu8edxROOrYwIdcQ66Jo1YLyfiXltziOWz8QoAZT
BLRgeAVxU/ZxVy97+fWKpitZbxyITmM0Cxt6ergcFPnjPVRjT0tOmVNx3y1tukps90QnFiTddWma
ugBMIhGgt1cp1pCgMSXusWBTHPvPt2WVa0BXHarI9S0GHUoS8KaaOyNk0ThyAM+0NRzMVOWn9BO3
yKgzGC5LQXOJ+F68GowaXINzobliWY/dhf231PTj/j6maD/XCVzwpu2ryioat6+CGyaFZJB3ZPW9
cmu4uFrN6Gp1Jeqohu5N256Nr0ovMBPvig8wDni0Yr0tjYZ6VdRkKJmlTtRZ9dRW30hMHoHUZ4X5
AaQxS/CppPsLuqjpslExrBWBldhTBenes0lfAopfa0G6Pv+gbmha40hzVbymUNdLmG/W1RsFE4sz
AFEfv8Ly61bR9yF4NxaH4M05Mz74782qCqMFTNGnobCgzqd2Nh5wUg867IHJKMpODAawTEbtRer8
ek1cze51vMb9vsbtsy2RgcKw6ZroQ3TKUlsIZqzrhhMZn6DOALwogxgyMtLNvsdHtfQAfl2tAl0V
Qm/BYQnFO+JPGOInWn4ZKz5TcFWhJY1U2tYBsf1Ah9LJPi0oeQVfPuYqftVlKGlLKzwo+KBBRkSc
FpA3StE3GHvXfjnZvUbvvtL58wY6senQus0MTOBGEoYuhqTN1jaABslk27+n/7lWXw+rnrh+/I19
jpCs4UY8sfaE2Mt1FOPzfe8r4HaDADuFUXF9qolhyoo1MA7FKlHi1hJ4JACkr9A8536ArpUMeWPX
0xTg7tC/g7wiTBowmpWufdP9pRQcHVq+lNlLuL5Bdry2ueWs1xoV7xvyj2g4997yhBXCU2VsxpdA
6HGYrgleo3DvxosKHsdlf/PLHxDzfrRBu0UVHt1JlbaagmjtJKZnhYl2GHB3+R4UXmvXwd6neIOY
XWMetLQJXh9r3XhhW7FsC0rXIy1Eh19VpwAphK6plvyUc/sUSHobusWqrLcCWCJ0ya991IakrLmk
C0ArT58NwQWll2Wd86zA+umBuiXSRNpI5nctfZfxcfdwh3piI8xLEn+dgLk8vjfjA9gmMgM7yhpZ
fKABNuJ+v+DDzb6d0gO/6dy1l+BjYyuTjZdt8j87D+pGNCHk0rCXbV8hHwfUHnK4VE9aMkzngBo6
skCoj78ajMWnL7bvaIqmr2BX03LATJweN+c3PyoYkPzfGroV+XYjU3fVSKGbih0JsXPQcdStBJb9
MWH4xHYF1+vxZSCWp/SeiHnLUUcJhZ+863pxDSJ9AK1xNVrU/tjanLzXJQSKt0DpOkntMpVsxeYm
WmDDrHMfZmPkNMnmJKWiiJHBEo/2dcgaROJ8vceQcOUdhApY8Rl/PqH0tPL+YE1ZS/sPq56dgK5a
jR3dj+IPBsdmD6KBKDHzFj/W8mYA1HxbcGllUa0ZWh48xLL/8Uxkt+Hw7h/KQKCgddbI+lqrq1JX
MXakRRzzn0ZkuDZyMlKyGIc3YqZ/qiv7idVMbVma+R3icoDy+zDpCAk4Gbn4szeKWPUmS14mEklH
un7+cPWu+JbpqcGu+kNlNGpKxjRxnmMz15XqUouv8QJS5yTLNDXU/IgvrkA2CHuOTfmRSUVP0awd
dQZoQDKsRG55/XtazRSoancjWTL//Drsogriz6YdUmqEwdal4sfHsF/3CnRUlL+VvOOpCXseWljK
/gCG/PveyG1kwDtmyaGEyLTGVcb9yIo9GpxtPOIYe84FMDpZAHfAoMK9JwM+J+IYtA5p8YcFNGvw
9ayhH2HVvSxCekpEXPNUYkvdUSCG4E4Y51lGmcHgY7LsOa8/Qr3btq+rdQNGt38ZwWe2qEb2WZKU
KVWjOfZFPWtGsey89xvsZ8bwHUH2TgfECH/hH0uwQlg6qT2hzQYDqdBBHrXbbZwHCM8mYHjCoYsY
1EPcJm6qK13zLlHfOfmmAUhsgJx2ylRQQ8OkDJlPC34LBCeYouvJOC95lmbvTdzRLZHjNaxSeNlW
jdnQyggDX+4qCs77vlEgDl/N/pgbyWgR94g3oc/U0EiLNMKkwzXJBs5l1psgQW+aZJv2JZ6sxSmO
jcyV/0BrVDB3RIEvRl8q0BJ5uZ0csjEaAbnTq0pzN6cAlYOjEXpm7DROzht4RxoT6r7Lf6eMWBCw
Ti55gzvWReeSX+tRT8kqTVh9EtUqvPfgmz5nHewqCDVUtl3RMG9vVqmN5LYKRAM8HsjsvwVCZWwM
p3lWJI0MR68Ji/xYv0RbfLZjiY1pRuTazvSJQX5LV5+NM+cMjaLmrWtNg914PeLP5eEQXm5IKKmZ
AnrotD3f6vzFQ9Pep0QyjDDxAfz5aqCZySE4GX/Yp4GS8cFJ7GseoZAbs4jW0VMj+bmeA+JCWMmr
1DAlY4zjc/jvmMnv44v0Z5NOaAjSmom9jVKDXQrSrQ86QPP9fxAXJuDQhMKCxQMEp5PyqwJIFbgf
qYeYSdhGgw7yw3llYtlVp1rjS3/gTTTHJ4uqdzZObTtOX9dxLa61AwQRg+KwTGzHHWGKu8WSYSx4
k6YqYkCMiIAyCD9ncccGTv1zRHnjvVcUrcr3ISeZBOdnt2F5HwW7baS/Wr/nTqBco1cpgWsjO4Lz
bzQBncJ9XqoZlRvRB5RG6zBh4S6vo9rcQZly/zmra2rHvuMHIyWNdSLUlSmDVBWIzaOqs6j2c8C2
H5hpm3m6ZVen2WZjS3jRLn25/1yGJvwJuvU0fyc8sGIjzQkloz4f7ShovK5VDnawuGFNkOvqntca
+GtohC8WrBrt8JckzSODBZkIBx9zlWG0K1XF1cnwQzqYYxy5X+U2YqfMry0qHETZjdxRuVHhdZ3t
ea3MJHvOyRZl757cztFdgDq1HXyZtP9x+xAQAdg2+6PDbLvIgX4Ya4uWbPfc9MJnCtXAsVpMy8eA
eluzgTt+mpE+A/bLtcXY4DxtK2uZ/EMJblGA0YF+Sp5k+gJpRFey9dkcokjJxZj4w2DmKkTXJSQT
cahJEyUDApsl6yCN8wUM2oO7W0/Zha+RMifxhwcha9TnJwTFNUwJbips5dTVTk794wIpa/ErhE9z
ZCODOV8HjW0snpgu9Fy4zuRRkwEq5gGNQc3caQn3A+5Jxkcc4ENnmye2JjL3ymuLPnNsLyRqhuQM
9TCeJJyLSTKv0SdqnTqW5rkyiHlMtyKC/3z8BLAk632sZtw5OSfpjP7iPBp9BBkyWTEzzXmT8aIs
D/2dIsfYko40c8GRimgi7o6+9MmsYrXxXqltq+iuE+Q4e2p+XudIRTq8hntTI6oaCXdI3zo2xiZe
J0gq2Bob/VigZkW9oj5y26PwveUJ+9gVAxJBMIPtuORaxm98FdDtCmS06LQswDC4wpjBybaay7QO
6RpkG5YOHVxQhbeKC2dCyhs0p0FbroM5ubynf+dzGgSGlFmAKaeMzUzWOj617qUFFsVeWtW6unvb
De/8Z43x9RNPzuCJHpvUGh+1UuJ661Nscu0CeHzvD9ZPUv4HYicgzFoQnfxQA/6+ldTAFA0wRdTg
b14cL/docD8/3xR7BXSL/bTMRTCnr7iicqUVJNMaIyY8CEdpo5MD6RKuH8s4eeK8wdK4Dx7+rLmn
JDT4WL24VAoTRdeBnilcdA7xkkiFagoEXH+PxpkuUJNh+of7neBrpskZ9C1d5AK9D1kRtNt0tkjY
C0lxUUfnoj5YnFj9f34qnCUBhAGm2hNAtTeF3Ys8O4bdfZrFcZ101cvZzMDfs/EiK6X5QX1PqdOn
17ElMjkyvZg9nDtjSn3SsBzEU44DGldfqtahXbNKvjOzoy/gzb2uyU5iE+vbI67rakmol2p9lmHZ
MBX4rW6YsYSfQc9XnWoXUsAu0+wdhhpGFXD6TtZLioefFQBJ5A31wvbwv6nM01z0GQ/btSZ7vNSi
lNuz/ivLrvRoB5S3Jtsyp228S99KyNbojsJ5+eyjL06dzaxqjZbpl7caYXWIzqkSLFGHlw1PvQRi
52Q9sPZyz/WM4P4Rau+jJTLYpedDlpN8dFNZGDq8d7+RhkZj0MEoZOIGjWUXpkx65iED0H4yDX0b
Exg8BzfHn9qW2++nqyRsApmnae9xoy0VbsneGrMjO4CMYAKFqQVrdXddpZHu0OV+RHV7MWY7fIH/
6StpPzK4zr/Yh4GOdj3rS03VcS9Mtl0VJqpU6717IrGN2Y9dgCLq9MsXDcUjoc/ofqAFq5lX4v9o
5osooAn4R1eLjamaMIOowKYMTWuGaBIgZ5CEmUww7ery/o/ri4C3lmd9Yvi2KAIS+dggIB7N/rXh
zBkaaTQY0F47BGCPcmunIs7xEnjCKKpHZdup2HDoHOVQ1w/KAaeLcaxZDyGwOmPw5ESEyAeGf7XR
H3y1qvSl6Hxp+lP6TU5F00SYMuTvpORji/8XaBzIZmEQSCV9ngjBIA4YI4X+FWSMJB+7U70JNKuX
MQuhThF6qMaU+D3tzZYxS8/9sA0hH8Wx0lmJyC3q/GeHoT0/qCW3tAxzR63Mhd56UrbFR9GB0Ixd
Od3rxUsC7ugXrUvEt6/OPKE0DmB2o60F3LPsL1bl4U58KeaaFAZeHBZ9363jIkf3VT0YVkp1iqVO
IYwnQIOaax3P40OroJNbSVvUMw8e97Y2aw5Ff/vEcRRcCxDMIZZyjp581FB6WNKjrNdP2n9XpB81
jHHgZEE5Vr7gCxETUtzv/OE+xkwArwvxDwUnS+p4OPV450fiDac6O/fwnkCA5lFEgswPGzM/JHhI
/uwnpoeMMYpWSwQVJxhJujOvV/SQATuq+jsztedssVFWLPGcfBMOidtjApMFdiQsW8d4WPv3yxJJ
EtfHzcGGp5c+GK5R3KakftzUeICZz4Cug2rCpW3uIdAiRi+uCNro71qcG2pwJd6GghaabU82wOyr
RkWW+Htd/St55EgdfxDgMWxV4tEim+CdOVNvRz3bsdWXtQUQYq8aVxNohi+2WeLnMc1/pEF94/UA
80BMayUH2YLhuCWoKe89hlAUCvP66xNz91rY/kt/UvTMdjIcDyLoZjM+xqod9nvK0hBGIZe6JdAS
A12LaWaOuyEXlkFHHyD4CyI3/GPP/boXAP/Fqxput9QCacqOA7H8q3TDf1itlZ8jJ71XsGdJbhfm
WLSHW2gwIO8MLJEC3fgCp/lVElnn07oQKodkC5ADSE7Pk3lA2s16ubDlMo7jlEdRnaDHLYw/OxUj
qRqwsIzRwJUwYS+1eikqt3X4tFtn2dqR1zXoUF5tZLGR/H03kb54MlpJ19We/Zd2lCp418mh9J1Y
D0po3iNm9zw4HDK+NRD2hQBPGyj+8QYjRyL6gy0dZyCfPs33SZNLaWx4G7wisk6F+1wVxKuhcI+c
7WY4XwSUcN5U5iXMqCy5rH+TKp7nIKIv3m2YC7WK+xC+QdE/lZvFT/I7vuZGA/PaEzk+YdqHfqjU
kBnBQDmvMiVbxgd1m7CMkN6B2U+NqLROmyOcbs9voq8Tb+Mjgw5qgYo/dfvZxrWnwZEQ9sRDDIAM
miIBEQU34vesq5IUwvMpzh0Th9L8Unj+v99mpLSQMG5vC6BR05Mmc+QPhOBkMhPv0FDg6g9EeHag
CniokT6gkIlM4LzfFkYRt+FZQdfQ31TGOjEs2E6o3HxgiS9P1SqSU0355IXEx72joQfjNMkHpEYO
In6HFERTQPZZCePDF7Fnx716BThurzUDSHKwAdWhGjKP3RMUnmLfxbZXotKXjvEdz8USBGA5Nxwr
nwdFJMs+9EbYeuSxXCQQREks0sKPjhVXFw234FXZWlbcUmn4E+Tv0gubbYeVRVuZD0yFs9fEmGw+
5SMG0GuYTxgdCslhTW2nHgMMOdK+A0sF2MnDB5faIjs5bzbVhDn2dwp/XIByGpQN3gsEe78EMz5D
T2QmK4gfQeLoJZn1P1SeaihKPBPZf4zXdUu2eFdoY6yovhGjT358Cqkm6t4sfikHpDg2aCfaCzZ/
pHtu72cqkitICdNCM4nfgtojYzM092rVKrn469ewIASyuQo6I+JydW6aOzEQFJAEeO4UouRpi4bx
7W/G4cbSeBvsg2tgD83k29KDEf83xPeKeHvd6B4Gr/fhvpYtzQELZrriiL7xgjr8upgr+vR8P+lD
9053xNiuN8+pZIgFPut2Em01S/VV9F9o0hOY/848wo7gKHFi1GS22apJwzmD3avaszyHA/0xiKjm
cz7CPmBJgzm/EQj4KPNdffENtJ8r+bMKkF5oNV4rQlBoCVghHlEeDi8r1IuAd7RDudRfMdB7LeVb
iD+m4WCX5eRCyqC62fdlH/rLfFwgDjCHSOxQNHYAP1gs4mpd/2qm6UkTypp/cLeEu9y7Dq7uSSpa
49CsxwX92FYbUwE3iDlTNRQUlDBN7sAFsOmFea7RDPpmxjg+Xc975KAPtyU1iXhrrFA4vwzpYptC
2SqEBM6z6yuXUeHpByYnp/yqljCISnjkM7S54gBxgZpWdyAJxXIP7G+m7ltI7ytmk0UISitwZVZv
NwIygXguWV4OIbaS1it0gzxKHchVSKcnofBZLpGTnptyLdcXL59peO+yiPQts50+aD16wMwnu3Cr
9ZYvInc7swgq6vh0YR7z+nkXxlVwIvlJfI4RzBMpKVl0TMDTJ3+b4v1tJRGGyQX7LXE7nTCSfLJd
MzBLFcqPqhfcs9MvktgwANCFwguF6zUecX9H5BL9Y7xW0ULtcfOdIOTSY0KuxZB1mZXl50rOdSTE
qhVwfxdBOMGu3Sd/AitVljllNfBorui41+5iyB5TBpT6E/Ms0MScrVdZkoIas+cKeOuedkyBIh9G
rZv+53TOXtI0qpiRheJuRaskWSWRbJDXbjtwV3lvaAUGrSmhJavDWMvd3IDfOPRUdNjHWFRhqqaT
p5rC1h217q+Gc4ffmqi9Id18gx7zgr6JQZpHhDxmS9wSZTETa912hZy0np0Fs8CliqaA4vZFdJaB
sx32IUA46unf5EEv9yIvLpDEl5xRvVES+3AaQmUQUSSIemeLqHqyGIk2bgcL6apMwglrlYEsV69B
uxBgCUpomdPgtyuDmRV0qzLBod2T5VuSJy+D5HORiKks0jdfPtxsrxm735ivp2fkl1oX8urvlXe3
NgNABXfvjzx4NheSD6XFGs4SynmPw1PgJ9rRAvRfruH6ltan/2L4N24RninHHWRa8mc2Jfoqjpng
NAHQueF0xGcv2u9JnK7hzKT73EGRbb+0EZa0Kiw3g7eKhmeMW7ppQtW6ke3CJ87p38RVlfSjVK2W
cqgKpmNY3ZhKhItC+IgxDycsYuPYDBFO+AAYlj2eSszYgi3LliSlakAbR0EXucDoX1MSS23LwWFe
sqhyA/vwLI45222/Y05MnyVxFtHTPm5iZH/yYNt+fZtAV6RxYtx3YsYuqOcfscsx0gYg8yuXzVQ4
pQ8a5DmsJNZXfsySTJ3vyGPB3KZyEM9xnbijS2zH9bsPotdrLV3MxfC2vdr+vlVnSEfl5T88Yqaw
6yBEBvmLnwm7LJJ2OJQjwq9BUCf6S68dvpqy0x7dBoRt1qdRuHTaex7w1VgfztiGz9sG2g/UACqY
0+EJLFdcDJDO7ZI28ovGe1RE9AfmzFLDV+DOMsr/E4YaA8hdcp8CrkfAgtaceF6SD9yc7yHZgzG4
rHgeeHJwhJwXg80KLy+7CDuN/cbC2gV8Sax3UgcvM86VD4Ml/rC2hPioibJ83AVqspgJXt2coqtH
/Tp+bHDrNk2pTKtJSwKvZWJRISy7pfrvD1gnqwXFIbNtoly3QHsXdvktjacFtsLPZYXxLtcgwKpO
/lORPjag5w2isPGBKI8veNKKSNhL0+3Lq9j3uvlUZXJ2faur6MNgq9+pWgvORgjygxpiMzAFiXjE
nmJOedzr8M5HYmIHyp+AU3y/D5t8DOqHVatGXjbF4Rxv60s3QPO8MHgKNzv3sjQoEKMBGoxdQ/Fd
16+iqBejeSR70ZM2euFwGZt6uwwDpN5ljTYMLm4Ftu7E/LMtGewXeGFwIacjnzTj/uum+pKH5Me4
nmSD4Uwd8G+c2sWfuuARRMpgs0Z7cg1YKR6WdMOCeaJ9zwmrMTYz5g6k3zqgWJ7T2siTTqR2L0KN
Chv9YLMTNM3Hy4o7lTA+F84tKZem8Ql73FdKUHLKT/NCKirrNmt8DNB/w+f/DreFhyag0CMmcon/
XNCN5Rigm//3kpZzIGQ6CYPvYT3rZJskLNbfxvtp4b3HX1k02YJrdbQ9bBKkvH9zVvmjE50aP9Tr
GbLvPRNt5fWMDSeVbS2uDVJ4UiwFblWtHYAw/8p5sVAh4wM6fhUFIeN8u4SqZdjcdDxJmjb6LVXp
qvtwqtJXjgNlI8s3WTUF8HyYYaWR6g4XpBAvkV3nuEdYlZWmKihE7XvFEBMOonsQ/poJVUhlKj4O
Gk6QiFxTt+xNE+J4R2xIPIkfdTv0UoO9NZ8ApnWgZDhL3u/xzWWVpmrqMs64koKiq2cVWmuG5+ON
Nnzzvgn+sdC8TCveQvI8gBseQDv2o7tDQCzd+e3i+U4GugBv45fwPfPYTng+Cuhb4vaEIXj5R5qR
miN8uVBcrFHr10jbwiiN3/8miJ0Uq9+d8OUteNbepoQvn85/OP2izfk3gFBVVGLH0zsDwcn58kWy
utcc4pi7WJMwpH+MrgDzJlegpXL+UzZbttRVL++m1+KF0MpiforAbjgJHzPyQRRjxznorqqueqtA
/VhNyuytky5Jl5TtD0KCOkN5MUE3rHrzhqBC3sDW3tPiI/KXq6cCYll2hUfDrepltTFZCQsDWF4i
eZA5eQV4LK3TLlsEMwKpgzQa3dQ31RGKBH2LSI5vnsM/rJ082RTipcBS00dMgEi5sf1xK1qn/wPD
AB1ooYfzV0Q/f1M5Bw62b/2J++VAjhnkIGnhIu1leqSQbQr+mDOZ07QKkZm+8gXe4JKsx/W2vPKP
lOr/q+n+zOCIJsVuXmyv+TLvXvxFIFKjr1dDebnXoW1NaU+GzMzxrVRPns6dURt9g+FDoNLos5zb
DWbAkWcCmq0UxGtXNaQusVMHzMQppz66nYX8xdry8oY8b02UNiNMF+GQmmtfUQmVSYZ+dkVluVO7
ms3Msuv6QRrQgNbWkoMg4Pp3NKEhUUO8zquQNUTnodZTPH9SjPlgmOtibMibWNB2T+iIodL5Scdc
BIjatFkpDhZzxq5NsQ3kVe5jw8I56pFZ0e/YbO9mhYlLIvJQtE+h3hqQFI5el/BbuuFvIrrDgpkH
TgOTsfLpGtWeX8I0vFpGuqw5+I3Ov3dTDBkdcuJFAc0TJI+RUhtZpZ3wKpr7RfcfjQws/QrWuSfZ
Jzeegsadj0DggK4SqHLdel3tsehWGUfqf+W8p+i6ep9ClDyJuGT+EvQ/79hmnrJCEo824pwH8DTJ
YQreDOFOSpnzzrIg/CvAlD1hTkoOZLym3+R7PJO+0RIq/9MUaBtZDT9/e81DqIQ30leNg5eyhD1p
U5kT1RFXDX6ddYcVvHPTyYENn2iU5LnDhTRvd/opGOPJ2K8nDQA3m61YOnNIcrjRHWqwPEwVole9
nfi6I7aKptHZWwtDTpGM+L478ZPFcvlG8qAsQwnb5197p65+FpkJlUeabFrsSTrDUbjMIsrDUfJE
icqwDpV5Xku401s9erlfQSmnSbXnbneXEL71qyQvSgAfUbZabjS0px9xrp99X5XyQ+DMjaJhN139
EtG9dxo84oTI93sLg147PM4NmjhFu2n9ScGEJnuKyjc9oVLRmqqQDK3GN25jhNNVlHiONhOCQwoJ
gYdBFhxLpXfIiRO2XTECcGkbaAC/QqllgilRUu3bPFp+iQ6J8kiXUtDro3vIJSdat/UiRTz1C/y5
3fSUx2NMTk6rXVTli81MPgYij3xN7Z73ZsnEPX6ysuoGsXCYrGXOV7F0McA2ZeiHBLejxr5Vk6M0
C3+DnoZ6t6N3eHJYtWsrW0GlCofUAvIaRdgNvBLfKwNBpQZmvnBZe9Obj6Xq8Es/NSIVgBJ+GF6R
pqtwiEFuquMLgUdu3f6wV2j1bAvYMgKRNYFHa1LBWJP2EnwNhYG9esLEMBcbSkz5XtvFHWCZRVLE
H6B0Yh9S0k+K5jbccis2nvWp4Pky0D4PhsiPz0BzBJ0hPBtojT0n2eUrnR1+rumny6cZGzr5w1pW
l9oyJ+oDsbhDoXADC9vQg9P72B2O82GB0lA13/2BFKSVL0/2j5eIkUQb4v73WWJmpr+M8uYDHgkB
tNl+TOEl9uOXHPULaORxBYgSOjWwBDVM1IHWk4Cog6RsqK2PsLEXe3enuUHvOkNe6xIh4aOL8/+x
SJ+5Q9FsoVuKyUnhTvNuXvtrGaRrjWipW4QEsQHw11umS6CNN/Iraed1YB2BFFfSRIdmdt9y91Vp
96uv4laR/B15cvIo3zAl0I4bq5/1/LBe/vRybKdS7ilzYAkI+t/mTkb0RDM1KBB4wrp07z+HOTwk
JpW0ZXCse71fLxAXAFCwyac81k/yJ2o5rqhGcZXZ5Yj4mId+UqX9BA/tEZtxoen+qayNsNP9wjdn
73N3COhqTJ2EEk2Z2P1r5LxbhzPytpHrNIVBbRLYJe8a6iZES5M3AmhncdPBlH3pxBdlmm/lJiWM
fjfg6bioy4ACbe3Hf1feFkOKjLtlHBE4g7E3Oje5P6ReSlCObW4IruTt12apcRFQIOzd3JdSveoV
TyMO7PRTeevEYTv1zJHa0+5INj+sYZ7feD4lfIr/FKG3d21TzlrFu6rnV2JRJExLzJ3EW9BBIBN7
GdX1NQyT7GCWx5FpErKE5Yv163DTMYZPcOo8rtly9sSl+HQd2NpdaaPRK/Jd+8evlhypPYkvXISP
XTK7Nd7026TlKD1YT//r8CGNDS/B2/kryUWUXhiJy4jrJzuPOfhzoCkOFXfbK5gjb/JDKzCV1nxH
CVoBTZtdi2HyJjbuj8Iw1XSGA4fUzTMCwJ39tFTdHEdO6/3IKU5Hc7bMsd2JsmlODknnM5/dG3XR
7iwN+M/v7RDZdbGaHkVLe6evjlvj/QIPMsdlm2YaVRI4S2BhqiwFT6p2gGaGrOFth1RWFdsAYs10
WMTUrvdy+sU9C74jcnhZ268B/XTyZzUJkLo/DrubpTcaKZ8++HZGhnX4omV7EzogYiVZMbHfPgYa
/kgJdYPUhZIfLId7CoRY88LDcndT+0irVm/2YXeNZye4/G3wJOf2fLrBMrDcKu0bR3Kmh3B8Ml5n
oVQTkYsa6WTFR5thUsoZWa86UiwJk9/zcBip6QZb0R2cviBHMf3uAVKg6e7kuzhlO5AHSTMeGaDY
07sPTBk0kThEHzLwlE/0CtMzsEb87VHzuSX4TvEBgDkLem2a644K/v2DoJ6DHpKWGFDrrk+ow9LG
EW2a4O4/QZGp0w/oN1U07Mnw5Y3YlYcQZNvA21TIeR16z0P39ECJ8qH8u8e2TYX3GYzVAprpco6z
TX+RBzRRPGy6Se/Z4UQKzciKqI+3/ckt9fVU3r4phpoDxjwL+sHk/gX5oz1uRmO7iUXTBl9FZTjy
QMRE2vBl0IA5TZI63IS+K+i0n0oYr41Jn+HIxogEkzMLOaowGe3WgiVSK1QA8uNT9NDiudBlCFXO
RfczxX5Bkk6Wf354j+RwqT06fyDWcLcxAkf6IFrBgfZOT0qD99SGrGchXg3u+OYwSiAX0BZx1/2g
tPT9X0sF2ozmfig9aZ43Ns9pd4D0b/nH8peujvA5xBtLSdsrmyyEtVUtf2/g82uxB4HMkf7JCEBJ
b/iaILFPvUih2MT10vIohRF1uxv3/xVIWMBvRtWyfyf/kBZ1x/FlldUXq0NrrMtGY6YtHviYU0DL
mDYUfHBSvE+e2WvjIe9o+J3qwFFY0i0O8jVd8156cRnPH7pEaMOj6bL2c2Cw1gA1OjB03jMVfhm9
LNMhvuH9c4eKtN2pO1keHBddPjWAE4USNwV3mxkqieHt5U/Ssz1603hyS2DLbsKE1gM06fYElFZN
n52bzUIrWZs7fP01qcxLJz24h/wTN3+vwgSWkg77gIc5MyR3ycvSEkCUJRK+Ae3peEtkhOJem3Yu
m9LAUQ93C7fPhV3+JWd/lo2tvnfo97gF++FK/4Wb39SA1d8ciZF+EbPFfZYLfL8zT28vU99qu78n
RkC8loP9WFRFJddQXi2RkG4vVOlI/XnStREvHhmJtwD0mh7EeS1U35Kav+193J55mR3RJF55uE7j
v/UaxqFpltI2Ta0u4gyKMlY+heyjZnP/SpFqmWV/sHofKzJ0ahIEmhOIFvs84BkTQqmgMWZD30hW
dJUdv61Jt8beHpXQszqYsLsuwsiq8jvorntQwo71xMj2Qx9ThadOgp7Dt+dZj2Sq8YhPmdintTKI
Gj/hyBV7+1FYT7qhI76/16tP2tBWSP92H+WpfptHA8fIIPrMFWQN1iHBbaz59bdb0kL1p5liUu02
vHNTIRjp42zobbSKO9G8Gs2GUj+55nO/Pbfq5a0d2/cBRVqi3A/Fn2J4C1qKCQx6ZdC0772rA+Km
/eSNNYZIfGJIV0rSzsBLVy0RcFTgZIAhXis71RRmJ82+FuMXsdYvtoSpGjameHds1DdclwN9eby0
HsVcV8aaXrjJcNdRhgk/nzdri0w5KgbW7+BKohus4j0WQCv1IiBSs9zM/iFgIkpcgOsbw84A+1HZ
UQDUHPcWwNhiHMhaSFsJZaUn3BezpqX0c+qxAxJrurPZZkNA1mcMvqVC/hAHntierWaPnnN1RcKj
OwsoJLOIE/hh7mZbAxZ/dGgKGOBxLZbkyCQIjDPT82H+RzAjUTyK+ekkX6A8hrQ0/WUGrLkqxMLQ
T8JZZiPaQJI8B+tpqX+wAAqSLORrloOYHOGxQoa+X18MJ6RmYpWIQpGZzZnBdIp9OeLEqR5ovZqO
Kk1Vw7YKS648v+7Cckh2DpS+slFZLHxhAzt0CJsYCHMYjG+f0J/BeYZSngJyhuKTO38ueee8TAxC
fW8BwtbWsyUfITAoKzTSmmP/U4g20XpjjW/MhUPpsTgh2q4qHOVT+yNiohe3+2gr9o5qR0keKNXm
p+zihVDfH9hGc97FC1DbQ+3F9kkO+f1JMEpy543ny27oIvkhTX/O0CA++J5o08lmEwNRzm/tuk/Z
Hb8SvmPnRgxPob882FrZSQxdCIcMpBfN1SjlvSbPZadVW80Z66Hbd2Ptxf9JicKwhL7ZPY/PrNuD
5G3v3MoNii261yAUai2zdTexrqkjWsccPMcxdkdgdlXG9itKsoYI7f4eDS87nRRIR9ozgb7o2jEk
RMTWvOwR7ZWFgX4CfNRgpP46g4Z8yh5zc2SKljq+gRGDjs+u1OB1q+4b3mXI57ukJ4ruQPqqEoJs
+IQwGHxnAl1klBpvy8zMraDVJMefnjBhSVbtXM8TXd3gEP4wPmuFXa47setWarycHkEIjZENU6/7
hMHoeECVWarNzm7+yh9UWys/a7FKNsNG7uCvGSo4kozOD+7eSMDChVf8KyE25FIdgeX33kxCh0zX
dSc/pmETbO4U8rtZlDsywWtlrFrNWW18ZWOkrZ9eltrB7XOroOxFsqc90LiWOZG93mXCs5nrxzy5
ycuNN9UYRHeZRhszi64PL1STX/cfxYgUeRHMbr8yGa8bUePkFDL/dIz1Uf4a2omjpAmFeqN8wl1q
L5YerTacPunf5FeKSFdJD6os3Kk/Pq49vdf5JV9vgeH7TF2XOuTgMwZdqBvkPwpM8bTJYJSLSse6
qCJYs5wk5PkBdZ8BVY6YV1+L+1M77jQSYRcxUXMdSLwljNEa9e7Ymi2YY5kthFI2P89zk2qWFtpp
ZflZbiKAz/9AkHGyvIO7UoqNnGV2gqDLS4Vi+Hx8eT4jeXDgcrrZ0mcX6rPzaOatWj+aJIRmjziR
YjUF/ItKIRZG5oSS7hsiLZbyeeErKXM1G89qeJ/yeE4Q5ds4mEc2btrPaJzSWQJ14zr6mfzDpp2F
Trzf9+gjh7YI+z9XheW427S9LizXE+EKC544OhearsiQJEiqxVvakuOcOH9W2lz41S9gD8pVsD/9
DIQQxWW9LV+nrdpiQr8+B88NYHDndh/slbPkWGgkb9kAkPg34SjM2wOkbPpwD1z90PuDVQE1gomr
CwwCOeMJYRAkassrlSoUXPwCdyoqaFHKUmb1v96u8tBckBRPctu46WnYHLB1lCIdyDfV7WC743AM
x6093fA6M4wpV8JfeF0baffME04oKo+G7HXrZjen2yPOEwyT2RC9HQMceemyXha7xgGYhAVqu4DR
Bu4gizcBr9BnqDAUB5LaACWbzVqhrASMCgLEkbtYmXle90KzofsBY3j2SB7/XSostoW/raPvB6A/
UmGeWEZqn3jzgLt2OB7YakVafs2/MkEmKBkm/ThjcAxQ0QwgRlC/utoLnrd2qfTayPUUZM+JJK9q
w5IcvwssqYB2q/8AmrRx6vUUqMgb6540e5l84ecYwjwNj4at9KnmfUBOY2+8puPZ6DKJzav7zASy
M7RUKKFGKqSd15ttsPbP92tJ0LOvg+SUeGAZGUBo/OvGbyyo8t3nOPofJcPtugbTreLSeDRBLiu/
4SaaepFv7mcH4euI5iBBf24NvOdjDyTdcbJcvg7O0EZ1WrgmeHdEq31x3bQR96GR/FPFrqE8Py4C
M9L3qKl0G7QdEZlKY89RCofqniI+slZdCGPK++KcOq21QPFNCJDZnVuK2wbaloAysJyJs2FR/alY
Osk80Mu3D/xOJV1vWptDgL2db7koyeL1Fpde5/LK/8//QvSeYB2M6i/BOU7ijTAFoRKqBg0hffzO
ZATeYr/LtdpCEGbO+8Uw7eYzbfPncnyywuwERWOaq8htiIhya1tMGPnSt+glWSaL1TBYCA17C0Oo
QJVLUBxE/euHZJmmvQcxUCF80+9nFtM8+tJGWn4lUMTDDgdua3HTpU06WYPFpUYDPMljRJlyawXK
rKNdj9gJTP4laPzqIpRebAsTn+vQ6BfhLIFzlPuWrdylele5UT+VqfAPgxWQ1TiDMyw+3YtYX1iK
8fQWHvHz3scibCoe+HY9ZY13Sv9B1UBLBMXvpD8oqTYzj5cqEuTi/rawh2uzUTbyaxRke9iAt5tC
kVVdcfWxhCdDB4O+5op52PH12XEW+W+/+bldwhaDWu0FSolA2ck5IcBihOEZpqHlxi3GcyH6Rs0P
Obf7msI3/Mrj63s+sOl1PT8RGhWriF8xQwjukWUNRq0FNYPhA6/3bSec5jXO7S4K5aQJJvbKRyzE
RKToRnjgwn49u2o6xfldgKYLawQl9j8MpaFChoDfN9XJVqchyGzKJyJhX5dsxdsEvpcmgNhZupmb
K+KgJCu1BUuy5pcWbk8VfRVzEObYn3gI/PSrVJKtipAmfWkoebOHUPZnWlRn9cX/I6AfTDVIhSaL
Uh4XQydrb3iFNdG6e/06RiZ1M3YiOF41JOHdMzurt2Q72xY5oywu6K8+YYDpagQ/q78my0C9cTZ2
wwDHI5vwWp8/5aWd2pnMT3pVye1Shk1LqG/f3yKPMMAhW9oj9vG94RLZ2KqXI4e025wIpT0jBnAh
I/pHAJgL4OBIpuCMywxrdkeW48rW/l+eidwRSCgNv36Rukh6oRtCxqofAkQt6PRYYrUlbt1u97QX
yt/QsdM64qQNKRiSAbZAlXPZSNyn/A6DDtXlXmLCEwTYkIfWMn5TmAscQUjJreQpnJvddDDd2ntf
CLGsgNhvcSn/SV8sUUdEG+Z6qiKZTp/nsI5+dH22cTl7O0X6jb42xDyYkF1FW2Vn2M/mx9UsH4Qi
XsD6z9/TslWxQLNlfa0kK7SwnP97jq0M9IUQ5oe77KKkfwDAna+U2YzYP3n+IqhT+rbg53Iu2gfr
flh22VZwjCb/n2Kn7Af2I68cRpJdFU3dlQcDOP+Ljll31w1VHlAwfOfWmEy1PYB1YRnkBFGC3jEO
x2hE+uI4l4JFomYsqWqmXh/wxJXafkPgyrRLULsxN8On2a5elp4yzoLmt/NdTpwTAIYpM0DGXnnF
FS2irnIFftR6XgXNcKKVpKJduWn91frWRA2xx6Bk6mqbtHk3krQsw3F4G3PFvp3Oc236EFRKVg52
XeVGIH1zNhj+DvyA3yggaVDUmd0PFNsV9CObez15rcmgjAMDH3/RoXbOkC0D6F6Q6QgBqeDP8lmL
wzNru9pCKcDnrzFkjzsUlMd7FudW4LLJf7J7/MFKjn8k1PrAc9RuH3T9GEy16YPeWauNqW62K3d9
ZA8v/Dgq/UDakg0YB3NGaTRIc5bxyJuNPtNVxwR4q+Gja5vcmbEGqqKRqU9pKvj1qPT/AU1cvy1x
BOPR1k7BltDNr3AvXszDCGDWD47N0fvpJF/DDO1fQWY4ppoVMGsMhG5xLRS0I5Fnc2mSrVfTlote
qSRdOT+5v0sk/YKQHd9yEAbEqSDL1MJkKDt608Tbl/cgcelxo+ThD/fQ8YkG7BUG5YpLwmrKyN1A
DFSM8AcPW+tl/wCiiKo3apOx/XNZ5kf00u6p1u5Y29I16A5S5IIfB7rE1KyC+PncqV7Ju4tpwfF7
y1hDqekfTI9q9BBGQLcXHBTBj6W3ZEE4mTzAEvd4fb1cdLFU4morIInSYNClrdEaPy6R91PFQ0HS
AFYv82gQlwltn0ZuxkUJBng88AsNA8OPnTpeae2vtfCkdLMeiOWgJ5mRkGMB/ck+W7KyWT89vs9z
+gKmxQvDyCbO7IFjoGfh28ENKfdTB3y/j9X2g+2B4qmS/Y3hWOtHvcmx2mz1laAYZHcoVYJAbXvS
F9dL3OvyRis5MlCe+2wDuMtCs3wro97rCsKEYKa7y8jQG3zOpZVnaET0hdpoNHKjwzBykijp5zj0
TmqsS4VF/fZurZiRzRZcxnNRko+Rli6ROXnNHxQzXQDIkLwVu54uzuGq2Tz7Rue+wDvg2QFxKyhf
FJfqi5/3f2caZMvs683ahJzlhUQQgP3H2LBNAqgOT/nBm+44jJqWDf/ybL2oBp9IPfJCEcd84tmi
B/YlH7igWLHzA3VYWibWTvgL18cXkBpNtwciDvAf1CoKgLh1Gi3qvVwyWfAvLJfAxfmSGtKuVKU1
I+dcJ2cz/WYh5NAHxzrBJgWG4ioqAB5EFlVg+HPBGnfj2Mf/E/OCf3M3kVYT7kVPRDbTWe0wnFr2
qsZI/iCczlMNwMrubJwrcw3QP3+fcqyZCFrc+FzX/uNv/5JSA9UvbszNXoz2idR2HG1Kb7t1kW3g
w2da2TbkXh/IFJk0H4HMslkKWFshO5rgCflNExiZqFyMD4efHAooNeCu/AGpao1jcl90PAVbt0yT
w1ifqudSdbBzmc4vD7by8zGJjrKHMgwy7NgwkArbphJy6vXmtdc7sNXOl85smijSophP2pg7h33Q
JgKBOhjD5u0GlZxZS2ui8MahTdK+zrhg3M96VsVU/hODMsRxxamwngdA7oCUrnB1U3fvpEsSiHEC
ngCS3ubHvaD8vAHPLpqa0cyrW07BLfyVY/mNBDl4BcHeyFMTLnmewrmQcLCHkqYQS74rginPfbYq
ecisBlvStDIGNI34/rEI1a7nLtPgWgIdkpCaBiGGuCqofVDjG6/gZBWPAg/KYrYvLUE4ahjlRiLR
LDwACnf95xsByGfBzYk/yZ509vioTnlYguiDZqnRip1DMIcAV27kK5rkuMwlzwgyqIG3OXh3iHJ3
f3GTRZEBf0WFHVenUPyGksG2HyIn9VRF1ywa2SrYUFFleUNmApmuc8hg2o+GwuF2RLLuU2/mrsah
f6E3VLItB+MlzKqCLGUdy/ak2/LTYb2tEKepyNi+STxD0BXZHJRxT3X5ybF90s30hN5aOhC1ggaU
6YiPK4naULiHqgvYcbEvJau1MJqE1C3qrq0i0fEoGHFkawz5HVMwEYmGfsfy0IGuzUIqJ74gKg1H
/Rop5uTl51GiJM5YKVntoj/5pBCyS8RWRyfJmxGG88LJWHcScOctahrgX8OX8vnA61zrled+dSRm
HCy89Re/Ze2n4ZSAV8UgqFUxTg0fFVMVR/PoQpzsRqHnwK/8juW2MHZwIUL1Q+zMXtYXG+DDuQ9+
fNq/mkW2L65cUcdNt2vIejnNFBT/LrO5oRjKdmELGybFK/w24HKSWqDEVtFrXt9uOj9jWAKq7fjh
x21pohHxCDSQlUGOSQKuG5koWLmmTvJ2i8oUSi2zaOAbLzIkgDxLGAu9GjuQ0DRvh/uX1PFboOx5
HLUQ4t5L2B9g6CMT+O/bm1YkmV0BN0nAc8UdeZguZOjDqkiYc0Fn7fAoXxz++qaThmKRlwoITE7F
jWRyL29oUFCecd2E6yNAtYJzwqZUGM+gde8D6RdQJYYLQ0wQHdKTB3y8OwPtDT9Fp6Csu4kZAJCo
FDoz+buIeAt2l99WaGs2I/DVbDpv8Q0m3UyklJKN2DH9b2PI4xe43Hf10AGXIAgnq3/Uyg9tDIz7
XYCUXru5QtVknP1pbJMA1QmKbjA46umjFwRkLNsdfqCdnS9zpPiigpRU9+l1PV3uuVu9QgYni8J0
N+YMbaeADYVwoNROFtGCw5+ljJJyUQQvoW0+XR3BFY8kiYZkpCjHe3WC3hWrTz1q4phtaRtKL1si
2YGSngEEjicJWE+I2f8LMSYKqqp+uZ7U9FQAxx8NE9takeK8HtuF3LdobXQfmBEYBBdTCZPCxiSh
lU/N1fj1lkNnQrgYmiHIT+LFlvgcm/5hNeF0nDNZ2rxqoNr+v6Bt68fFcKQREWsm5fzLD3dMOR08
Z/vPk/rj11rZJXTYC5R9ca4W06u9katHpF1j7//UvzLMlO1xL9ra05Yhr1GnS1Qm/Pg3VENM0tEc
WyGMBIwziT8GaIzwSK+HVO0TfLadXyrjpW5PiCROLXhWWuzvn+dSVsxinnDHRLGkTe3etYWkVdLk
5wYtyW4TdLa1BmQZNUQ4Sh0lqTuN4jELA/4Y8PPw0ZMQJZCQBFWLqDhzfVCbfFIcbMUjG6hWsLRK
Z8lCcj+3atsWLfOFH1yC0ohVaCd2YcVprVN1LG/As/ghqarS0vomL+tlPQbYr2BlHyNLumSJOzyC
6UtdqSyk2h//f0R/p9wR+sFhNAMDlb21Ns8gWnw8YCTo7iI3sUys3n9CdZn1/qJdoO3r0sRMnJF/
Zc7F8TQxJPave9+9uPX6XNGtAWuMlytSTcn+LFN59m9nzQQ/HRcLZcTHVKlpxYBKOgSE2nYwJVJ6
MLt9pRwhnMVITaR8T5+EX6I7BmrL56lmUbT0loT1Do2rVCMjhfBr7Ww9jGLAvKmpwJDbYu2FIjIy
RI54t/N9q3VyZvZi/Vr3wJtkf1hq01/ZKEKiY74x0V0K/FvHI3BwF1WfZO2DlaJcMwuOCUoZGdjh
59UqMlm/IhVbRbfqzfpwOkEYx2noe4URs00jcahXa7dWUprjR6BX4UBhUtEPObvgRPXGu385AM6I
j8oSZ723FKADSPRaTtdgry4c9OIAuW2ZVC95xxFE6c15rVlFxNdqmVoiRZXKEqt7k5uvJt9m4pQ8
AfCDHoGmpTFfoIQfz/cAOs1ZLzG2VQTzm8JnKTyImSszoge3LX57x2wpmNwNI6THJvRP1NYAkRWB
qsAV3DbxyRnMJ2eGQVY+/30lzan2rp1WUE49LSHU+IU6FzhqeyOps35vVJIw/cZfK14sHt0G2ayB
HxjWYx0g8BiGpuBq62c3I4kqMM+aclwUgtGWDw4k8MCwoH1tsOofBL5rNr2TnDKwhtSkPFdiXx9N
2S2EcbJE/El6XPpt2gmYiwIAs1xQ+hDlvTtO92GSqKaI23HHHfrvNYYIY/sJvgJICxvQa/f9UWTX
jg1WyQtE5eDCPZVR0H0jTIlcSPAjWVN4h9Y/UCV//awvlTex9xdNSAqfFmMpIn0NN0EuSIcPnKQE
6Mbtr+tOBqobVbSjQVphegty+etiWU/A77DiGD6JlzKCuVkWFJzRmkUv7Hlf1ESCZ6l3hBMtPj+N
syTeUlUSEioJnK4tCc2idBb78agG1UqsVGv4aWHk4zaslngGLwQnjnUDoDj9bJH9Q1FRGh1stBdJ
/tX+5JJzkSRvGHbGqtpjpVNIVpshSjTEnUC7CbEwxPI95DwvdHqc5GaH0IxVN3pJUneSE0fxe/bQ
kam0/Sv1BQe/RQ1liYcgMZfyoTLyNTRvEEXE58OUKjkJ4tgnXYyNH2NW/tyFzSRaYP9+MVM1iJnv
E/54L2iYGhVU3EwJQSN8a01+39LDtn2pKNx7XG9bTuIiNwAYuU5XBBkhrbVSY16UQAK+5DJjF9as
8w6kkIa97RKWAeeJGDd46KLbhOFYm7hFhZct7YlCksk/mpvInyPNEqSdBZnvjC9P/daFv5FxtAIZ
pOBplO+pp1jnFIfxmdsE5VvCkXRSYdgX5OwtkDTeU+qdOlA0T1Y4Q2DuNtt1HAC1QpuDGsBdZ1Px
REd44Y8N9iVwuXiHsYnTUkMFujKUbXylQmkL9CnLhfZs376+jBV43rzv478ehkPIma2BoFYaRl5+
gVLSzgFOeQBCw5pk8aYQlEhe18DeuxC6UsF5rMjxhOA34SYX49DSSmucik7FCXOY3HuI8qlitpOq
t6suxvtynxdHcz/en+Vq+G4KIYo6ggqPGlOBCmN1utiUf99pOI9PltRlkqLlkWV3eoIPgxRow53g
zLgdvfJVMsJyfwQmGLOcSXKH3sztaeTP+boBQL+0SGZCWR6Hj8CSFExSm5c6EpJYUV1Fg5a/PnFW
kIrJZWIx5G0rsTi8EK3hPWdSKn0LtKA2cTbPh9H3593dVjQzEteGzoySsHNHNSyH6PIC35+r8Y+Y
AopKv9061y42LXXhE4wCtvHQQcB5KluuSiLHzK8AJFncmzRSkGnTeSj3Vcu9AeNnF7skliS6lQEz
RlVfOuMENvvTntXsoMDsmIF5RlxrBbdgoRWcyTqHIu6qkGLEKAl3mV7AAKnpYpY12fdGDpDUPpCh
7M6wxf3SvbLkU87wan1Vnu+0ugF5PveBuBaNpKyYQdLgi+GannpMB5WlONMh59EnNR4k3XJr1dDj
cCv/p3Es/XpMNguBnodimLM3YKAU92ap9MxHEuWQqiIwA3cjo1QEWUEzsteajLo/km2mqtxyhRyt
PxX2KzOJwODWCIMCGjejsBLMbxAZjiONRoqPsPi0pD7aCa9tlRRxlTuPzh6Ou1EWbOhxN2DfRXkU
jYX/1dqs3dS6l/cBCe87Hft4dXh3LCkrIhK/Ytw8ZM5tLLX5X4mEM73q9zlhPaVBAU5GphiboJh3
yGxI1Em4dB6wUfZ7NEkvZw6xjV+VVNucfGu14Sz1e9BxMB4TNB8zsLoY3OdZtqY6FCgvQ4Qj2ar9
xVkpzBvY/Ikt5gOcMhlibFRvvIiMAgAjm0Ev7hJ4k65SS5zNsVAuVNMy+H7RfiF/fpb3Mi/Jwu3b
JETyC4CsYL/ER1efHP9Ku5fwXEgRAQWtGHqmpsJfbQ5nbGBkT9ryPsaqKGfaKTtu62HFNIcvGvGM
ncgqHjNO3B0xGDWHMtJb3BfcJydpL3VXCjmJLlMrhUBNM3hsdmyt8CHHsIzHfdiURLVm73MqtLtG
DTVtp+qKrsaEtOQxz8UgL0AVFQ9KwxejC8ZczixcJ8rE6ODcikw79Y8/twBJhSNAUykGCAA8pDLl
EuLKqgFir2cGX/B1DtWQG3stHbTHoBaZpejjNm/lV035TXzyzapD8h7z0Y0pECy61y/TACGooz8v
3/efGh3m/eX2LVOUzm7Qxw5z+s+wywE1Ghrv5M2KnonsyfaPnAYEw8Gwd4LUXbgSEoFEfGROZJWL
tNvs7YJEOUE/a51CRty4EXGxkBDGFE3ULsgwiA81rQjUdMZpi4a57VrHUaESrkOGbtmysULTM78c
M2iWvE23Ez8aY08M5zOqZ7PF2KyFpJe8XXCPxC1P5/Xy31v4EKjIgE2San5WVu2IQXI7UG72fTel
2ilT5llDnhZmNua2Aw9OGcv3sS+Dd7VozTPUu3OsUKdisnX91hapzlNXW2TauawWsnLFapdC0vfn
aj+BJChFGee5+/DK9gkSGjtMTFwCu4a5SKujtYTW1+FjyJk7hMHhi0iDcuq2TWZcGhiZHJCl6y2M
kbXe9HTpNoLYVM6zG1r0fBnvIG5REl4epxgQbEM429URY/iJXlC+sR9z/2DA6qKxiMi01RXDOlS0
q+M4FREKFx9GIG+YkFCQtwfgKXXHu5W3ueraS18L9q90/EQtlrSSvRWOSc/kjI1QMrEUFRuzaQ5t
a38O+yamW45clyEr49zSkKgb3ThcQjjOLg1oDXiTvUIp8Umrjky8wKk9AlvbzcsdEPpGdgLFNlFB
R4U5Ysvfa004S3ei5JiYpGheio2txYshUVVshHXLPv/8BukH34Pr20zIw/zQPY7y5XT+/WePusRv
drgXZjjmsL7Fyql2WuKND84zabMM5R4bQueRd1WiDiC+MWndfIThDSTjElrulr9boUWsnS/a8w+J
39/kDdDjSWHzeKJ1vdEg2fdAGTTjDCU6vFvNmW57+Ky4oFrIwU6Uv8yaXK1X0L0BvGHseaLSPgkj
I5XJ1wwbM6AaUfWiXz0hhCUrCwNAPZGca02VK7/gsHcR836d97JQY182aO2J+IMbyc4GSnwXfuo0
yJB+XyyFLKAm3XxxmknrhgNzzF4DKEe8paqUvumzouczbvetVvhkh93a31+PW7J9Iqbx92gcLfu0
x0X9ya6isqSwX65RlpMihGo5P9Uqv/qhMuP6JAw8QD2roj/oWf9yCjqT/zbNriwnMyI+pPeQRKp7
7v/OmGwVLBUzvHlhxFDG0ggrUELVO9Isk4HgPVdlE/LRXe+g4aVbsb6kfL/wlJErDZwSPIjdB/Rz
QcLTzUlnQkkzqJR2kcZ9bFl9GGOEEy6+dXpDqJd58J5/4+/8s9c6nNmeFjIwr30XUxRBnmgkl14f
JqbXC1nHDAigTw2aevoCQp2yVR/xeCJ26UGBE7qcWoku71bLdXxPTHI3XpZZKMRuLHj7ZvvSEipn
OKQr5Y3kgjAW7SzrYErvaLUb+JFO8eO767k6KSlP8yvw1TofCMNHptnjivozttuBT9zOY533Wyri
eJHeJvmB8oa4RGIyF+/ObN1OIBDvmR8uIO+r7cLoAPnfOcDtGgY2AjvxuCJNLQc2wHAioQih9sid
rmvVJzQRaF5WxY//WQw9dq1oMpgDsYnC5odR3BaeSbFO+/zanYom73LWiJElAdFFzdHxF15wPr3b
MaVuuey8GOmYHrFuNn8MX1IsooWEvnvZCFstfJ2d8FtohyIIimgUCk0tHUAUX6SKxdm+VOSnc9MZ
4JBRat4UxYSq/poIbJkD1BRH87s7RgdUcqEYLxqISNa6MgPkkLiqq8mLKl4X5+bbQcnKcARxmucJ
qqziUdXiQl2y0qUR1NgCT4Y7tZSd7M9XrBdJjLEVi9ARQxD0MbJALVNezzHN2zpcK337UzUw4msa
hHk9ZbMWzEQLG2Bhp3d7FGXjZiiKH70m5g2uckpVsegeyro2RBakWXWWoEw2LUGDa21gMEND10mf
xNqX1u16bvWHS67WoslThixr8c6aRApbHO3SswoGpAR4APb8gEUXRvKoEp0JNsbUfJ6BXg6mQF/J
/WY7Yax9vEyKdCXDKIdjfpT/RcAbt9mDBrLJJmgBcg7ys92P4iq2/whh9gdmC7lSUl2yqZ9sY6QV
aozPxWGSeVETf/FzezD/NuGsKAKUdwfAZhFoCkbczK9HhlNDrA5vonaUSNDPJn5VEEjn3cVqezN1
gpkmJh6dRfU5X2uGRcJpZBcMfj0bt+waP7tXa2CrvjCk7HpNKLVRjcVYEeFvrseyk1JPOpiSeJOo
x0ml4Es6wmpYjK+H54fempeictciAnE+RYsNrWRmCIUWFkLkfEeOMirB6I13LAO53hZl48GPhix3
3rMWzVUAMPMA6YiCJvZxMDrbxAR/KGIYzQvkRb/oUK+sCrfl2Vnr3CyTBBmDyMN6v+vBKqPHKkhW
rEfCGRmvaoFcWWYD7yipZTVOOFDfuVO/JpEEembz2k8i4QPE5wNCPckqP1HtRKJwnPWq0z18MlXo
Mko3EhfCPgeie8WZeU7zLnV5ExawBfSttmOZ5TEn7Ay7UjFlagBRNn1xbX1Vt5kW6/478j2xRrnJ
uAAyAdedcErrnXJ4MWdkh9qVtyh3NguM9KGrFzKutaxhK7XkJw2Xt+AK1nuTYE+NFhvd5PjRdCRy
ieyqHYg0xHZVRjOejFzESSmlPJuyt/+c5d5s3Ba4CpZS75AkkB27Vi/vW5g5aU74NdOgLc4UsvCl
r0s2RmKiuL6mC5b9qUhiM1GzFN2/umdvCi77bm4HMedwQb8u+WK4uUWKlrZr4BH9dEykDdadmTs9
zsNmT2USmeACLrkaBb4rdEJzB0wwDBG5xmBFezQmxmukQDBnoLU02/MSAz4M3hb5x3EGMPHUBbWI
iLmAyddLZ2xZIS/BNHtmYJ9XBRrRj5hWNC9YKb83qiyDKZTeO93f5eFkJZxkZTW5dLCpG68HTIQu
j4yoIa/YOhOCzwMU/tW3oav4r7pZyKMK29E7dTK8kUetl6CPb7XQlbOGUwU9S9sy9V//Eafz4K9M
3A5D/wrIUKK2ukNQmLOzfbD9I4WiJdjqn+984UZBz3ArJKwP1dGBIs8zTPB/mDmiSniyuNZuwD1N
Ka5fuKKbuP7OIGn4LwI1ryMSQ+RdAhbL9xShH8k5OOBiWm7BbRPm7Yz+guEmoTH5qtBfXOqTthlS
70HkLU59Nrzu0mjtnU8DJ4KW1Vxrzc2l+re1MB30bqJc8xrMujRUEVZ4Vtvf5nNrI38PlAqQCLa3
irpiOBqJ+W34veh1PrjzIjO+VdDVBNTgyR3UknniJ5AruHjRAet+QKf4H696kXS2t9LyeAYBb0bv
jIatl1sN6hOOYx5YlI6OAK2i/55bj0nNDvS59PL5XEc5Y03L9PJhk4HS6OGuwkJAbJ0FkRRRRRR7
hIZkeGh7/5cTNyoBMCzsm3n5qmCNaFeBimi9E1CmkcQLSr0vAxijZL7YRxQyszTyTLHyF0dr8uXU
SOjo367mxWA1meRbfB5hi/vRcX06P29+b4oOZg2YNqi0LDzN04hIznn05hmZmi+sQYDrtw0Rkc53
o4pTH1ejExb5YFetAbpo6PYDWdeYRlGPsoNE0IKUylldKdPtkN22eYk71hQ6EIBGsqda0iiOqZPz
HqVL0xQcTu8HGvlyDImbFg5NgczZTbDxbA6Ri/ZY1RYqI6EJ8+H+TMhUBleN2V3jmWnVDkpgu7yE
PKu39SLXyWiPkQ7TYMbvpAmvowCuSKKPwGzCwfyfz5XRfIUTYq15JZaZEzjuthFH5rV/SjquQA+R
pHutrLMmJhM5F1QyMGe0t3eXCXEWBP9wPoUa3pZJu6YQPo3YvQm56V/D2qcmaE+jywLycb71exoy
Kaav1AFuwUvg8Q2AwcAN1X9BxJRxd1KJidWqKhwVKlXZ8CJIk5Jy7oVhJDquEsvDy/FhFADoqDHv
Z5yqnG0qP8559GUiEBi2wbsSw7dJWV8sR+U2pV29QMW9U6BTUcQOAa402PBu0Z/gVcMkxrHD2jlb
JFrmoy2FBaj+3jtgwNOnDPSlWH3+EfSA/pS12e8lD3/78Ntps9XtaCbIaqTLamv0dmYS7YAQgVv0
iSQjboWlpmywZEr8V2dkne3RDuoxA/3+F3VdAkgpXFgvYnzT4uYTHQCUChJZtZa7vT7H7mClaZF4
Il4VFi5FSifcqhfZBupZPqV1H2S0PfdGMgc59iOrLsv4t9bu/SmLzJVJrkCVUxF6+nnhHa/GEXtl
/KPwS/NgcAV0M3qjKoizjK5zAnkDNg758RRbqHQNM8Mpf24pZN4zgYVdBlVVNU9bsA44QEF5O7C1
coHO4Bch7jeQQ55dxVs2cBASlbpMYkMOqO0lm0juIx8egp7vQbaofX9gngSw9Vk5j8Z/wX1Fyx5D
77wDkaAYv8zilAh6aosaWvgW7TH6At2xD1rsce+MKHnFtQthx5xD0907u12fI7M/ptxKpCIut9Im
yhTU2lwHAmOC/LgHnqEmmwdGWr1WQMkdrCEV/buvw2Eyd+1vnLdrNfDtcJytsQ6Rp/FeSFkbr6+l
K3ElKulxf+LVgGrYsSO5ulYlaegEaWw1N0u7MHhUfHfM2Vy7SdjK8cvKXOIaeAyC97BLw8hUCuS7
gzWEdJnVWHGhh5vie2OqlBQQKN+99OHngeof8MJtmwgjIUGOPqJwvgoSt9/3166QhplaUYiwVXER
uyfEeazY8DGB4FyjbbwK+sePI6J2skZl8Atqx7MqyNrCN2gz4HQFQkDg9EuPXGuLoMwBLtRtOTPA
8ZhC08/iEBi2/y4fpI9L2IK+IoFT1Xljr2VGMdomKh755gZ/4iS0mhXOMVivWlPUaXUMAgHCDFpG
gdqLG5n4Ibjqa7POPdhG3YDr91fhlnnodnccbkGhhx7X3J1ahMEzN9j+fzJMcdk9t7fULNSQfrsJ
DKBHkkYw5PDKcWfqnC8bGRJ1kaSFBaZdD65n6NadcsnIxvVDvLP/OkJzkV+p/8SiLiruDsHUoUqd
MXz99B9eScn02DXCjpQDR+s5tI8w+aTLteVXfndPw25FPRqbEds9EUlajlHK+/vzWG8Fchpjq2yx
mo3YymP/5AexfZuf7bMq0CP/pUVLXyBT1ZFTYVwWGcS9UURWdkM1yjvx9usRPyECkEI7rb7z6Eb7
ZeCY1krP0GNhvTo0wl1dneuPNFT4x/ojBUyczCEmr+fzUHAo9v5kgXhble8E/NkqRareYZDil8UJ
xz3bQ9EyomitQAV24fqxIfocEbt0sFuvsOQdD1tjsjVkfmgy5WUEM4tIr765msOuG1dklOAscy5F
6gYKguPpjHDBiEDstu/habg1tvUMReeXiqF90BK6iC74ipWxX6JiUli/vgatR30n0oPP9p6d0SBV
+wlSOU54kHEBXM32K6DH6xuE7jLtdSujc7kZMF30LqDnCjzDOqtUb2HYvLsGb0bmiwWaSNiq0+Mr
iTqI4Ej2rFaRxe9jTOmcAPlCTrQj5RxjP6s53qmqLRzsr4MvUL/wRhJLZdPRKR4wu9niOPvHv9CQ
zq45ZBB/36qyOm/qYGx02+YeootCNAHGcrvlS86L2LVC3cXroCX42AN960R3ENmJyFL7EHw7McYI
CAWnJiA32ex85V28qtbMOkTsX/F2HwCLqGELGz3oQAT+SZ+USy4mraUgu2l0OOjBCf42kOBVQMD7
SYPVHwPTifRY4AxvbyekmleP4AMW+as+tkC8K/G9SNHLl1OTFxdZRo0jh179IdKOIobhACz6Oyh4
poFC7MHdY1LVxYw/rFL9Ko6grsmpmATcieUA87YQwLTycGwbRvHgDX3+6bFppRFh6TORvpsi+PzA
Ys/srsZ0WDoY2GOuqdQHEp0cL32NB1oon0YHW27YAqtZm3BFgTkuZSGhbBIZa8gVP0xcqOr1JDOI
+fnNaGmpxZziaUXflxScrf7P7AmXGIZ81L3Qmz5ZvufsRelNZm4YDbNtvMD9v2v0e5Fc5I7UuRRC
OfgVXwKEDX+zLQIQgdb0OsN8P/lMr/l43yG09unceAK9BJvQiSWkOqG3VJx2EkQOW5i+weHbwTBx
k6xWpqOFab8EwKviQs77jxvE/PLDs+OPEJwuAnnsfWjymc68H6OBi/DkDkuO2pSiD39hA8dxxsQo
0fP9Zye8NXAuIESHouKhEiRsay6a2NWBBonVkpeAOqLR3FXWS4dwL5fTL04B9OxcnYJihXmCYKYU
DwavHZMNAIDntNCcnYy4lncao4VklsxDq1bwXNRfJ6gQZXZu/N9w9lIHkaX4y1trSq+5g0TKA2yx
gLrJWWENebi/phW4F/uzeKjNC/QLK98Wf1IS5mh/hy2LzIfPSN6oqItWEEUdNPip4PCeDbQnp/5I
kOgV9CZjBnULnGUNrHV7RZb1njMq0AynhntthaCW251tzmec85kgOmH5zughrMeWX3TPVixt3jQw
pJa1r3s4FFOlF26JsCXabykC+q8U4wtHPNLumJNzfxCv9fo34xEw0UrFLCICHCvdyf7wPWiRdNHr
oXB/ILQE1N+qGO3VeuyMVDce71nzfyUGNbq4zsZQH1kPq2g3T4qeT4tgU05WD5VWOCC3iPMEp2G/
obYPEV/F0ugDxSZQy+A3qa6AhlngEUBovir0lYfXMFldSZO+P3/XGeuZEqNCSnsHRLjCAep6+rCh
V73mJUhx8WqSPgx+1ApTj0hzZTN9T54olb/SfrZyDNEqDz5TPxKF1NF9RS7/otozlMv7mfsADxPe
yPr4t4eIjWslFkQG3lODrdFCjIMJkmtlLr/bquLHsL50indbpZjdZS0BDcIz/X1cSqg1FvHX5qv1
6ksJhrzLzCNfMGotYLHgnmdWGjJkIIzWfviicVtP1EGGRxN+TAb0RsuoVolCyFOf0JSadMoYjcs2
T3qgbC8kiWqPJL89g48rHMVndDuCtGtoLONUv4lUdzkKKkEvEhwCbB1Iqjs0oKD0ofZ9uuovAS69
1XdOX53hDXzTZGufRfbzc0GjU6bUHNELi/iIp8FcIqQ3y4yrAUmG0qqRRq5bSHoqkpTB2sxZX7fT
3TePBgAMXmFesTc7Qs0nKlBGWhiZQ6oYWR+V6zzPE46za4op18YuUKlW0/cjeJ/RqgMEU07W8H57
99pOKXGE9AYd8ItWbL2yRrKLSDCzkgibLllxGuQ4ppIlbAxep9JDBqEHx1OmzOyFtd8vbYIcueOT
bDeeZeEoyJChLY98P3GA2+X331xigJ9VP6d8iVbRE2VjyU19AI3eqVFbhuw2qrSf3P1/gT1zBmpm
AKppq5FHdU1dOGNQQcyqnZdt1/qenu/W0jZzF0LTJcpi0CkmJteHMCpJDpk4PDip2MSHA2UUeKCc
PaXhq1D1b8VL98Akf6IRp8+GSSPo3CvcSoMf+uPVsiR45WTZ/eJiFvcIrKGvTllu9/42CxTRSWhc
htamh5A+wf68LGv7wbI0d96eTNILR9+H0dprP9IU0E1qtcOlpeHgB//z9xGStPtX1v7LUtQaYAlI
HnKz69iN2tU1P6u0ABu1QhO+tfFoGBTO52xjuxAX7LjOgMeyYYDUn5TO0qJ8GGXZ9BTYdcOjzNQO
vskv5OCr7jGuzCkpkCXwHQ8PAkqcu5YnSqMxQ/rvDyDjqE800E4UGwe1J1gzfeozvaQtX9Vfw8ja
psSDuTRvqEnppdFa/8aCy7oTZC5Og6xmwOBSsi10IZH2qLfBm5sG1hi+iSvXXfmb1lJVi+5PELn9
NEkULIWztf/G0xBwFZk6YWoVqVmsFEsJZMb6cubRVIgJ+KtQsVl2r7cz1TSrq4Z7fZY6EZNV/Z7a
NMH1UHZ5YRYMuohx5lMRwjUnIpJJiC3DOlOeulklnmyTGzj4VlpHU4YFc3gKPxs7YbfSAsDGFEW2
4aAMNAIwq9PFfii8Meyfs1G3OtvjrqUiSaA65lM5vYMMgtPhtzYSqTHTKOLP1/59X+9YBe9VLhyv
JSjj3Nq2DjAAE6829QMpWy/mlRc4wngJ48tdlFxE0l8vU1LGHx+oH9vIfmDnU02XkLSf67JJY8dF
qKIzZmZznRjGaGqWe7Fc56kybQl7J214Sue6+47tW9vvmqkEzmCBkbXo4fJ925rl+UdTFXdQ9Ojk
Z1ed4TNnpk79B1dhcj1Wbkk1WwzvYFHTBllc3+crJdcfR7GMFXP01S3rsRKQS8q5J1d1DHelMbwn
flXx+1djwVMhoFBPVCnpTx3iiOx4VyBklID408+h4rwcEHm85WX3SNU7N6QMHCUu5vuzgfT+uJiE
Jyvt4s/z94z4x+jvAbUhAc6mNDLiGD+Aibjzi1ExRmWCdWyu/4R1dmU/erKwVG3S36cLqyP/fvGX
DzCrLvc9o1aHCn3RKvCu58tcvCwnuu5Q8UYUK7SzG6RpQKyx2rI+dt5HUiQYf/UX0RF8zFqoxaNy
uvRliLha5JdedEJ8RD+UI/CUIOFF+iyJ2nPd4eFA2AdKEyT5FiijOyUdCQ+VT+KdhQEfbEXVwryk
iXEsTV5F7oBh7O+J6NNKgbaABVv/D+urU52KZlZu5i7qFYPif6AZtmaQSdI6T2VHdoDLzZ2q0dC+
8sZacTWP/hcPM3nG0Lm2YNd4H59pqcc0f0GeHVeYTE5jz6V472YYyggkFK/Lx7LV5NywYuzcZ4ZH
ulkRwyaW0xIX+LFoSxFT4lM1o/aPSTT7DX0kXtTfUb32g46HB3nvYMKy4iBoHdGAtGD4VDP3kR0k
TH60tgbhaQQirUO9k9RNNYhsoLbSdfvcqMDlguPyLTHLM1AAlM5LsYRYX5WEMBDLa70t2hoUvGMH
d9Dqk4gRi/4TzdLMpwPYTvxQozNbzi7iqXTuCrh4m8Q/SlR7DuA2e4dnr3DgLXdWN5M89TmnS3BQ
XlgRxekZH9iUioxCXqcJ8CwH4pcexJcVdSRKwT6Zk37LlyPp7xzqR02gK35uXHz27OtS+kZQnKKl
VuJomwbBpf8RPDznMeSk8waR4qc1E8zImVyr9dEM4143TUwPMwsiZfn0xpuJi3mbuxfa2wOGbAks
qLwK4Soab11mn+3CxHKxEncfuNW0qqcffwQMeNRJOn5IMv2z8AtGi9TumHZMzVXfJyF44Xl7G3oK
7o6qkhftW+h4ehcZFD+SGcjiKSbCq57SU3NleKPHwYMSA5tZu5RZw+Z3uvf14vZNv9xzoRIGsM5A
5JIXQvgQpJAT3jRwjn8XMFNn8Rpq8KF4UoRqazqyZiwKTrRuSSPmZCDqm+ub2/M4rIwOLiT/fpZj
jUqsb6m+2ipWaX28AerBW1PmXi+bkLQlhsjUF2m+ChQJQREbOM1LfD+9TUCaq6cpMHKwi19ASULu
72TW7zClFjqHkim/w/d1FDe3QZMHwSIefcPct6Tq2OlQ90zdQVwXh7jqfy6tqzei3Jcf6h+BttNE
zRcNaWhFoOaJg9EekqhviY5CGLd89lrkbCv5wXanyoUg84bgS84BFsmJcKbZ8V4+BrJNCfatAaIy
2wP4647gvQNzFQ4fMyOsY8rjDG8GGM9PL143d6BOKOTgAM9xHnJ1oUgJbeA0slRnNnwbE0Pejhid
3qV0aK5iLerXZCKKlrtr00IcXjyMFAuuALfbNaDf+eMXUOUb8tfa8Xud672rYH/yS5Y0PaC7aQWG
x954g8qPOxLTqYbjA786m2ZpxLK3zll5Clcw4oqcpTuGC/E1g3SvKKl405vfWanO7cDGuV8R7Wfe
jGfM+QKAiPLHznN5pqnHuVFyxRbWsjDFW86EHEyP36morPRMmkUQOe4l6C+eKThLGuJnQJ5UfNGT
iGrOgJNJ/XVzQ0mIUzFZ4o2Y0LWONULZobLeOMgqbXVphUvFy3jjbJlirjSfFkdnFpgHX67As3v5
knjSrth3eb49bh0HFYFlckbAv80zklF2k8f8HaFyfnfgXcgwA0MacnuJSoI05DbNUtewxZd3bwJi
P6sg5fZpe1lObEf2dKXblLJsD4r5qXiV3B+SpT6F3OTKKO/MbwzuaCI7ds1kpcHHoWPJQycv5VEm
nLHIKHpjQKXYYNjBMeVJyrYE2DdKS8XjcoVs/JeeysxJivjL9w9QvU3fuWSFaPUW7WUZbTqYa2uh
Mhai0lFyUg3AYh8XI0Efs1XqBYyQtxkJ4CExqIWEg86my6oCIaqGw2R+5dkHqAEPpxdUqgYXb6N1
UAnho00+dXAVXiE0JrpmRIHNzDAn3Vy8LEnHJL8TkLKufbcO5mjXgpmBawmZ56vpHGoI9JMXUxuq
cU86K43RufRrIniXM1J39N53c9am4Ym1/NmYxk2FoYA5L42SiOlDoWFXKVCA0vVkKwgXCCoLpscv
TAXOIX3jpVpxwRbBL+zZzwJ+aefHeY1wvZyJgcAVHcepp+e+dGPcFkpQDp+REy3IprWt1wEGV4sB
t77t1vAeKOJr0/mesLTAKCjAxFOB9MMbtLtjYFR3L+I4pd77AMMoAnbE9jjlTV9JAi2c485h9dXv
9lmUYGlqtdL5m7b300X95iihyNuRSe50mYMH/knTNlTAlvErU7Ln6zuCqo2aKCh6a+wG3zw16+0s
lZNyEv3b+QzdeE8QRoo4LjB7cgxhcNS686KMb2aWYH0YCtltgwttI1AHDTxRaVblscfmNAx7WCGt
orz0b41DxGcTtqUmf8u6horNuQ1M0fDWh7Ynz8If+3Sz+FmoW6LFc6agzHZ/sEmJ72CmWYbXyRya
+tIbH0JDwHIKlgCwljmoPM8Be5Xv+lywslYLRmNiJkAXr93Vat1h4XIlXoyS6X7NtCQxW69u7k2D
dUv0FlpP7H6BjbFzm3ZRGjlm/2V9ZUnubQKx6++Uvp4UNf9XcVylHP5Oxbm6gIRprRIUMxSMgIGq
Xua1YGEtOOCsLJMNTuWJbaclJmZwaRM41vUKNxlv+TyNfB0C01XOGJMat8mU6dwX/IaMJ1pSOkxy
9B4nFVPcjkjYDw6XQYgYKeAxePa4vgKnJZ/vb6Hw/ALsQbgI/RVS8cd+WFx0ZdV181EkqpQPkf7O
dMvlaFJ/2gwzBgtNlaze5cstzSs+3REqc/NZP7/Uu5/emwht8mZRiAl4TW/Cd9knlDQMW3Im10LT
ahQrHQFMl/+OcFUxWdqDuIRZ7P5qAThqzSOKyMDyam5DqlLxOee0/IkJiUBdHxuXd61Er7SPYJT6
vSicLXVWNGvucInbEPQbLIKe2u1cARiOSdFxbwdAts0U5eBYZvGiU6c5koXPNSb0mekNQa6akg1r
xH2OvdS8S9DBAZHXqG46/5ZQv1vy34Ib3o4YAjVnkQ5VEG7Oytkc5KS+Lyt/MS8K0DDMxGq4GqgL
1yTow39MQxQQVZcN3zaZZ18E0qetfIozvDDS+44k4WF1dRVUMeb/QGwNGEKgQ738LOWjrHKQzlfO
KJ+64yh6pg7jFZovaURPCdrvNpbadxP6CRZGwTYKhMru3TF47vn6F9YYa3nYlxTEVeWOhrGXEjBV
ft8bhVADpdYm57sS3Wna4yh9GfXe8uSJeLBwIuB+jWLt/lvEV3Yf+5pjmS1yQQFotupUOZcwYDYp
lJs+aIPNOZoF4pA8o3KolW6XYbdWDlhXaSO9T5ad4rp2si3ZrbOwgC4PqUVFcEPjaP7YBc75DXJ+
ZIsghHZaNb28fTUFWBzG/B+tXbNGyDl6R22qMkcXfRvPMn7Fvm41jnxS0+Pd19NE4aPuonM9mcrf
SzMmdJpDw2UDBsgkufhtKw1OM2BkBzg+rO/Rgz1bsf5uSvAab6EFoQxT8JHIgeURbqdtjrbDEAtj
zf8tSTylP9buD5+mn6XBkh2785VJVaU+lBu6qfuLT6B8/Sk5coIsz1FAWUEva4uKyLjVwRYaBm/g
tfF0DZxR6kHKIJCYJf0om+BpUkOMiqPmEh+a2V4loadPq0ynHTyOJnaT8OR5NMtj2amwsfh9XaXH
WYAzomNQe2jgc9a9Er6392AlCSpp4xGy69pGoixlDTiFod6w9R1doAHpOUgbh3c7OKON2PICBYU0
QeKPYjGUmiR5c+HNz9QvyuBnB6aX+MC9V0mbYSrJ16zUginnGzdCEj0YEWc7SRdosHQUkCWPc9uh
g8RD2qPIiCqGK76M1MtO8NcFfuVIr9bZyQyNtNScZk7C4zFGsFdr0w2TqGgF2MdSt1RnfBFqoHPj
kqUPhETUhzzMJTyTBK07lWWQufZpIzjcJu6BemW4mH3C8gTq8dMPfOBAXxh6V/zNvucoKNikCmFM
4/675qiGoYogcDV7X77IRDcY+VMwoEgeQ2xx2f/7S7EoCoQ7ErmKNLckenDT7rAranIg8pzdkOOm
e3p0q3chCRXeR5khr+BI045A06sFOCmCRi0Z0s+YPzfQHfPvL7TxLOGrcQjl18bnq5XcjBiZ+5f/
RrvTCY1TWm8oxzav13q8XxU2Ewx1t0q2H96cOx62viX5pOtIdRk4P/ef+AZVvydekg8rA9jCGyR4
9f3LADMp2ncKBozOahYgl0IdO66VwSPCqhtFK5pO87GXb5WEPc4oze+BXGds3xmtBCp9tmYdbuGg
Ik+JhqnvHUDz3SXlkDBZHe0Vwqf7NAx9soahqBPQLK0tJTvYCV9ggyFQlyQCCW0U3ewjBBwJRpOt
hpyw7VEF6ulKON/2pka91NzNKLUDqAGK6FYeLxBFy4y4Rlg6wXsGXROYvbvh25yKa69lmyx9ZYnh
62To6GyW4SFps0siTg9NFlK9Ap69uWWFX8ag490KTSDpn3NjbxEATNHeF51aCzPL6HepZlgph/ZQ
+/Zu7q2QdP6CM1WD8CP52PIJgzuwnXP/fhroQ+ku9tyT2NfCKaQzKuYCD2+wNXEpRPpzSRp1Hdm4
NVBUx+Nk/AEA+ooWLYCSpF33LGiPxlS+P6SFhPhJSqyvXnt1qFvDjjU4QpLQxl0eDeEmKwrpeREi
8NdCSaJ7xKQd5GI7tP4ok+K9TA3zyJjKY/dJfrFogjIFIECIOlZCU/Kdu1N3iYujhlHok7tEaTp2
olICjdUK8Rtunyz10btU77uZ6PIkXTbezTAyUmt4Ex7+PCmonG96UUNA2SN0TYI6i0IKiuzPHSms
nZRhmXindLmEcegkSfpLQZZrQ4n6P7WB63HD4WATuc3zIGD6AWrx+eKdOZ1qH6nuo6g9WQk3W7Ki
7INc51Aztj1TBf+YKbHBoUVs/14AjB9XyV1Ic/T68Q+5XdsHupo7R8O37PyWtibV3zLioguH03Wm
FU3XSx7jXKULSW5+1nEIXOb46uOPYk00XYoJynvdinAiZPpFT5HYFOXJcP0WfUfdX0z9oAx8rMYV
QCYw5fp5MCkHz19+h2pHIZ2rSvYBn1Pn7MAfUS7/nlbd+66GPlQxTZpCODZlKUKPUeDFM5LiDU1W
WFN3H3qw7i76NzM2WQO72/nkw5EDzsOwLmdivcbX+aelSJtNbtzrbk++jXprT7aLRHdObNsr0IiN
OwpKKJ0vkOj2G7ldx3GQIn66f3dc+YpeNLM5b8BY1AHE496QWLeae27qOhv2KBGvPLjh0RMC3y2E
G+VQVmXEUrxT4bCK16rqZ8iKlPl6r+vZDS9WIko0mbJTpYaTWhadJ+BFpSEYjZYm1+9Psra5qeHF
mD1SvDil2E+IxZhdej2gbGUYmRLoEqa+p5XsVT4IVCUyCHGl7SondVpntBUASE1UeavvL6dfCKpA
FE3WSx6Lsx5VHxwFs78JBpFxf/c6ZfuNXD50IWxpHBVZ9kEo0fNEgJlJtLHnJ7dvbwUFyqQbFLJx
SvP+GF2F+JYKSghVNnZHuihScHwXw+Lt5HmBwswhuODydGPyTvGOdHgYtZCoV6/QNhAGm26xd+zS
LFivw7qCI5eGCO/vhqcfqL8Mo6lZwdNOIy++D/36q+ARgSzHeMYOTDmSKLMavnVAzzJpGT1UKODw
GMPlntBSG5MKGh2z4fSeiS0V3qglOYEKwLjjr6S/tQQqFFiTRPKwn77Wd0eZH81S29SoUNE7JaZY
12PR7Kyd5g7UQDIfx6IkVvKJZUUvHBw+80q0TNIA4cQySNN+q4TioEaBy2YJ2wqDCliTru4b+tNt
M/t9knJvCeYKMPdoWbycnJkiXLlbzQ5JShaXg8LwBweIp9s8ymKXyNMvHHa4QakTGiwinT4U6udH
LNsY+Zy9GYtbJge/BZTezpdI3d6d1M63S8bVCdHtcggUW4DeWgf21x2fJwhFyJPYvyy57ApVDygm
VlIPMW3oGLqTppXl6waa3fGfa8jHMzSrtRDzNper+QBOb8n1GHN47EoTzIKhy50Wx2zvDX6dqv3U
orvCTVvtoUcZyFSEl6tKNfyzgpRc5rBStMdqcAZgPSLlMBwEiGiPqrKcHHWma3Fn0jn+rNaQ9rJe
0ZbiDksDWdKVSEgKcbZrcR65lTMP07P7Uv8ZTMpqZ5XaWeDDMiZ1HINGgKq/Ob5F44CvJjPvHZ6e
cuPMwbnrIsz0hW5jXjWcpindfWQN938AHoO0wY1fLswphZBIfMr6st/4ejQs8lQJWBx1UdbDwVF0
zwNe/eChGV0lH2iHJ5ijquk7H2MKwg22vTlEJZhVC4yWSXhIPpRHwlsJLqzl2uWAjzqbnM7t6rU7
XGjAHuSmr8CfetSxpvBv+rwNMEJ/t6Ap1Dx62KtR+vhMU3gt5ONgLGoFSuN9wm9bG7vSNAXHw2Yv
2gxiaCvwWVENqVA3+ZqrO3f4v0Jz4seTcqWUxmurRE7aoXy+ngNO0WHNvsKLL4pehRIZDoSOHcKn
kInMu+KVixF0/UNMeUEfr9M1d0aCPjfs+nUgPxzACAkDy7MXfMk+wCy7qkDxj+iKjRJk8hBYjOwR
de91MIuufSSmsv7dvkOLT4UCeNoFCgrEXSnuSnkgFS4OJWVK8p8eS+xtrO7K5dOBKE7IFLjzHVYJ
TlFyGn/eYofPWxqi7goIH6yGCnTOxpP2H1vIBNh/8aFJBaT0Fevv+QoPJVHKi9ow1TIU/POHfg7I
y3UL2Qo36uarHbjkZNgHzJvOboUU27zlp2HKGKhKIgJVzibyEDlBIBlTukjJGxkNqz8fOsceI7GS
lgawBVLbv9rezPXCPPdlv2OVdxS1hS55+8NcLRJ1VpztS/nfGdAFAbnTc19Pku0i9SVAlnLev0VS
iQ12uTUlSqqsy1XYTSPdxUeXRJEEQOThfbzh1m15EGOizEMQ+RYz++1cDZeF4XumMBSW+FD60yvR
NZ+je3zNBGGYKulcfLjDd4HrLCMzoqmO1nCm9BqwHGjzvd3jgiMzrVyx+oUgO7nUitQHDc8IM7dE
1gYCzdHkPbGlI/JwBF6iwBXPfLYqu1Rf1vL5rbE0RB/OSi6EHpqlv4fi4a0yBllcNpiXzisA+BiH
5GZSoEnN2/XKcRvPjDB95axQCWue2/AV07Y0x/JGXZPqMKgloaaWEPDXZd3wGQOgZ5oAIVCdPjxN
m8RTST0xDmVNMFe37wXt2xIp1dmJcFFXfrZQENvjnQ8R4A5MWYR2fpZ64kxYKeng+0R4wt61IoGz
rd4TNfJek6DL+FlrCzJvrJeT8MGhWpw2MRp/KfSSv3agX423iPK/3aTFoY5gSc6WXCwn9JftS/MF
ind/M6I2WvuPBkU94f4HuzoqSJPQeRqeU696finzEptP++yGwGMPCYtxK3e5MhUyBSnLKz8MK9ZQ
ZibQKJusTO30LsfN4Oe2sA5h7S16G2gZClR7rWYN17BYA+oJxbfQbA/lbioLk4SX8f1zNyB3d8C7
UeUpXdvgCiAhrLOkusZKxkymQxJLFlkwQ8n8i5F98SugYfdnXehpEqdZ298UfCeEgvYM2cQpDonf
eZMT6ykos1sjE6nXj0biglLvnF3KvtSv54tslYzSjBPRpRnb3OcAL9cDNEUVCPMpaMOQVzuEmSs7
Cljr7xT0MsNQHtyujgrERue3KzIFGb1yjoeTbJIqw16aZkkTK0fh7Yi2jgiNrNszewpvRjInsfGh
+qai9FNeuXb/WJl4sS8lgghRWjN1Byvk5pv1gXVvgU/QdXQNZ4ZqabJwSgPobPg9PnpvoLswsOa8
JV2BOWmcyAgKEGrupFqFawQ6eMB89DAHxxxSL12n4S1cX9zVcXZ5fIyYQyfB9UnTgBDZNKdYXVo0
gdcG2T2yNKn4XUZIDYY+6GUJ9UZnFHimhPX4rLBtyFCRO5M0nryXzCSFEJ0GTHMVD/tZ+IpvjPug
Q8xWWY2lqj8lHF+Ow4hcQFZmccRWXj4MbqKVOe0QNDT5mh5PKrMSEpKe/JsgvObuq2K5YvIAmEXL
LJbZxx++ozNEqBNRsFL6uS1ZgVBxe/Khf+4BIXk0jun9jQEx/vXysFn/+uX1EMf9eYqjCvrxtDSC
ll+T4r0g44W3yv7fY7y3YDTBGdKjNWdWE7KndWDEeNJK9ZdgX9re1/I73VHcKtATTSeDEv440N3O
6VrrCiWk1Kc7db4LqxEvG5DM4/gjazr8Ws3rE0m2p9JXjYW52nbCh21V4J6QF1UiPt6VZBBNLd6Q
FXpiBY85AUCDbWjY1PbL+Md4g0OK6iFEEMNMgABfBKQ7nClefOmb/Xk+nQAkMCmGwkkWWriuJ1cj
Vs4O4PwE2IqfOI1YQwAXS2pKePxEL9Jk6LqWeRWYkoyiYvTs0yA+EFMI+t6e2HOIIKGEq8IENY9s
hTioMAk/wDx8YsEDzhg3aSdAgIcg1mu/Nv5w1npYUXsv4mdbw0KU8mJP4bLzoDmkbrdougvUESxE
4nxxY12hqe+1Y4d0jahY3t3z5lmG1cJFwXEVzuN0lOIhk9ezIxWUk0lNM0GvUZqHtleZfW+mQHbU
Da/ydxV/jtqKh0TvNqOUV+B9ssUUqRBhjj7XB94/rSXH+YZEmnHGi9vYr0g21PSr5S+pKBVJVxA6
XojZYrzY3KRxJL2V/H5V27xpJm9oyHDW1jrl2B7ttKdzos7YLgGDfQaQUuQyb81BCxi88vFPEU/q
LjaE1E2hcNDBa/OPukz88buz13CqdoMKB/zyy393FrqU3CvzIacL3L2W/xOeakz+1uxzSqsFogeU
MR/77cVTAugwX9wxrTzPYG/8Nv9hW5lsgKMKVlR/38yjkzik7p16VtnjFrKJ6y3SluqLbyxm6g8d
BjAAHJ5OrSAquqYqxxJkXC5rYDwnCIvx7uQhd798wbc3/sgwvKvcr2yKq3uQe3gGTNhyMrcG2tlt
NfdhNVPrcBKbVTVDbiPFZaigcJ+XJboNHOI2l63AAmqsq1QjJPzYlfSXo3JTzWX6gN90kk3ggqzw
4pAxhodpkzMr1ZD3jyPK9rK7FmdXnqXEAoiIDH+gQsL2HzB2F0lbB91+SI/1pxaLn/PnxJMuUkDj
HPtGgUHFPRjb3QNdL0/OyPK9OxXd+yrWzm36s5vINQPYU4hWit3ER+l4ToILeBrkow+fxecdQirs
EcMp0wGnTqwfzUxSdftreE6XreSd7t3f4TQW9oSeWwyVfW8Gz1JO4WOXmj5bo+kmCnFA30gNX/k0
p3+GmZl9SzPbQvkFQXK3xS7kfjW8ShKm/lb9HOJtX8DcX2M3BHHSYxKSFMi1l6T18EfLYcOLxkw1
R5sDG3YiuwGvqAfJ/C+9NfI42mnDiOiq3ysoqrtKtW9LuVwJ7VVjIEa6mDmatn4X8RpCuNCA1YSM
vuRFJM1hjMElENwD62vGLXIcLmv3HCzPRl85IXvf9jPDUhMFjep+62YzI8RQw3vh2GAANZR/t3L4
NQBFZmS4dtnIIXu1J31a1woVtpZDfsoSZYyE9Rg6o9JSUWYLhSNlm2d9GkHJfPi17tpoipwL66x/
Bgs2GnhrSa1UglvhrGQF5QnkRdTmsqMPgrqHRQ+ZpOjEYYwYC4XB8qbUWq4rrJi6SeEVAAL+Ixvz
QLTLpk4K3dqEQKDl7w0bp2M8XaeTDhtpU7v2SpNbXNWngjTk2SK7nPBtWI+TDe+QOvcifeayQUVz
EJBOzN3zpxqccyrc35IBXw4XL+wrAHC1z8U4aBQJyg2makMa5Q77cuUjTNlsUiEkUqsSWSePLJmG
f52S1UW7FDO62txDjth9pnzqCGefLbHKSLe5clv29nrs9zPchmbmjkDphXBsrlhYmYww9x+be+bH
To0PQIYN7aYvOzZtjwki2lK6HNyC6tAJQpMWGAWoF2n64MZ/IkPTiogbYr9Bx+GswFleHfEiXlnA
MoYzisVMdAitSG4g5+q18yFyJnUcm+oDi8xUBEL1fFWW+hCca3Uo3/0Ou1HGb/eQUFEMer3mejGt
O6dQ2RGmD848PvUkuh08kycrW2H20U95SAbObvFjh4zXhkOXDwc347HemU9TH6/q8P8orhGa2dJH
S3Sy8u6jO5zUxmTQChJADsYPkaapxSJlMQQCDtc/Bo685xOJg5qNx1ZUDPLXo5dhuj0rrDKN68wp
ykPZgLFGOk5NCe2NOD0h3xd2V/9nFx5ZR1GI8aDMpO9rT4eh+Mi7KWwaC1fldKjfteFW358mXwUE
09/i2iN/9t6T5f0aF+W8S/qnTYrHFd3M/bG1LciDfh8/wr/9pLjsMhCt/0hwsIvmKxmdHv5adSMO
6FhF8IdCXYu5SUrqvOuST/ePJrWJ95g8q4zjwylU7e9FKs/sEDo5OiMOTT6sWRYCOw2P+0bj6Lsb
ceDqnWmevuU1ZPcLCxnCNPtyHR6hyWppV3oGKc7gCqWCu8gmqJQeVcRpmZNP7MBAYn6UKVof9zfB
NbG84NhRY/cHYlpTox/Cf8VXsvvmKGHa8/ACb00ovd8RX6iudj489wgt1XfuSf8Sa1ruQPkOPWHu
KWInT6rIPxSYdv1NU43YZYTvsj4kaTyy6fbllv3E76X2+FoRpPC5gLnGCNhQMi4EyzIZg1sEwX3m
e4FftOr3XieEInXfhz+jOIaSvbMdm2vnvIgCCi8PkinT0iYWRU6lKdeeWJZ28unwHnAYcspWfDk/
TTDQru/DmC+1bugwzw6RjQi1ZL5yg484COnOImO4BJY0ymYjXFSVvB8ZKd01PxVezGH/ALC+YMrm
Lwn+pPwrg4oUh4/nQRIaWsTCKAN9gnvv1cX2PrzNTr/2T5AQffhCWSoNz212FI8ZaiwJ5lCNO3NO
T06/ef4TshbfUR401+wMizfpoqkxGxF9U4puJTlus0gHrwhRMI+96x23uwHjgUcaStrfz21SdvQn
jN+gr4ksM4PgdkkjMV1FIIIfU+/uG+SrmcdYKc3eE0fKPn2mt7eQJWVukdhB/abL+VuLtD+kIO9M
khL8UchTDvDiZ4vMyykcUrR8WnV1l6nsREbbUWZR1qtr0ZJzi7RTWYu3YB8NiucJ27TFF8+WK96L
qWXoPXnF9BT97N3eU/nnvcTcaSGUITFTeYGSLfVZB3vB2HCPy65VcLVjczHOwav5M8KUqPpevfap
UYrHx3VKSsZZmkKeATgMnAOSF13P+vhCMlQDST9n/ABcGNuqID171UZccA5XnK1z0vOA4tiVI+LZ
zx1XJvPpz+eQ+zjXoRm50lhvprmMaNCmWmgIPZOABuD4F5/4CU+qfkaajtdrj+4j6eubi4vQgbeH
j/FwiZxQebtzSzx2wi6PadLGNoAXESCW9Tld2LtIHG3d3sxCdKPN7SHOyYiaMi5hewIKBwguZXDX
W6b/bvae/sEyW7va3YiXG22pRTHN4mGWS1RRv1dRIY6PYZ/IzYzQYVVvjSuoXqHrStkYRcJqZXl+
73EaA+EtfgBElO+jP2G3hY2BdO8vU/lyJN4CFePLFKJuBMT25OZ+/1USRV3vZg9ZFZDDAnhwtKrS
zhUgPr6d44Pbr0dlB0zG99PGzsEXNJjtNiFs1kYwyo+Hdn1L6f2g7cdfS84LD8lSmkYoQwXEadMX
1IejiidRiDZ3s13msl7VoOCuRuWzrX/x0vvdyyIh3vk0jw2KSNklZVDHOeoRNIYEj3UFbFxAglEr
b5B9sv7ichskInUADd8tP1Xc9iZIrG+LCO5eYsN7PHlTybsQ8In+rwgW5bz0JHkwe+3iWiDBCzg5
0+SCFAUPz6WJmzdaoHtU8yIN09+HlTDM8FO2q1OzLcg0VGpTsxpE+K8T3jV1X4AtaMRmTpWiA5tQ
pPmwZJotZcWZx1tFqr0AW+HHvHnL7+HUoYllqmJOpmZDyG90kp7nQCfN1ri9pJKXyeyJq5+1pCpX
G7WaQxqxQXHqi9/nT1CT8bmiibLOyDhenq7mibsfL9wRvvuVZDwhkCh5Lp2kGEEyy8KlNpjrFilx
1E1HZORk99YncyqBRriH79KYhr1AVHrgprM7VNmwSH6Ep8arY+dUVI5csv9gA62xIaSE9MvksMLe
Bax/Y/WWhdwTJ123rc90+jkTsIY1EHaT2xQstnU7c+FKDn94ijxChmiDPUp6lXtadpRxMsoBDiuU
WgTSC1WF3zE0eT0OzuIDEttozPECUvy0ikFZexxwjtKBh6lQPeLU1bSzS5wNnkeT7YKE8XCVgwHW
q9u92klMcueUGTeZk/h7lIpZAGSd4OfNerVSUI+IUBsHAIUJ7mP7n7lnR0nZF25sxcq7BmPk6+i/
KXReeTFOX1In3/22C7ks1UWGuwbuxKM50cEL9uKxaACnrI1B1NCyFp9IWf9yhv0F8IkItK9GG863
PhZ2xMQMv1MzOCEEkWEoY6MZwvhfURb3FyvYA29hjZGdRfy0iKURdGSh8RO8t4bxpGCbQhE5JGE5
LY68WTYqkAJWSlnToarOCT7MnGWBXgQSdse4GW2FPpQ1eZ9A6tQ8uXfNZCVfv4+CqGr7CRHy09qd
o+ROuZMLWYoVn5HSKEnqhAw9E+s28BIFgzkhNC5ZgxIp9q/0vzHqthFvgK4sY0Ik/9X+FkrRZ0zC
G34YI1Wrx4LIER7Cjd8GFljJ5q1Q65gG41VCpWiCXL71kgZzYKhl6iv86EqgiODny/n8IfHsZhLj
nRD7C26O2EmbYaekFBggTuKWI7ZiQDSAFkEwUL7iA9Gyc39jH2H65XMVCBvF1UcgSWctqNKyelca
ReBI7emta86rxasOlltC0gznrYNYdfSWrTBEMrsU5YQ88sXWcss+6yGkl4rbLdkr8qJYjKKADXWL
6hYsGAviS2gxvjaCfkdDt5edHkUYKn2hP1gtpjCTt40PapGb1K+gNeWgiiQ1aYM7zG2hOnvHJx9u
be1iNsMafOdsaQUUIpMH8jw9pEx0yytfeLKcD1tS1pJdk4iVm2/gk1RQ3yno8cfME0A0MssAM+ed
hOIP+uJHFZ5RNJAwLIRXT+Dtvn+Vw4gEy90e06MWvFrRxnkBQlgPridac1auEbxv5mQLvMjggqh9
DwhWpWiuBc8+owFGPr/Atpq7oNNdviahgBFKMNKzTCLNJN0bMDv6Tx1fYAUFqNLwhlQ2w1hWnEQ2
kLYgCi/iOht6vlhWcNLWFhcHFw7BW6z1g6KrRTNNRvk76AiV6+XNkb2nHCff0t/ZFKx3RLGlSpUO
wPgBeUqXy0163e/ELjMZrUYeHPN9Q+bfWONIV8p75X5gsJLd6Mticfe1QlrT+dtyX6elZ7YYxJNL
zFMghNxXD2zep3sIHlVLIVEoAA/sEv91jVgK6wQvvsZAfCIfCHmLyCh83EDsP+yowZheCmAxCQ8W
FhXWu9fVqt962c/qRAM4uqYGXja2Y7JVR/OpHyRT0K9izqQnR/2Vl79+gWAa4klU0dVo47svGqxA
fPEcalwQAeCm3NmZcmQUH2tnHje5tE6n4rHxDAiMXewGSSnYjBzWp5JRe5gmlvN/iW5y78wRj7GY
BW26yFhVyoVK4p9zvPh/uxGYeZZmMTQabivVqi2k6/fgRdMMJriK7rvCuXB5C9wcafHA6mvLJCvB
TykFLDobvvBEZk34SQNd0cKU+3inrXPnjtHUhozDC/lME7nWQvKuUNYWrtmN1yCGO0e8xTuLHcym
HJrdGnCEF1rN+zLqVFnZTvkf6ODT9ViZUjje8x8Sf8Zh61axVsqmOGPpBO3kLj0QUp1xJTfF2j7E
eqpOZxR1G5xaqq2Kfy7B+ZENLRkLeLg0XHy8GCf2rdy0sTdi6juhJl9h3YCfMhTRB3/2nxl5gQt4
yyQeH1SEfKdP3viP8MeEZTqosFzlyTNJJToh6i0qkR2xH8V3smzHUvWMJHORhMXguYHGaaldv3R/
omKVJc8kcWOMornPPgvCuhzjo9Sn3IJVn5lratqx5cBIi2n8LHrVP11bcQNqXl072t1D2jk79rdC
Zpjz8zC51UDCK+Ds+0JjyHPL0Lgyt/FrHocu162HRgQx2HVHIEw6QTLFWZm131g+ztiyEaDtS4Ws
dnhnSAcP5+WU7kHcnrombIF/9XMcnyJQz0N8s6BxUHtseddVT/OCI9OxhCVTvtshNnf9MuegSvqg
H4QgL0nLVKOlDufVTrAx+mQR0rrx81Ao9eS7+RhaZnI0HvaPh2bO7ptLAMwJaja/kIESWOwJs4bl
QwcbycY55C5WCFg8YYHwwrMdQdYDW+YoErAmrTTHIrpRiHcgMv7aB1UmYK9QFrC3XhuWww55shgq
+IV+CEqbPliu7u2BX7xWCC/4M1Q7Ft3ktHwkmJ/XcgdufJ1mtGR3flK6Io8LRYzmSKcNuMiyU4Vr
rnDvNfjywKtnHFcwhTTTrfhJbfAZHTgtdmSc2nMjTvv7RrJi+wzNbY6AIOPYKMEqd6ayuCgmgvpY
hDEY1hXJZAdfTHGUF8gsl01CTx8O2dqbd5xRccMRAvd+NX19BqO9KznGceWtd87MtH+JUe5bIVsx
tx7sEw8zHn0UCU44t43/5/LSgfw1sJLN3pGV0wtF/jNIRv3z+jkw3Usx9SOLpKj2bMRpJpJHZMXY
ZutqQ4q/2OHik//UEl9HHXF2i+cLVjfn80RvTcpEfowXpQrpZALUooj+DhiSwM3lSfcDnK3wsqHe
jAYdw9bWXSLuehZjyDxeQVfOiMc7HqKr1aQ2TfsUxCz0b8ulRnJ2pePTecZZxuXbuDmzL/pjZw90
GiNetNI8abuaJSyOW9VCPMcOjEidSPZuurSdkCe+RNj8aJXXsozvcoIJn2QXNhw9OG8VuyazcYuK
BWXEsQJo/axXpPRbJ4rsbJzApiUvgu/j07STa3XCjXgA49cZV17/ij0RRon86EJtOmbqnOUliJh2
OOSrwgym6rfblXNceCXXVFIPfkyroZ0jGdnBcxmHgoEmi3nx0570nw9zUmwTK0jc72P2toGhld8z
6ZqeQ0S+2D45gTMhoeStyeXgY4D92hdQeK63Gx95IXwSYeRWnREtvTZwMs2V1n2gsXMCNipBobZk
8D+xR8EE5Msyp6SfDppjWjpXoMI21kaC43670rQcIfAianxdBRzwFJpugVPWpuY0mJwJdjoDzReO
cSuS7Fu2weiioA/EIyQPUF87xyUrrgKayzmtG+vQ7MB3s1SugJvVS9GQIpuCyeYjhXSGjC7NToHm
e6mdvyl288FGO2G3t+vhY/wnzEkNpVX8MDWNpmF7voCvi6qcQwzaNYOPDB3hnh13w97lmNwf4/u8
vAzFHMCPzJbGHIV4v0uU18FfkkgFvarFFhjxhqgnM/UlO5jxPIO6KSvzrPDT6uZcRt9nvKrgQijN
wZl40XXxpr+5ggMB75Rf3RbInBzcfOanzuqva3DkeM65qtbmLJEU/q4Lx9zyRQ7pf51qfx10Atz6
uoUo1vM6OOOMbiJmKjBjQ99xzT8tGLXUzedDWL4vfEzZxKYwZnU5GEF+QP3tJJnr46PWUOQOOhAQ
l5UFG3Sodw2IdjHVM1a3q4sCYULIOuCBL7eNgxTwLD1waLGBaqqL3XF2S/yuWoaxoKq1P25qdf39
TKQ+YErrKpAA330gwSdiNtZIrd/YJNhVdjhKLAlY3YNNcii2gsjKp2QSszIqWMpTC+ms12forwSM
SSq/ZaVCJdXhZRVlwSSQ2vZ+oTxdhGVyp1v2bidSFIuqzB70YSK7QlEgCVkbTnUrCjLhwyiKUD39
Ax+TGaLCFWnMFmS6FWTt0RdxDCYt7Q1KPfeYdlOeNv1Gn6Wcni2cApkthKpQSzz0EJPbu+qQaNa0
8cHts8PFDdlu1EEcFwibVzqtOkqkXtz/odkMYJ+fyhHAnhmjM1+zr/dx2YIor1KoN/xNOtKUNKXZ
AyDDKgvs6YPzJpOCFlAwmch2ByErCt78RxLXfc1Sp7Na1JFY1tbTeA2n/GVGX80UgjCW1y2EYyS4
VeeyPVZsvPYvnSoNv8h/Bme+D4q4cO1f3D3IRAbvXOEORq4HNIiGJJNp0aLP74beP4jFABvhykqa
T0XsU0cxxMyj/T2goHFdsmSdeh1R4oFyuhTNARi/UMShYSgP7MCzq4AA0W8DUJu7tLrAVyL0aSA2
KP2MlZrqS0Mb8Bn0sFhSmgr5o8Wbqm+4tmOpTt2292x8p8myLfNEHizCLf+HX0ROP8cgXTv6vGGe
DbUl6dyy9btIgnTHzupa8KdjYafZN4xTXdeFzGQBJsG9Ea+r1AkQcPr2oe6Y+edjYgeXI+mlG2Ds
yvXWnMwiAoseBHyyIyLDfT81nk9XDps8/g2BdzGM6xIQH8WqcsE56sE8K/qQe/MFTLQcmxTwvC05
eNA50cAwTL/W8Bl0fbcpxPYc6VCk7FvonMfsAXe1MGGOtOssFP/40x0cOzuPhP/J8JMZXEohtxqn
exAhx51QX7EQtCAkrNtDqRaB5aAiEn72jea85x4pRiuOHyNPowuAninDtWyqtbwdYCX3PaHfV4YD
EjtYPlA4aIzZSG8pdRJ/34X3MFMcskqhrnh+fMUY6P8hk9DCc38Xpeg4/uD+UNIlHBVA7W67ZxQh
lqW0kT5MYoXhM/3XoJhUzinnOfLVJlq02c4I9QQuWuSPhHRwS8LSx6o5cQWtcwCT6GVK7RRG9W3i
uD1MJvsZF+Yf2szfaRSSMXTQPcWsB29ZqRUMm/8sXUTul/w8591Tu5I8PDg+tuuTPDJWdIR+oEyG
bnpx74mxQsNNmf37ytJPxzCz0593DmLpRiU+ImuHOLsOJyc4ree6rpVo9ryaQvlrm28ulPd/oDOc
CBHIxzSfJgIxLdxJSVQz4Gr/XXaFtSEeWhjbdmiBX4juijsXpDEk49YtO+7Yzy8GRJiamNzHe+b5
kQK3GuHBei2yOHBenQAyrEiPTP/pJnYf92eiV6g32HwPmdfG1tr/PDTx8SvbCyQxSuClk5AWkAoU
RQQSWZUnACGPHS5Hr5PKmGSNKs8mBiK7XN5K4zXVTge4UCZhysrKcYhBpB6vpEGxl8qKRCeTwICE
fZZrVwplcyKgrIGasa8r6Uie7A+4EbBy9aswSqcuNfnfncgk/2Fv9Im9WFNM9i9/gB9SQCE2dRv/
/I4U4V+U/W6KZv7XsqhnmlWC/fjJkNFUfPgGBO8efVXbpFYhNGX0eUWtg0/g/b0hxV7hT2WQnOZ1
bIujLXtGXZsCOgvsD9X16bC9kE9AN/FG3x7OpzrCmRzj5tt3XYyPFV8T1pCFYRjAAF/BH4lgERlJ
2xqBDEQsRqOJhIu3GY8dRHFNQYdmp2P5kltYceus+/JfT08CE8rdxT1QRf+O0lcjwfwk4QA2b6Nv
Lynpo/NKsSOE6qaaw6b+8K3LCYvAq1HmL5j3pDWhc6dhczzP+O0qDw+biWP2CUpco5IrLwu/TR95
mx1TThM23E/ajMZgozJBZG5moLiS/UDeDXjgTgANPADQCS7FZWDArEdpKmrgrsaN6Z+dwL0qOOgG
OtSFqq/ZTHsJotstfLBxy/Cx/OY3Z29KhGO+s4puLLnA1AKoIBWGOpy82izNpf+6v/lcel1bVNT/
pWKCHWnsB1ZNNvBTj3sp0/0AWCV5jiu0epjsTyZGAlKdKzqowK5WESB+oYD81gpGtMfw+LtRq12R
Szk6eFuMbSY93b2aK9qXN2+GPOAIfDpiNfy3sIm4nQw8vGaLNnnTg8znA02Wpn0F3fzEpXU0FJ/G
TU6LgiMSyysLjOyQQIKtbO753Nfr4nfJmWBhP7U9XN6sYeYz1nNRR/bPB3FHLU2Ct7XoJukvwtqx
K/sJubBpm2/X07jC+afu/WbvJlRt1IV1QPlYb0czDPZKTM3sj5lrFcYbJ1RB2a/jw0elgMR5HYAH
soW4hyrEqpdmiyqdprIMMX0Fdcwknj7/erIYifNKYIzb6t10wzU+Ux+KzrIyHFm6QPDjHKhANdbq
G0mj0MOPqMklDq3I6XIOmpgV4Qy2nb7BxiQz1t9XPRTbPBtHiLKTqvuTg2MoFfoq+d+GJrn3Mto6
Rt36wg+5jPiV9HyQpLD85XzpP6mrCekRNNuLhayEYTHKU1NyErmmCYss0/4pNDbz5sprBQBZ5sfT
ue4XKjbpVAKxfFmY/sEzfnfrmX4u6xaSSx04QDlmVgYHqDCgFY+h7wLKXXTd8FKoMfOy48yacmZ8
6Ejr4FiTRDL5ALBuFlUUHC6EHLXeUyEYqr4XOxtcPbYncdK7b1crPWUnxLHT/4k/NKBz2hu9W9/M
oSSHLP5un6nUy2AhGM4TkB9M6sjpVUu15Y5W2aRQCAY+jbgKjkk2ggxCSViGw82nOBFJZiNHQC0j
G+885u63heN9VV8GprmiR1nYgUrYOpiCBVl+eXXP4YZ6bjdBnPzg81nE7DurRBWOyBTgwotJsypO
TOa2b4Z7SrSx0sCL6+S/amswgw6/DlgdwMqe5tIyDmNR6NKLlwQhRaYuEfKhbXsjnoIDgtNpvKze
yN0WZjXSugdTWu4O9nqHerxQFuslVKEW9wb0ulPC05Jvl6pCx+nVK5NbgiHSYhi+hML3yIeGPBOa
srl7JT/ILFMUY+F3EpFlPBPDoU+T3RFn8B9R0iUOimYbE09yUBX6xRmDafeYRtvKDBKU914swpCm
Al3RChvhoGHE36+aJb52SOGfyW6IfqV3koHj203Bleh95KpUHKOyd77mzgRjcrDynVplA7swTbaN
9kALY5rxx2b8ygHDgM7Fm4FjKqJFK0Bt77gtG6kRlcDSZhAwBT2r19QQzlmLA5mBD1eOnqEkVqMA
O20Kgn3ovRt8wbh0cJ2Nbfn6nBF7RxP3T1Y78vYW5BoFNhGd3bqaiSp5lwvczu7MEWB3j1HaasTz
fJg25UPEM5GtgvbxJq9zBEaOaqoK+eBYpxgQ0mm6MMvODDHtMUhDOM/BeBsSPP9I8gkhJwGLbiwZ
9gbYa309Gy/GTKPJc/t2zfECunm4XYzFmkbdzPU9rkwGn8mEiR1iti31vm4Mdkz7f4xt/Rgpa7Uk
cH3DhJQKh875W9gdhyoF6FtGfXvi6CPR1J/dYUz+9Tys3ULc24XIUoL0XAjjWLLqI+QnO5kW0KAG
hWpKiljy13VvurrgzyOEWT23E9E6o80tWuV+xayInvuweLWasRpHRPScBwxooXQoqi/sXxG1HPF3
SlpTd0xpGMiyDLnO9qQT+EnSYLYVg2gn2cmvDnD2gecnlInrb1KbmaUj641UxmDfvDd8oylXrX7M
2duuefHUYv6CPXoapgGixt6BFxZB1CtrpqDJ1wu09bQUqjcAWJy/SVoTMGU/tCiaNbTclOucqRfv
aPlGH48SYTJG/mRt/Ue3g2Nf6vFze6jsp2l17P7dDuA0ZWuLXeguDcVvsPy01V+Md/ZYuh1r/PZW
JIKDLFhsY5mPbIALOeTmWh5i0PTu0f49cUZjI0yziL1M3034SgCKXAt8unz1pr9mb9fiD//uMdU1
tyCKCRd+3yU5WKaOhLUSgMhyfcry5UE4jdvxZA52mMYneajb3Cgw09hqeq8kDl1PN5MFJg5RM/+r
gsfqhHcdiXiSNVIaZexwnKquGvcFCjfnzRw0PJQNm4bhts4CO39mdrLzTLwyDuaUy6w37PzIthtQ
eyYJqv83rzlHdtg6YkeZKnvlD+Gx09o4lpXI21rxwD4ji6okbCXcL1z03ZI7Sht5TR7jCOyDva5w
cEFrr51SzWrtDwfCOZjorvqHg9f/cXS8wFLsq6wkTdiR/dg2oXh8TRZLx5WT8yAn0rV0ACXwk7M7
WRQNIEGM3kiY/qjcGXSL39xc/nmIolMrScLVK/5oocPkayMuwBR4tbCkeEDexSEgObYY64czVaO6
GAyjb4kIcLguZdb4rK/fw8p224bDSNgz/gFqbM74hjIOH5HLXgjlvInufGdVAwAY5MM4F551t3gH
nYls2EZDMUZLNrRtLnxkp6byyfchN6p5GB7RF3PYFDATq0Q9PIKpdPGrvFoxpORYcXOqm+E24s98
BX3NtUCBKptAocmMbD+ALKOct3jM0naHavhZB9BcLdbw/c+3AFyvydeZGqIoP+dOIO2LHNajJCjE
qr19ocyfVONwDMVlJMsBksAz3GvRY0TnO35fVbKHtHa3Tw+bIcQ0UNEx0aumjWsDqCVq5um4hTIK
SwrIC/LL1ORvbOnMcDgqd3DGjzA2ln6X+QgGxeicskyefbb4IUClEdvxVdnW7xtgEadvidFmXzy0
ItLIDvSNuOCV2b+3KPqUO14jjdqzVxUSNeWN+F2Y5fWHgKoxxH8gtMubltDMjmjyIbZjLQw+q5Te
u9T+nJuk6wlpROfM+CyD/bUvS9bkN4Zu+WSfmMtjpigWEik1wBZbAU6Ttd3Laepq3lvmSXcHb5R5
GeZiuWlOkDVo0/9t6A+STGUbLo5mSDLeTB+lwuY7y658vVst3519HRrGmgweAradu3SNKz15+gQF
pOwrHq2E5TYE3MO6h0A5e/J7HhMX3GztuDpEziL2APXXHAEVs/+IWYfjJGSSFpO84sIfMhnB7dm3
QrIZqMc9U65XMrr5p4M4RR57KiHkt10iIKWFZzBlhac5CeyBKAujh7cVch3Ozu9vLBKH9hLdOmIR
fAHXmShD0AsnIk3gQMBx61eE0nzRLT5HAqp4kSrM8OqRqqUxTypvMWJCOfY7zda9N2XVtw2Wo48w
IsSBvpwq+ZN/rPRQ1ln+TbByZlvv6ndm5msRzo4ZAhFCnTJwYu/Iv0yeY9yJ0deiu3YTJe6Mg4mx
YPx5DQ/xwmTPY3lYmkKE3P/ATgUIds68PTiyiu6wvhD9hWM0fnaL40Kb54xmdxSZLpjVGTFpU1fx
GXyenoClZYEGpBgW1zeyBsMDJtq4Y8INF/nOyW+AvWWyoe8l7U/HFG9PPsm+YGALHOt+94NgHb9e
4yA57uXYEnYMjvpbS7F5/lYN0QG1W2ntb2kHUKPbjdznuu3CCi2PYFQYaqNVjCUqLUQJ7BJPSXKI
zWaAHisUggjrZcE0MOrM9wd+RMPkOEArLdZugI4KbGKoCuwvvrv0E1jLvYguBwPT1fi2Ut+G2DnR
TPSX1immPFzQNSayHgIbMIk4h6BY0FZav065NTBMPvdWvL4ParM5BG27cwX7nFcp/i07lDFgtD9i
C45P8srZYRulPabHzxAcMx/0zIQSTlTYqw2Pa6KlObzQsRCleg74Q5awiNKS79s9/sKiYC3RzK2b
toDHZswvgQ/nDbDQxSm0HkR9X7DkQnAje4vY1Ynh5qXg3FW30eBeDSG2wDzwWYCyjaF/FvE0/PS+
j63XYLNSL8IhMWGDn0hmStsu1XVFNulQ4s+EdJ+bGsZvZDtnhNdmoIsNCikS3m/NIHRzYYfCKNZ6
wQHblEzWV37WyIl1XBydJ3pHnwwdVgQ0JOcbPkgj3mdRPuCKi9LzkGWm74x+PfANFfPE1HdZM6wr
ydDvTjvl55DJeeG9KbVAn5CeeVWagnr2X/kbUuUHddulYJvFQ38RQpvc+Bn/uVbQBtg8OsIZ0eM0
dygm0eAcEfGHorDKgJYCwgzHU8k31cTTry51UFsnQruQu3RJ/wEo/FNvHfOFVEWLpe0haHtNhy0w
eG6EK78uElqhojAo6nXvj663Ed1KCa9N9Uxejn74Q8ientgdzbcYIR3HfNSl304M3ICda/sWCtcs
vcR9GcJpDU0DOWtcmDil1uECa4drkXp2waCdMSTiFduUzXiKx/kIX2wqGKgHhx/lkoRFAG/SFaEP
PCjMvUIB9gIcdxbBW3U8lFQuTbYSBFJsNm6+kulRJrRjzWnEcgfUNMQMJbLvC1ErD3JpCMm0WBYn
ql4qoSkIsbrd+AU2AxYT9hMb0otjmTPHi4bXUxeAqaAdbBLZsPaFEEzwK7NEy/ExtFH52mXtrc4S
dCNcmZYX/bkfIqKsGgq7m+2oYuinT/uTzZpBYy4pKaF/o+Ylks+8y4GRr2E93UPxcQLy6vKjS8Mq
CksjOV97G31eykHyR5O0vw45nbRXda9D9TEfU0vMDwEtGppCekDODZTw7dPW0MGWQbc7M3DkrN+m
6IRJbz/OL9xSPWo+xBzeXQm58MjhKaJwdT9oNjBlrEDjXs7g8qzSrvSpmIl1/JNm1R4YWLUKivn3
/c8EhMC3x936q2ko5xScS+LodoG+hnLfFZ4KVVuoQYc1SwDbrVk0DicEEColab3bAeT+dvQ5dpoY
/CtpC8ceHwkEgLEAwXcBH7y9hqfygAHC1VbZHFwS6C/9nUidy009ghk6T5sIc66bGkt/kpneLCDU
/YFQfzEUVNxEDM7rfhgHS3WmYVe66D3lVWGmblhUA8zyOsPyMYJTj4Tv4tkAihdE4QPEJTFoAGZs
qUocuL3VIbXqfFYT0xYLJnnt1SSMP8CpzHUbSlgaE8fjVpb5nERBTVTY1sqG9RYwtPqDeYuIA9cE
/COwb5L85iwcsK2UG3mciEW04kJSeijENLJFGNGIXSxktrJyP1COck5hjcCNSwCYlgyaanLIXT0M
4EoZmzUMADwner8CdbZELZSNKy2JEF50+nBL8GOCHTWw77x4m6JL3TUkmKtKHGiCsmd0DlXCcr27
2D5byRv1EKOSQ6fmLQtDgWSGOmxodsgK60FMxFEPRd55YZmrCxKOCl3jZ4FXEj9v7WRCRmuWIYD4
TEZZV8hIjyJ3+9D8lrFdixpEst74gIRxXkx+WNknNDlbWfSQnim8TOV2MbrdGlz1hoHtYg8HhRsI
UqhctdfaBhmLT6qM9GKcWxMqBmkUF0Ct8d8geGc0bVurABp7Y6iZpYAnH7c68WgbAo13PCBTAPxM
YLNEysXnVWhUfUcOyKdx88YPmfEwL8SbTcykmk+qDI7lBa3XlO6UcCo7ySNDzV2R5GIymIIEX0h8
+e5c+HcL+gbVFwVbe+FjOAPbKHPDSQZzosvTH8d3UcatS0k1NWgXQ51NSLstNe5/OXexVhTi/qgN
6GirXW9yLXQLQUTUNhHML/z52ajisc64jj9sc/iy0s45G1MtnQf8OcEv1Xbq6TUJm/IA2S0drV6J
/fGWJQ108P4PKszRnneUoHejlkBAp5Psa21iB+ZAM7jI/JkyoDS+qbMncd79Ee/25nftPq8EfSPB
A0U/uv09T6iYplRlo1I6Ywli3Fd48UxhI+AyssufmGBG4XtWEhyRM8k0Fb8FC1HYDDZchc/gRNWF
PQfSEZ8TNd7znl241GvXqkEVERB0sG55i/8YTsHDwC5Inp/INEVFsouoA/Mm3GUB3wXcVxCD5JSe
ccIdmraDrwwERqS77Re9JWhbRtokqcVuQo0CsHdxwOEuaS313uqy63LEViHAZhDn0Pefm2xbMK0v
ItQc2VDnfAdhWmeDv3k2kjlSrkdOmCZfdqBe1bCk2R1Wrhytnpk/+RzERL1QiYLdhXSVPN221i1C
G6sn6BQzOM/5PXrQYHKjMDn9KM/KxpPerxDq/zaVG0QJ7sADWavVNT8gP3F8W2rUVO7YWz/oP/db
i8p4LBzASc236ZepnWstO9yjkCO/+E5S8yONtvrILujkD3IwBVEl7YEWoEQg15z9kyHOBOuOOz6J
sH/iLtjuRVAQRSltwkw+hk67SGjy7SYLZzZYANO547dB7vmKBGCayEJWYPu3hxwPKNzSh9J47NhS
RToH+fQtg5Dy51rr6Grh0NKBb4mTnwynkV0bvWzDDzUh+mZChnog5PYtnaE9WEjdJy2QDgqFPq69
UcS7CC1OOy0ljHCwho/9rX1IpTImVyrjvv9UXVs2yc/umwiTzVm6XdQrc/blJTmG0jgOzweAoDJi
A84OEuXmGEN6t5SWpzBjHCIBTSEwCNIRQUD8VwHNYt/q1550C+mrK0mMLjQwihyQDJh0FFUjjvJT
1fzaQItVrdbVP2UDwvyAEi3I1yLBen+Z+0tZyC5nxQG/5mnARC7MgAIKS9A8uwPJsImgBKC8yB16
n3DVlzpS0/PaRNMpN+tJf+5UuPEMkNUiCuuhbyHNnN5/s1Q/V8fg3d7pxDJEDJZHZ8zHB8nvE+bu
ihX4brKgLejMiasyWfZwU11BfKAVtk7hOAlBeSD2ctNtCtaSN2pOqshNmwljOBeoM2V2q7qRSgHA
RzHvRey/6HLsdt0qukzmLL1qKm46dW/jlsXMiW/U69qvfJKRqB8ON7EdTbg45hPB1O0fi3hn/BaS
oJ0NrBHGJ/+yv2Ozp05+VgDjTTVP0Q59FW+Tf4+hpZRp02JZjAcHaQGCYAK3/0GBMak9w9s0sjPO
fhDfiM3Q03ySQHsVaCyPYTpbYMFX8DBRJkMoic8cLxy7rhp/jRjNLm1Om+fkWx+W4CwMfJFOqJoF
CNYsG4uzGQDbo7XD4JpAigGgLWCpx5gwyH0z+UksJqsX0D/niY4YB07UEqIHvJUllZHMfKPxJFzC
z1CUdduS9SQTkEWiSebLd+pewt+Wg38FzrCQEsDtzqRlpNP8zKlZ4VX7CNBHQ995YYyhKazecL1z
y/GaFLnZ1DjDdxzZ+zgkqjKlVRc9LFoz4Yv4j/5+9pfkaSLy3t6JgIqWrhIRvWfGYybqsl8ID83/
M8KSNQgiiYR7mOY7b7XZrbmw/WhaXcxQxmy+dHhm84Kr+WXf45fDp7zrO3wTP3MLKuiaNdZs9DUQ
5IfZsPEKX1wgMA3hEsW6wstkBamE99ejalWgzt8sdWZIrw1Dk784ojR2Yy2WAgZ8cyTFI3wiiSFu
nptrz7tqievRkvDG/Mbv59Ra7LjIZpF/nbwXoG3m0+FNhzwtq8UoDEsc2iM54DNjlXKPwIAWSSQS
sUqXlUJ+IqtHNaXWWU1yrnXK7K3TCaju4a8rgD00gI7X2KbSrvDnsnbrEs2ZDz5fnDOqv7puQlN0
ueifMCxp18ISefq7oxOlBgNxCbdjoLIg9KK6rqMcxFzgPpMM9DOeB8CqeB85VGftSiQlBlXTrk6E
Mp9E1PmgUeRTPr5EzNJwp5Ec4VufnkxvQO0kzVJy+kQmf6rMe8TLkA5SQzv+/GQMivDGlmoU0gkV
as5+yEs6TLEelg72ibVEou1p+75fEQFkTiKFQJA/1lYD0YImxb6Od1l+NoV889WxESVrEYjKZf3a
Ufk1zH0QJLd3tj6lBrawMhuBakgbcATuHD0CG2rBL1MwbiP1+IKXBV83H7mhG4mZ/bsDkYzMV1Id
tMxXyxrlLQd01ybmv44EK3845IZ7t03qMEKZA0HVyTYal1VzpFGc1spT1MPsSQilTRWxUGmMhZ9p
5ScxxlrM4OQKstvcqbDCW7cG0/k/+W1Rz/D66ROwcQO0rczH7fSp4tZvhgmfFH2T6kWBWB0mOe5H
+VlGYrTiyN8XJ2D+Pr8QYELuArgLO6YH6ZgyWIj7C3z+6PphzDg2a3aajTYBR2anZ690aHH9ZjNu
keEMuAdAIATzHz56+NGu/dNpaYSIyAsnD0fAITI+8WZevTO+vHmJ29zqs8Y0RrS3t473JxGZQPTy
31xS3DvcpZWJ25Vog0JzeJLeR1ax8RXCxXe5QbTpSF9uVi1YTOB5Qt+eI26UGPpKrLQe3lLc+D07
iuyBUQL1ymtqOa24gpDKSnfoox2oEPZ5z7olvBm7pLO6n1XafAurR8fWRDJp/6A4WnhoO9vTQku2
MAIkNJYK6ByOttfvPe0K98CkskFVAtxE6IZv7Vb+KEjU6MEUZabkOArIICzTnrwqynZjpI/SSdRT
NoihItxpF4y2P29vUPcacqckWnbXdPwP7bAw5z+p/2R4KdNHigTGzOHnEj5eYSBLYJP38Yo5tehe
IszZS9x+lH4Llay8GjhuiJVQ46+Uruv4AmXC5EkRYKzuLyDKXmnN8cu3YqtuzSHQda/NNcB+mkXD
29NFGB+jI0IpBuK5Xa7g24q5MEsvBO0HLhdyJqy3s6UWfKSqVRy/tSgUopoaL5qycMq3fbIqTq3Z
PSH2xTw8iFqJO9+MmglCMum+rhNNCtYJ1nIXoNzDmr0GkhDfl8IL6SiYhjfbN8Liix7ww+vVDEUp
3DMlpSNwrL6KOSQLhBV2zK6pYDe6e49sfuPLVKQWVTnd3smWj7C2jvZEbxr9WwLlJC8An7D3nZ9K
sbXu9yxkExbb5UGljHrWOEx7AO9kHuAGQkWDaTaYWsGfWthlPoForlvn5IIRwD0YkruPFbVH9XjT
6JLiYN/G39Q1ssMWi0sunEQNgVklKL0bm+dmzbC9IQOVp/BZ5lIrFhz8WzbT81ecsZg54bd0tvK5
IM5Mkl2xoMnXc1HIQN5vGABfo2WgC0K4gigUDqCc2CMU5Zy7Z9KwnM+hNckS41Ebrdsyhi/RZxKs
BawZXrJPbnvgTbpKSZlOVSI57MluSCmkR/d9hOxZrjPP7cLQyEaLTRL9Ow1nqcEub0t0muCor0jT
ACMMpDQjk94eE+gqBIft1jYFMUPbW0PEr9Qim1/iyFb950B0gCqsMDXgr0g1C6kr5VUZndVNbRDl
N5apLxf4RVjakPfMEuNOQE0g9yK0S1uxLfFklUAwgM19SCUlFEEl4sR4QV0ew0tdrGSuK9v37ZCu
qNQVjWa0M48EO0fdNByfNW+8zjDZ0/QOSdp6Amf7DD92GqMEh0vhSzOJkhwoyAqaAc/8Foa0Wdno
3MwkTP5G08Mjwn/QDTvZFYbF3C4K1C/vySBoGwqEJ73zvIybOyrO071U0kY0mvlpSGfLb8zXGV8j
v1iWWaAIMhhcVpmqsHDgiii7HpjXDrDyiJbvXido/zy4/zMnVQpOWPm6EBlixD/mH3/vhHRYBbQy
c7R/3IS2SROl1V3ohV1XF85uYEXHhD2t2TZrrdEO518wEY/wYvMCq/jWIFJktpI4G0Sk7Z9sTm4h
uEJswddPT+7JpcMdcJQC7tY7xfaHUaSexsjys4M7i+QZdsiP1BEhhjxjO94tttdk2kOqEFnTgt8g
dB1c1gFhGNSgymDl6AZr5SY6aZeoaPZ7lZOcaZr2b+Tamr2ZAL8za/DuTDf3bw+z75YBtN4Igq6z
9mkQxK1Ba2YAyfOngFypnquMsTOZlJGb/TvYyn7iatM1G4NIcxQVA2+Qbj7ou2Gl8hcNtkGilSFv
am4dHzRDDRW1m6ZHVV0BjaLHn+kTzrx+JTFv7Qy01nEjnFIqor9awiiGLxZdtBE1OA/zbBB8r27J
Q0Hr6BJsqeHn16pmmvdRE6lrKXfm5p5CZA3FLpmki6Vgmj21/Bdop9REnupULM8bV4q6YHzSdSxG
/94NgBI0h9mJ6GbFFXMzGD4w7cjoS4BgbOh3bbG0AXdLFgb13EwesFefNWyrZN7AN4RHkzDOtZNc
sGY/d0ZVMVF3cRwpAECmhgaWS0gTSbDCeE/fnRARlC7LjdnpUUmu1jfSnWvaMrhtFfikKMmRwKfU
3ebZnqDio4p2NOBFsFc8UW/UJEAe+OO1qNoydUGM7MjCwSjiGH/s3j9gr6D0OV6J6F59bVQc8//s
lgYTsASoe65xbwEYkI2y92peO6Lzz6voJd0J2ZsmCj7YeQWqvdMv5vvrWr4GwtDLSJl77fc2A9a0
iiFxN5Poe4i7R9RHIRT5GX+x1wmFSSA0p0Y61hCvmvyBQ6Uvs0bL6OZQTKanQAsUCkf9c28TveUO
SVoYkCny6LMBDNAbgnnYhA0hZleckJClDicmYrBnSUaKSzsjQ0VieaXtwXoX8UffW3M8cYFSLjsn
/+akZrmmPIlcEB2QUT12nwGgIWHCUCNLmQWcrula76Rn8cwAZl53fIyiz2kxde6qWYsfai0Y9KP9
KaYPFQ5s1NoZMWZr+V66rWq1rhhqv6yyb0kWbXZj4YZyXBKlv18XYUKyWHrV2c1ZutX1vcY00/Xf
w1M83Jj2assVHmOtZ1IizmYsV/1a1N2d1ZGjY8NfgTc+bPlUSTzZMg6Zlxd9mSjnqtk3j5h+ofEf
61ToHT+wMW9Fx4rQ71M0A+YvWnD8GiCsk6XhOvJlAHBqevmQPJzGS7C1QH+zD///8i1yO8XAjet5
O8gMYLM/3un3bRL9vZ07m/mHCuIfFFeY7L8FttDtMwgLK4KN5Z6p6VB5AoPZRbRm7DBvsWxkUQJI
jifJE4IhSo6YPB6BvMleBN+wuyExOpZtqcwUl7UvCsTrP/Fhvlx0I9f4ANarpDyPJgL/qOwrFuMo
kNKZl5Dg4+QlPp/O1iI72Z/kOpqQpx2TUzAtk1jTlk4qqCa1JB7CtHHCr2fPL5xHWdWlry0bs9M0
7oG1tVJr+2yHMuPw48Q5TrfK/p2tRWcD3u2PG4x5m5/Kw/5ywXiKXHhBjccCnxPYqm5nIq1UD3Ju
0tdcyH+XLp5oKTsuFRCXQzJ72iSSmucC8fRjtyOF+POCjJM17iYsqbSwrqgFdtMr3QpYra/DRaAg
i5REJl8Ae2J9cf50ifbdOSFHn/+aYYH3afS6vcXS9Pb+pzDKaiF7xKROyiYjP6NJljhhZJ0kxgMp
WEdQO2XAxm1k1S6n7DxLn+mNrJgjpqiKny6fSia7uTUQo1ri2Ptj/ye4jZ20s4hvx+59OV1+rEvG
JpjAPwgjQqh8P0XXMYVKbhOM1nBwffD+h3Oa9xnpWqbXb9M9o5bBqhSATIFFIjQ2ITqVUjIuh8bX
4IvvL2GE1nvN0HPQHIo9sRn4GeTDuJT1ZFQMRzuGCk1AaBN2UMekTLzAa1t3oxzhOt/Tkqlm3dC1
bVlrYvuBgN1lF+jdJLb02jzPE44fOfdEOJJz6dgX1mQj2+pJAQXuf/eflZN6njgePHSc/ELfY682
jRpSlyHwbOLy0+EY1Fdci5Q/MYGKarxQyajYoOc9aP4eDPc0Bh1TJzVm3y0gWTBi2+70Nfsyt8Bm
1eIiUAku/REK5a8yGLurXoyL4VhY8MnsyzrNk3KbXZ9wu4rfuDuRdjJtbYQ47dURdENv4G/+ld+Q
o0/xqKHzrPxiwLt04TMFTd4csEPnF4HjrTYGF0PT1Z4NDrzk0EfFRpjZu1vjiefQbuXVsEblxaLT
WL3hFtRDgaX067o/bwwfDQEbNsx2xUMMCVxAg3np+/U8/YT9EpK4pp+pJCm6M8r5qN2xJPVOdmw6
dnXovCdeFhETYkSdWlyaWgfhLWjlijOLLYjNqiCi2WOyBtNBWyXtWjt7xVH49NfTq1gxtFOcpN+t
cGzSKkuLVC51b8wUPXoTXTxXxNgGVzhn9Yyp/zr1L5E6Gg1RHKtke4qZsZOTgkTDwMOgPQkrrA1y
Flf7umvYT1JPyMP84sCHDkUnN+7LPuPPTiyKUV37Fsc7hlzXiR4TSUhX5aNbGyA7xP/ogiUZcdtp
QXCHesPdSz18tVKeNFnyrSp9h6aEw7pJPR5pQvl+vL+j+aUeTA05KM/sJ344izL3CnYtBB9s5v6J
MANdIXZ2gZkbDvRHWbGeC7skQNc2hLXyHgACrJOGvMsCR17j/GXveS4c6S556S+qKXIDk3XtykbJ
a2ENCnh3uFRCLYsnjAHc1HC+wl0T+RtjYoqPk/xK8+E/pQfQkZwWuCoaMuWMbY+P+z7xTI6plrsF
o2AVjUjgyL8mlzH1P0fKe8stbzw0ZM0APDzr+xrGDTI2a1L3Va48ajXTZKEjnwVrC2vIdbbANsuc
F3gNWGJbVCEb7uvtnBLmpKZY/gAPIot6C9PB2zF9FpwzlCRvJS9Z5CVNQqie182ryJ5j0t49f5fZ
5BQWqPI0bXgnaR4f0OT87WbIy0e19I0UNI7sbtxgJG/RenrBkMxRlN5GbE8//Sy/tjyCLpA0QzlD
gNL3rx4ElCzJ55Tf5/ZwDZ0wT+xFPP40z4fxev78Em43T1rgdv0pf7R1w8jiq8J7BA6/TNhQSjNN
VE/sTLOEQ8w/w6nRJ2kAEYsQIx2guSHuPHH6vs8Ce5fXCiVDxXOk+dZ9s7lz3qZbvMfDD451s46m
xvilfAU8bssGMVVSyOO/98XyLfSeoVbCr7kSOFPzaFkQFS5ju0M4nRDRwIpkZuWJGF1xD82eS/EN
rGdZVuwt+3H8Lr0hul+IADNR4eXDE8GihohN3a173mRDT3DJG/2+908zugp3o6fjQErVyQhQC4XX
OwIG6/+hj0Li8O7FEvf4LRKD3B3A7ZlnvKIGSD6TL3szPF1oimhsFfAV5+ocGMrLZ2+IC/PnJ/+s
YcyikG6eyxORvNLZWE961Wklz7q2+3NLOU0v40rh+ZL7eGozWmoGUcjqyptMxoV/Kj9WmbD4Fj16
ZS1S3x8aQ13qqb8DFvWRMJFIcaLIYpQMV+DaKoqv8xuk6x61FNo8qrxUBEUEX6p8jAbLf4Q4s5FQ
YZONabwlh8E+yZzYKSJ4zew2L3Uwi96nYgPgpkJZdCvsN3DuZ4ujevZx6+PLdrNrN1lL3UfGvXrF
Z+prMce3MLYT8uo5J2FMiToL/qBRsOQcDlFn7vIIM0/kKGDx08o4z35ItpesueZHs/ndqKyvpwkg
bxT785CjXK+vNIKzrPpmqTvgjzOKjtwIgLp3cPAFTd7Vn5un14YkejXwXw2c/n7UDQL4hdr15H9R
2tE7eGAcVWyrGgzMfBp99qzXQIznZxRPW0unmApR7G4gILWIfAeV666qtpNPGta9Pim53kaqrYrK
25hkR3gjXGWvKLFZeVuCF8unM/NzpTeMso+5JWDU4OquaW13Lob01d1d1fNRRfCxuiz5CP0ujZ85
FSSSZOBnYuhwok3/gbpdOSzz/YI5RPvA0RtSS4T62Z8NAbj0TramPA9mbVq4MRsvyJxiIkAKl9pT
pzdPZptbdoUX2L3otptLOssyL6zw+OuCD7ft8lBcPOuBZNTwChOWVt6HeIipP24ktuE+seTYnZDF
3WDycd0KeT5l1df2U2NECIFtaU8r/ULE6yNUEZrEXs/SCQ15w6s/TruGD/niBw1L3aDDSo8n5d+K
wffychKbA2yxdIsA7c2CI9xCt8nM90EbWTnoDNw7KbI3E1g6sKAXhQKnlDZE9T11C9JgXlpvyAAV
WFScFXskZ0EQnG/BQJKal2Xkyn29V2nFeh3PnTi114DmSvYLNJpuVdgO55wA6lWDATXycFELGJSw
VALDwIFPCC1uP2S2ks+rWzOmWr7pb9WyLavUzWr0d40H3fHKYF/Opv5K8/uu6FRWzHy5jgpsJkPC
QXhRp9iiiNCsVhBh41mU9AaItzzvCjkGzl2g+2F52+NHhvsj5fomzk31XOaweijRJbrDrbDle4Mo
8E4c+zfyM9WBDzHziZTDeDo5HGymMOD2yN/jDRPJHtePdV46IHyKdMllw603zyuMSIKZvMQuDVZg
erbKRuk7MppYspPE7mSDUG7h6ro2HBKMh4zJtJb1kRZqe8QN2EGH76+dSj7BTr0x9BAP9iQJHw9v
AyruLluL0iFje4CR8PlvGZXM7Nm4bWr3uoh4RpbERwOs0vFfz2oVo5DsQVSeMvTP22YxO2IQHmqG
xazCTzK3JSN1MM1Sb06WifVSGaL6NKEDs+lWBmVnJduJnKZZazYmFuT2ugnndBNmItPFkGl6FTbO
vlg+uV0GfaFCk7r2RFGHQCR+4yYarNIAJTZHSvMk2WTYYTO8oIWj/8eQL0oHBJsPgn1pa6wl8Ukz
P3dBvvOK78VxDLgtXx1+D7zM9g81WLCaRNFtwNmjCY+rQjT/Cdul/gwEFLEHYnxhlMR50lIN/VP7
0n3cKLS97SpbIw3UUvh6ICN24au3KGzMvvE5JsNWL6ABet9DCLQ5yS+obNcWLeDyFu3Qa6ishMfa
AB+n6PyUnr7QdvWu/CG8gi3SDVjjKQ3TOooBrokTS9TeepzFhlOUaMa/hOPUfI3hEHaBs3tyRxgA
HZlZ5Rg29Syf6410kL0J72IJXdINzeLRO12dKuIAxAH7KLmOvJB50J2Dmz3tmo++Kwi3FAFuA/wg
EEDd0sCOfJZmEjOUkQKTvYTUk57c3wNpX4gD6Xs/AkM+nkp8GRMqidYKI1TlfRUsFqV9ByXstGwg
37C9R+Ywb03+AWvjuhnioWaW0gKQLEaqmCoEWtzHIhdV51/GFAWMs9oR8UlKeh4fd40QQbVECexw
w1Q3/8kqg0P+dmtuKtVJLIby/bQQpI/ryQH0NiZVaHU/Uhu36UgXfs6teBmL8zaFIieGDIS4VJEN
enPT91XlrWebceUiN4MYGr+HQ2r1yUK/pzlZ7h/086AKeAL06+96v8I/1AvHaLqiGzD4TLCKWgDR
TcvErv+eo5NO9OaMIFd+m8ZUmldFn455Z0uN9FgCIKQ4IVrso9u60h06Q8f1A0C+2iFUtF9622fA
ZzZTjhk2IJLEi69Pfr1FVx3lnaPAKwKLST81ehI9A+6C3ux2AaJJXjmXZthu8aNqNUXFMpZwQjKE
mIeNifCgKg1R7Qy0EyNXzsGG7y0rsq/vQiZfwd+xKMFbZ2q5RYpAegaQCMR5QAAFbFNyx2PCiOiX
WZB+xeylJ5q982JNFPOQx+DvGMIH7CMUh9H4WRv7invgydJwV24h58QBUCLuYrG3ll1ND0+rmW6P
ZFWaejCKkpwFrAU1P2ggkzbT0H5FUQfwRkRPW4wnacjCvmyByz72oI9qGg5CP5mEdilBvqZlngR1
k8P43kf54lFYpqczrgVK+6b6X0eOOvOaqvKAG/yQKyHJ3QExPcPr4oMaXMnsCLFicrKkybEgjgyf
FflRhdaTMBlG6pewRexIyNYMzah4zYMaV64nqIC5FgPHJiFK79wfRZMa+y7i9BgpS0Ga7zxbX6R7
PTqm2FbS1qlCRYhfEFY9fIjriI7ePQnJHCrA2ZpadwwXFvrJVMpT9nkR1Zcnw4aQ+m5x7FP8G8uj
SBsBa56yguPwJOnoRHU9mW1uwCNQFfGFTGCJnLl6LzahF1ek8uhV7Un1+2jMGmuJ8b2wAC/agGTC
eEC2uyi6FNW5QhIWGsSo9NDwIdt4tBx+qFk3Urkd6jJ7QXPtrp7ss6xJfpuwqZkfTsPGjEDQ1QHH
GDZKKUrrAoF/e82nH4V1xV8B8drs0Md44iz986s/OP6G8GIqy0nCjvRmQlJzgFVGN9jxbP6GsMfK
0qb/zP4DF7ZhUNGiZNcFN4pI+EsnM82SGCualFHySU+5E1JKO6mLrm60cCpI41FMhrUVZ+UKq+j2
R5DvwAArvjJefRUYEDUFvp3M8qBPpPx4PdIuSKJEdylQD1olcw5SyCvaIWDLkmALHfCy3AEa4Djp
wlM6Jmg1q5UeejEpSsgBIJpl41tedb1XJwsUkk1IK3pecAdeJEAfb07R3/yehEw1EuqetmivXXtH
4sGeAymNrmW8SiB2FUkbigUoHvglEEUu3dFRhzvgOiIyr6qyfXCNdcyyzRDTf/oMSD+A3ngPBwh+
wrxpq/gfJkaVraKGQ46bficDYa3/PGXytvd9XJGezE1/Vyvzb8tL54DTVVYpNPR8TLHSxaXyiTyi
ffaO1HJR0SBT/qUSj7c9mP+nYWpumPDP1B54NKid9/KUio4df2U6gwkzzpYlN9qfNL3zvhut53fk
DbyYzeL+r3H0Tpj9UiQZpryVOEWmXvBX2XDFK9MEvZFL4W8RsnikZJugQsb/CiX1le2Z3+PLjs08
CepLmnmmKjrws9il6CCxvK3Xvfl/fuwpreU/s6iu+fJPZwg1Q9lH9XP/btbbh7EC146IXSfM9xP7
w8nJKl3vFOVAmIllNQ7QHi0ghgqPc7QXa2fsD0ZGpGumwCUgHlpaq4OLFIiHKf5PqTBgynlZA/kv
QZ2Zo+GDeODORcfvdkGSvoYHBJAxvS4ub51RFpmWirC3EiuWwB+BMlrJVbhw/7yRcXbX6eeJ0veA
XCcwgCrVSeu1MpOhO47M11MJQIriPFDbcAQlNFcSxyaO1EjNvUxTo/Jd++k90fZfhcknJpKVLCSY
HN+arfaKS3y3+evAmyoxhV5ysraRNcAGPAYrWDA7QoO79lQnsNoZED6AUsnwcYQmgi++d+7Kxkvv
Jd0TIZrXTwk8uz8B8Y9BBE2EH08htG1ZA7yzu+LEPSNXdvziAHL/dux/758gE1KduFqKXnE82S5q
8D2XLA77LFzuXaJoiq95Os+ci/M1QDIeth3KNjpbaAu+Ym0IwzEm3mrACBcfUjHobC18eG9wD7zn
NDp8xNbDjjloloohkmWu0xlEq1hF1NcMzbQOKoJtQChe6rSekoZg0hAOvB9VjWNE2ZTzZWC5C09K
RtXAwbloYz8NCUTvgw30GNpISEc1fPI6wGFyNhL01U7e6iq93ameo76kvkGbP+Y+i/lWbu8N6Imd
4EpZcBfuIdum+LJ9wCico1hmp4VLR1nrk5xpI9E0PQJBvj8I8BcxgwhRD5JmB9XQ3GcqOLYMpSta
OmDn7JHFSKHRkyq4mJ+FqnNUXpHc5Z6ITpVe9OzaBfIrCCkB69tJ17TQKoh96ZWT24F8gl2YVCXR
M7tarMJIBNReb8KAqAfSDh4beRk7gDxQl2DAaPnkVyxTz8Xb0x/iX30TYVMbsI2GDOzzBLkNcW5L
7FuWOZpnAK4eHCZzwI2rrz0jw3YM/zWHWdO68IoH9YB5kN+acy/MSTmf+r9bOfEejmSm5PZVZ+jd
nre1nnjPVt2GodTUwqkCU8tsqVgegsthQ2kmTWeukACWhPYqmIJQNe0PvItb34u49iH6Q5HV0eFQ
hjgBxkfabC2dmP7XL6LU/BgtwIXcSp8r0ctIAWM119ezHaYc32SRZqKiZBOv1cfPejab1onU+fQw
WEtKx38LFoQsZYKQUfYKcbI8bx50TxuLRrAkUaMqrfYZ2h54j0NNkEtw2tR7k1oftr/74kfR6QEK
FY2wGDiY/bfMqwS8HX9wxT+FGj0ASMu1v7ec93cI1bY3H4pqHW3zo7vpIWfLCPSlDOTsQboyucD6
JISB/tbSgesQA3zSuWafT1/WUdtAHaMsH1smQnKCwJipGHDhCwuLw+tFHsZSG/gcVhQzkobZby5d
K4guTnhGzSniNdV3zY2JudiYFzzDl4wokpVx6zSg9AS8HWjaIzR5xuUf0SvZ2VBdygMFjCDdqicx
IlexmnWu6gJ5nht/BnkCD4XgZ6pg4sVsvHS5Qygpur+O49f8ddsra3jKKrbTekmIDXe+8AoPB+/f
vEFV9Z2n74KPKf0HV+zJ91PtxOIVAxWLOR67bK15KORt4j2taMX7GoAHYbGjfDYwf9cGKBEWzVcZ
nZoqlMG1GQsORjj+dOj9ilhcjT6vqrXftMkBbauS+3Zwll7Zg3Q3pLVj8emOW8G9SKhXzBoFTe0V
DE06kuSSTB0oENx+QftYqN8YZFkzhAdTZhI7xtl23RbgHk79Z5DTd/TQdm3fNR44kp+BfyDiFoih
+iluiJrhUKvwxM1tTAKgveDMPqbIP9uTuhi04zdPMsIWafBT2jngekTPsVEI2OTwT7UVQKaGVU4g
NVaK+enUrBlQYnuLRrcozRUp3o4CttdV9XF0qpf2gI3+ZB/sG1qwnIhbDqt15QO6Tyh+dAJzN9Mv
kBmU1i6WyY7z59vbyIfigHvouRswjjkJ3n6rp8I7HVVU7Z3MMlvImRaeycDzX4vOmv2zQi4HNPkr
vjLGXqajQWVBqgZikOl4XrMHpmZGoN1Wy7tfjM2veFqqs0g0VlajEhDTnK5uOR2i+oSipqb/HKLu
uLCwHA7gn9ocWF7gqFOGpemlKS7z/nmBPkNnHAGBH4/aiJ5h4Il0hEX8FU/1Bb2zpnnpRUu6RlIn
RMLCMpGwhuuhUjiBFoKZ7SZFwnsBg8bHID75cuYW84LiSYOhz0J0unu+habadHVgCzZd98XYD10q
SGByeeKOT8BdDjVDXNq9SuduaNa9fSZP+fATURIXQ1V0GJa3qPViVoUW0z4ZfnfOI68xZYzOMbwX
KpmfUBSX2Qlze8S1Y0XKiyT8iqG6M861Vyc3CMsEtf+CsQ6JaV84bSROBSC+DFJGgfxdj04qcv9Y
3u8hvTIc+b6dTJNuqj9FAXXoL/cogryxPMMu4qGtLFpY6kbJkYSdlAxKuLLRphLvBmukTA7x8j1H
AwKRhdskAg+FypkqqjYTX1Tjyy+UVidCvE9uNPPIbps+U+7tuc6RMWmgajbYlF0jqNda4bJzfgkw
jIu3pmWQCw5dCJ06ZZ5fs3hgs8O4X83Z9lW3IFWsMVFk3Yc8tXF8ECrhGugVXQ+3Xvwa44ZK6v3M
wy0pT51vE2CAIzE24p2GNWbroOBqzLuOV4yBCwu6W5nhHbzNlm+ZzsskOWB5iIeU9VX+O1R0rRJ/
WF0+K9P/9u1eDhULNVlgc/cBNUU8mfCMhu7hauArDqdclgrqlAii6TCR/AFXSKSbZ0xwb5h3EA9t
WPy5bu71wpWgdRZT9kZWxVS5hcq00SWrOXVC7FdWKmkksq1vQX6qDmVDxgqbTg1hVdTwb5+f/zYw
bMeYMreR8lU3jBUdFAvmUYVe5fZyuamkq/BcsPQmtqn2nwPu1sYYNGJDoiQPrzg9z8ih9LQ4rpiu
xUBbeINJkddeo4CVbg4Bsrm1w7Xrq4wkUT5RHJpb0KxfFvmrs7nFeiaP7iSU4ntGgc6SfdWONAo3
ddd+9ORePZHl2mtlB0FhGRTkKfwQ0/1ZYCHvqwTczrHjd4I+NkQCyD5idjE0dyxRSA/AorjBt43R
xbmsPwYb99AK1VMo8iH1RWmHllJMGH6dA8Cl9ZpLpxxFsjNcLIfHu90va4u70+8q6wIe92uYU2oq
q1flBeUfr4GykSrMxMTN85hLFbIGI5wFl71QjpKxoZSWJ453jSSjzgE8tHWN5y2wjsDmxu+5yJfT
5GF6XpjkfyFHUtzcmoAvHRTjkmlOjDv9f3l9p0Kg/ot3xRD082O+Mg8Ow79hG5epQDFtUE7cvNyz
mIiW/XmhBJDNiJea+VRonBUCpMD5JXWsmFejvLJIJhHoMeE5FMjo7lWqK+oYTzPNTLF5IbEu0C9H
Qbl0g7ry/0iwmGV7XFPEZ2ISJDK1mUSrvAk8Z/5Ip+GSCy23TKPqJWrY2j2k1HZpDJsQW52RYJLc
M1BUKH0gtZPi8iwczdyKTDGWwGj2VnACfGyYTOpzBJV22QaCJdvgtFUDQMZUuZkE5/BFwm7AaOOz
y0VzhSrMYfTH+jbPU+vbJlLpoq5lAukx60JzvQOYd12x8AqmcyEF6UlDSxAA/sHTAHDA7o8YYEpw
u8d1qloJcCAEGP0U/tSQew+VwZgUkTKxxPGsoQzyBV/VRv2+KSqmvo/RaBdrJ6azy9Z8veDKml15
CIiShPz+SCRkM7W+D0MoEBzrjnX7QRG3C7EBnkJ1oGTnCr4xieg7jxAIUWPkX8RPO3E50BlY+hYb
8RMEbvfwbgRk6zetHyyjMzUcGswfAAqEb8x4BUC9GCqWAqO9o9GK/g8tLL5UPMzsK9hkEi4ME4HM
zlOUDpYKtWGR2DkgH3p+GIo0tgnOjtvj068quShyieH16OM/Tj2z0uo5aFqCO5qLxJw8xSWn+pPt
HDYaO/LrdAoNuoO5Yavsd4bSpVZSTZ3zvPkKjVKh9EW+2XIe7VvTyYPbdTH+2tk5Ng/5IjFNF0Q1
lonTCaPHziCxfXj9Qnbgm7n0lJvQ/5YnlJkVaTf8OlsAy/DpqPwSys9905AcGO70tj7dnhd06l0s
nWWelsNK19m1bM2tN5aufiT6hdjBYNJP89KxvBRZ90V29up1I3TZ0+nO2f6i500pdwjhAFFDlDJa
x1XVi9ypt3S4/XZ4AymUWHCTDXQs6VrlzHzuGelzOIIBz5tjdQcD5VN86Kn6rUGNy/ffqSFdXmvX
e4+ZM5xNFSwChxwxlK4A/X9+ZnTxrm16X9Of5kd5CC1ARyRJFJrXMA0yCgBlEdse43djJbqAG/xZ
bcvTlHhbklDSY4B8uUkN2Ln7jQA3Cl6nVqY15tezyY6rUr2/dmMg+KQS2rvLAU8njxZIY4ecRdmf
pqVJECSKp0WLNVQyRaJD2DxMmXCxVFlDDVwEN1Ffr81WcBW2YbUi8obJrTPPmLBU8vnLkpkG9dmT
2D+/bwMUrUmENaBwd24TRNYFIKWeDbCi6OC0YJj1AXy4v/zgghB8TzfjCYtYtgvK1XKjnlUnkXTH
qXIkxNkbvG2iRyRxFOcfGAwEix3AB8CG9yOz4vB3Hjb7LRHyiI/HsNcKe2gaHVIsS93T4uIXYiG3
ytuJfQV44GOUsWHUziFFVz7vXF7WuoYSd1B1zH/W/Hx1XR3AHnQSJVvvwxW1vYCqVIIcSt5yLMvx
4EqGNXZK1PksrDHUDWQCU19X0pBm0nFZtwHEExBrSwYCdubDibY5LUrW0cUsKrextaXAchfGuyft
sQnjJ7A6sHtgKVk2TDp8Cbpaq74d5YToLqcHAsMIQfWY/bemvM9xErI2+OL63jRSMARUaG3/ouQp
GtZQH72Gn4e+W0IV4oBj0NBHXMBwIhAIWMyU7hL+prW0bcl99miYjPBSww7M6ewnXog10a33sWC2
mmcee49HYnSvQpEjdiqOahTly2ctQWDSoSzLhQBxNHHj4ZbrrgrUEmtdKud/IN6yt/sfrVZs4q+F
Z+ib+RvQZywDSY0hzprSNp0YiLIXfaVv3sLnwH4wI7zqx/vj52JKYdAjrQW8w79UvtbWoH11Vbql
zU9NcRYQkFI70XbGo5Q5GPcPtfXavTN6B4VYbThOLREbLnuBLArlOokvUqMSYR4IaXua6E2DWXBz
229NAA6bje+1V85RELWL8uE/rOWb9JQxJGXFiriu4S7Vm8N0X1CYfK7sqarh2VIl9ZrpIebK47ic
RuR6qofnZEnUi6VwIaOfEmCWihJyJst9Gk6x6mwYgyhfWE0aYfFdmwIfGVSqxugNwjf3z0QEaoQH
DRcw4xxdmtCrwmfhFYALhZL9y6cWIoqL5kt/MGH8IK5wxkjEtHb2ONK8TtUMeRXXdFDDch5eJaNO
MGTBOQWRutrhInb6gdCKKCZ2pUAOiLP4CJRP743rbIqMpSd8lmHwY4VCEHY36uxgRSC4iId8N7qC
VsZQOlnv9P0pBq8fvwYO2Dh8Xg7VtFdZW2g8VHoW9pdbPuPPd8yDn+v1wN47hww3zCprT9GcQfjN
9xIobVwf5Lu1YShpnfQ1+HsVFsNRuoh53L3VEU/AmwqYkU4tVqkmj7SWlXh3cgQNPfB0LEC6Sr3B
Vc9ZZEQX5lO3E1m7bGXEdTFhNQkNv7ZoXHu+KAgD5sihiTta9hRAj5+nonDAfY+8COiTbRZPibob
aBAS1qaYPdzWKLPiGBczduHCcuiE3ZG4X/gUYCPYOhtuc/x1z6n7C6eyBizCTkf0Gtx8g9C/TmM0
PNT9XM7gJPNLacTFVXnc9ARWtAxl79GLjl3cWRUd+q5aGcMfLzRsk/BR+l6bu0PpB9OMD/426gUJ
65sCNjJJc5W0pf2PHBLaEHVmsA36JP81boh3YjSLzzNzOI+L02LuvyL/WeJBt1o3YqOewxebPABC
x64F241P6XcojyVWqwD+1XFNV5BMrKgXAdgu40yOc9W0ehK0eHMtZ3XphynHiaxXNs83BzRW0rss
vv8tMedJOgSsQRi7KAQDI6UyYWH02wu3GzwBUkJxPj5JJ1tYltvUfbf5cEiyLUP0Mje/5ul+juEQ
EZ8e4KYcEPLsb/pzNS9bJqW9LhBXGXMLNbMaTukRUZVo09LbPHZIOjsWNDKNK3WjR1sW1ZVtV1RX
RmKIw4v4GoVBBPO9uw46kT0qGcgkgYa8HcV6JixQB0Naqwa7rYmCS9U5fgHi3xiy7INuh6Vuw6z0
2KBm1etU7JHx3vu8cTerOtlIheJ/Y2NyLleLA9dOmi6JC73kjkN0YHrvgVWyHlGin+s75q0PTAuu
uyFBLlcMZkVB0TV5SScNY77QPJA+e9M+3P9KRH7liNx2GrPWpLrEKvAbCvddD7StRn6yV+1BJwEA
UyQ3Ax9YiC2u0ZSs9kewl1W94vn0+/Ej11RJJvfRLNHPNbQKGCZyTZ8B6kdmjXo3HqeTIVMkdcZr
njbzannGZ9iYKHuZPQOvfUfBow+CLxOhyKWDAhSuYNN7DchBXZ4NvRgocbdR7cmgGLn7Nrq6KW9a
c53wlz6QQeWDU3AyMitAT6UV1ZPHrWj1MpYIPtqgRG/hrY/uYztGS/dxJiQ0KDedtciSz5zCaHs8
ticsXlenQ8AEocS62XGU1R36TsV48B6WLwi8vd6GE5Ht4iBI/OyJcC71x17xrBm87GYjZXUsYElZ
kEwJYa2n5Imnr+xMpsTH1Fz9b03IpzN5JYsXE+PKLgJJKUi7tYXG6C1Xkc9fbecy+cv8AscRRhTD
db3+oZkObARz4+r4T9fVut30sHYoPA1Ljkzxhvm+SaCyyI49HkHo2BIwNAc94LX0Nyeas86qosXQ
bgOkF9pFoPy1UNIVyIjPbbJGhpQQcPb6mw0uEWNvRlCzXScUNmyH2MobQ6SVMn8j6QjjVWg9kTrh
3KYA/qgzlN4R+hRAEXtXBhVpjB0JRjZcayLp5BDmays9hRQhTfSQhQEclYoGQwDQwwttSK95ZUA8
iX/+UcC155eq0WSaIJZ4HZrTlXynbYo44Si4qJjKBkoOoh5AOAK3keUwogWKjgnRJ6ZZFrL500cc
J28krqCcTHPaaqtk5TNz2c7TFjsxhnCxj5WV1FwAI8aOGvTMN6JoSGhMEWOeHCF1NrNVz+8vQymA
MV3Y3Y4YDUoQ7bCT0tQoRyZbWmdsVKT41giEv3bNvkO9tOdtsMwtnfLdUgNMvo7Ou49cZiwtsyyL
nfinC0gpi76z1T/1PL1tcAX9Ypqbsq8BE8rHuMPQEWc3sOItAWAg7dQmE+q0MhfAovgTCLFZpzPm
9xXPf/alQLT9lodakmzdHPTPSl3MX0C5At2U2lpFPHqbGNj/RqS+xxDFHWrHdY/E+jrbZAEFIow8
K2fLXpEiugObAheJEeoQMrve0PVNy1WXQTlIwIX8UybvzRiJneO7PGpLf4rmyjMpFnN5wpevbAd0
wsKn9Yc9Bz8qzaJhmzvGmC5v/3AwdhduheO+xaujv5Upo2chZyLC/0+qakSMElVB8Rh1J4xETfnF
Ohx9vKwkZBI5K4CtGH3UbHJgWcBVAKGQZhWBp5TIxuOK0oCrjRwcIrmQzc+on2feTy5M9lP5kV/2
EkI0y0w6ogbJWgosuVQ+91V9uHIqcT5BwwJy5mldhg92moPScnGlLnMAeNcCSwH5gj6RLQxe4fwL
Z7DurSUm6rwcffruDFRWWkJgfMkoxnvtu7VtualaBWyhq2rcZLZx8/HGSZuCkZz+zCSkivZnB+h8
tN/aFZPxto4kYtg92SLdlzB5doOAwr0WDnrgr9HUrqGacOeSEe1BmwgUkm2FsBHiczm2SwLtwq7Q
Yv4tqsW8mHZDdQKTKk3XlOKgiJlcOAm9TLcEYoaEvZ4eskgM55PnHI+aPWKuEH/HXnhoa4JlpkC3
WM5XNLqgnyG5O8XgUi0KbPFihrM++jeghFAEc2FSaF8ro281fEDWcr9yPmGTGGhaT0bYUqml9EY/
thMsAl5fWoTBnXoAuepKcRFtJPTNbmsvWv9yvO3cFEx9YUWwgNsZ6WKQ86Y7Tqpz3sddG7iROTAT
G4lhXUC/vRb86OqABbeDFh77PUH6zUoQIGWS/ij4Up570sKFMpzF60jzyqUk2D17Di+vMQCC1i7G
76WCmR9W7b8Nn1vaNTKxB7U4bEeDHRO9TA5jl9p1l2QI1AVGmv2LjRTWgjXQdUfpz8/l8pQPYmi4
quTbx0wxDKn4YK3q8QN/IDvMA1Mt67DEvtyg5wzHFVO/f1UPUU8Uvjd4RmcrxVQrUI953p5TiDrN
Ui1uSzI9DVwfcpgOSi/3/xHFc2RSFnJBRu+8zTSQzTqfKDwl3bL1IHeVC/oMHM5sDsMQjQPx4nd5
mvwuNK7r8V4dVAqkE1x8sNFYSxEj91KbNpHI0kON9jRTBCiuMRR96s1uI2qiAPBNOInVy8pxqAPw
6j/mJ39kkYT/tdrT9Zu1lnLDxy7q0Ewu7EeRV/twrQljchjOHX4mqe4logyP1DK7/qx32Bw/6tae
2eQVEFU5fhHXG9++/aTk1vVAryyR1lHDjsVAEXmA4FnDQj8916R2YCcGWAwgLI+rJGYIE/ukb55Y
01cVIDPzcjxL54Tsu+QSBCk62TpjlPbJGmaf0N3a/KiGx5RnCbLKOcsUAe0DB1HELiZQtTQze8f5
n/26m7ladj+kmFdinU4vwOV0YInTn+GZc4CRi5HHUpRnvA9Zt7rkx+8140fT9hmmVGFlbL8RSWeM
spPkbrtjLF+P8ReGubkejQXt/orD6Qsn5MVxIANJOFQVb8bIi/zgZDaSDWewTkHkqpVk7YjMcpp8
gt1XyPtLrK2B81BdYQ6rs10wVTTWEH6N+DxkMgTYSP7JEk2cg2pRva58Qrx51x4jcsJP1JClS2Bj
uUsSjIhtj7TbCK4fuCZPJBgAxgW2MRRYTk2XmY5aU4FBYo0uB07BpzhjDd99yI9eWAD5Inrb+pZE
9bAdi1s4Gip2IF6UmCT1jASunnVkPL78cYoStnoQEfNsZWD0z6GVurep6XKydUdrXtP3X+mop3Jp
yhQT+d28Mn9Q5MdWayz4OmThouHgetCnKyjatGDBJn46/CP2YXmklsYGDgzvNz+GEeaniSpJY5Fx
r6Hnow1OmcL4q6FOiAjUIx1BZKgbA12v7ORrrEbaba0Ykh+lCz2t71mixcgzs6I2adSLxEw/Ci9p
e+FP4cCWAu4C7zG4Rp8iDVI/o+6D6Ev20Rq3z4YZtNBWIqztZBKvh2nNeCLBkiLXhOfOl4w/4E9e
82mMUZsIBjfy1FvtajX+nu2PzYqznHp/4eWekZW/bUl1Lhi6377ItyUcJVMOaZv5DhEY696NaGpJ
yWa0mCFbyrmpWNy2E7ZMEFGnXAIIkTpqQlhMOtgqhI217A+Uo/Jw1XI/U76fRQNlYa/42MTnalLl
RFATP9MsHippXYeUfu3jZrgf6iLfFhsR5RsRqXEXnaILSWknRK2jJ8D0YuW/4ypv6z7IXyxM4ATh
UhHcWmBgQOYWI5faHxTmER4glsvTiJiDlyjYo8kHhdMvUfC0Z6wy2qA3NSNqt2W3NHtbmUm2WeGy
3OQOI/LCiwxUyTsxTxJInYWcqHu8ahGe0IV50hF7G07JEpQvvRXQ0oPjAIRFMvA65AVx7Hi8sYu6
Yq9J2nyFGARGudDitezvK8/fsOeuoChqnX1XCpv+QxcgPKA9w72ZL2rPnmttxIEz+I1wkHMQz9bd
BRy7SnklyU/+0e3yLnzIMngP0otivs0RM/wj+wUP2roEZRijJHyz0A4En2KjLIIltiwDX5DvHZ4N
rJQs3hiRXp38WHYBiYslSvGRJsEhwcwiqN54Vp5o2zIKq9CsRYbAoFLCAqu2CnhV0NCEDZ8H3rCv
nwPcNYX9sgfEtgrcMPytW4rcwdPzjCIr9sLGuUjwJJgk44KW7UR2LyjyBINureu09zFjKZv0rUm+
hv/tnkfYcgFieyfHYQRff1cNI55we/ddY3AhOg2N7qnI7xLZpg7ww6GsnN87FTayl7FJQppoREUo
mrORooFt+EpDdoFfwY2w/ugwRCTQD5vxXkkIscaFeFz3HmA6eHZ3/uveOFQNvPncQSyPnN42Vvj6
QFwh4dn02meLGRnFpXMbJZ4jslOH11jpD4uc0Pfbu6ECKxAB43meIrvjwaVhQmOCZS8PgOWwJaiD
8A04SP5VmD8tpdZzWncD2Abo8hxZQTbZMKvXfTf7nNsUcvfQ+AwNPeKr74uQPf8izRvu3Y7GS5yX
IgbDgoM46FH8VFWE1An7sgRGvnQ79iMn4wuaATju7Vrjt+fNXWwSoh2cRVMcWSdq/k/BjRhlxesl
HyUB+EIq9ox9wEGrfE6SIrsU0xhISssmBMqACYAfc6SR1p7ABY5TphdKS68myVJeZBKegkRBJPkd
hVSGYqGA4T0cYDh10IiyiXQodCDPm9uV7TQ6LXf4xDnJX15ZtlsyqAMVeyD4vRIaWk7wJSLIZMCZ
4vM1t64yjm3j+kwwE9wGCGlzKJ1svBUqSwlTi0P9+S2AMeiG8cAGWAXX3PZlTd3P8DgEhWEcimUN
CoJg4U+MBEe9Cga6Vek9dH3tHnpmeiLnqL23+4rIo21MVVxrCehXN5n1MI+ZyPdz6xcHWy3TPhPM
6XdoHF0g5Lrd1JK2IR3JahX+Zw314hLqwfv32LvQ7sJ8OIslOLUwjf5PacrV0ISQtZSl3JmcYMBa
OD4YNUvax5PTb4GmHTP1YqBbAE2stP5+VZYL/4yV5m41/aSYjqcVY2LYm7YVC0PBrjDWDCLHoqE5
jT5q2u1ssfboFoS0qAe7Wb6LE9oXOAnOn+r8KNHgvNtmPROVi2pEGsmFbj3lpulkMWVS0hT5kBkh
h9yFZ5wBeQ6ORgyqK5srOEgTb+eSzTWj4zUib3SwpavrQUJ1NwzwLktR0FuYn7b+PixlzIssLSNd
xPMCoyQnLlvc1FXZtNGByk6RWuUzka6pahenSDfQKZ7pIBYdTgcgXLrRyoPquDOaGR5h7wfAtkY3
D4oFAVlRyRsFInG62dyDFy2+vyWTjCijF3xnP4i/z7balEPl3pNMZZqWnXXDb9773tpz21KjE4nY
ilFPc8RhnDZ7C4pkaW96WbZrTzCE/IFB8tJsKq4YSk3wfF6DH1GFsCqwN9drwDpy22dGMWBcKspx
/T7AYE2Stvuw7NyxBpSoFv9jaNKlf5hmnNBeKxWVj/GhVl3KF5tY5f+nTWd5ankuUPbG1bWEm1jq
ZCC/qwGeA0qH4Fibh2WyWZtU/xQWHs7sWRkwQ1qM0xpsCQq7Wclv5iT2dm8EJKcZimYKre8LvoAw
VWO9kki+O/lRuGmxJUuZDJp/dDgFOQ612mRt6DYVWaAclqGwdUWWv7Ik7OHt9MLC3+rHdJyrBiDx
0QhX8neejs479lcyR+I7BVxvb1Mndz1A/0NhOtWLg31Rg6KNVE1szVzOQjqKv/PHsmQqbFRLZ7Jk
k6IviBS8QXa9GyrhDLnYeUhOCD721NsfD22F5MKB54/pPRirQNg1n0IPjIyok1dij6dmr78/a1QZ
qUiZriIOaeYdInQzno5VtvkSDGIvDXS6RHZFac+9XvydhKXYkHceOeFUTLDISAP2KrWzpqwIlgOt
XWiGtztP3uAr2z84mQR9jrO63lx8kX8awvpAwEYhHI1GgY1SST4Z5310StqG7FU2P9oUgtg4fl0+
yDnBPQ+Y9stUz7KTN0sRr/SAwOesTMu4fkUpqDOcEP0Q1+67PYbUDdvy8sjn22L1U2y1ELrkCI8v
fKBiYDpv2Ek+mjpbRgq8TW0DIpEhTmxZ9sPO3sxDvNtdOUyFNBZrocSWDMOTCIM2RsZNJ2OMVsMc
f+suCTPtop0UAZ819MCznirLiGi7YraTF2tkIRzIMWx69rce51mw/QdrKLosFqMWooiEKoDFO1Ki
HqlgECHFO1R9H77yEoF2n10iMyx99xJKUY6d8xeRGmctQHTQjPwAAUuI/K7waHsBsDAjDRTItHB0
f6vD45sWTEPKujOxguIIdXyKP01U7lJG+3dMFuXIrPh4a89r/mUuxJfbhyQngRF4vV2tv6n1+F6R
VV8rr3bC6Gj3jt8t4oBzYkYjwDmgX2+28sqOnK90apquC+EY7zTWoYrZ9Xo5c6w/aj3rO5n8bi+b
4Y7BnJEtlCQRRk5HuJ8BHPys+ANRoY/ULefsP/a8a7bXB+Sopvv1SmSW6bqH0xz4zekYKOVz6dAB
STgtvJ+CyN8yeu2DXhXdzVE/gDKrwr/BsEpMFFarUCfIwLepzE0UGJ7o7TUGdT2Etc4sC/evDUvv
aji7nvrfhDtub1qq0aQ9A+bDFDRmJKy8hWfn8kTm+MuNjLcESZPIYWU8BcwY/7AHDey28vtnIxI+
tj2wlkY5kMK6ej0QiDovHY74PGOvaHyWyy4kBiYj/NGZU0knIMP/c0AQ9PN0JiESnMSVuptAskRw
Y5tFlFonQubgWqbBGyWtz1388jFVyAW6Jtjsf+8d1xipFX6KzoVpEqklgLKUW91NaAX3W1QREejP
CqXQWqBu0M9xuGXBSRmhvhZZMBhUZpgcdt4loqwIhiFUvN8D8jNgzaIraVlQYG6+9Ss8U+w7C0FZ
ba5BJILncGGNAp+mbSR3g++3unJesarSyifZMNHvAOT48J8kMNhW2Qr+OG5Iop8vS9InSgU4+40p
qlEuExmsNQG+S62j+J6jS26y+73TJhvJNtN3GBIXbrVV8/EN/7Yt/FPoeV8mKW3XwtQeLOXfwhJ9
FK8CcNV8UJDdooSpzxuRCHbXqUCL9emK1F5mVw1aTyE6ShHcF7CWxTli6Uvb1OVcImK0LtCiGaR0
nOSApQZWM00iTrsCDxuWSrC+6dD3y9LA/wX3YdI0C/l/RHY7kqokWOKIly5ysR+4lsEvUZNYz6ZT
IwvKIXcoaxxrfzhXDKIWCYZzK31p+Tt3f25ET+Nqqsv0I3ABqu2s6bOYw5/0p7oGYqIwrFbaHLLU
l5imOZruZKI6t/5MdpCSpep4oz//4+cT6OeA+frtqVS+UMWXGB5QKwa4kYx8Djusg9+v3s/RPFgT
0O79e8nfO9ZM3YZ0HcEhir+e88/n5K2r0vUYqOytDOy1rMRYpsKvbHt9+itn7G8FbvXDa5Nb04cH
FGWpBJ/zTTjxtNhapaoQ68DGF3s9qnGYTxplXyT+cCgsd83i8Jfeu475/8K6GSyc0PDwSlCQqxVh
TdwQTGTU5xFRTngryc9mssdjXtScuOFmG0xRhXBX1WWpYyzWqVz0Zk7U7pHZvoS/d0+qo+jzCikK
pLVCWVtGGLe7TmajKBVE3uXwr7kreHaz11REIct75SCE0vfLN0xpuq8LDsnkYZhfFIpSv46NREfY
mrp1gL5EkMfTXLEsNggVx03oEQjigyf0mWqc3tDIZARHz9YQ9Ylt1bNYyv1PAhioqUO6UFWRjRqV
yMreRL7OislhL9zgPV8M00B5LVfOcinsb9gxWHKfywLMrUzVMDa3UaJWQiSIDdSPZgmZNGNJEeHg
GpPkKzSmykpb3+vhrWSzhHLD+wUnMw10dqopx9JWeTgZtzn1EbfbDyGy0D2nAJeN1MHRElis1pJM
+lsCuEsV1AQVpJWi682Ao0lv0dneFYImCybcxVMAulsZsBI2dIqJBe9kTvZyxx55hGlPn6aAk16r
dM3ztLmVkfIdiIyoP4U4lnIdBEqIQkestOtzQEmisuq0UQeSFE2/nwdVz7r35d+0+TDT7HfglN/P
Mh5sgfEy+TGV7bt1bSxNwZpcDmRuEQjXe5tj0nUBPemI/R3/esVDfwClPV0isnURzabGPeoSnMZ/
J5HIc6hOZ4yMk4PAt8VN5Dpvw3K0K7oTBpvT+mRrVLfYe4fJgWWetEHvCCp+jp/Us7yJPtPAFmdv
uE29WJsTiP6Ul/K7wy3loOJ1Yzn4AVblxP1/7/U8fOckCh4+ROrmEl6++vf6WDNWnlg34BXxd8aW
FfczI3ceqp9F4e3qzS4hwWg8fXfvJapKF5mENb1+YZy+dKkq2LHwhhpGaCaBfjm/u8jsy+biLSTk
mxROvHSLDYBtsfTutd/pPlWPLLc/Dt/fd1Keqz5+nntGEiHWFNy8i1iS7+Z79KtUOvuOyqiZouHU
tbEAkydy5VznmV8FuUDJhLcW7fSPMltwu4mcazFAiNQWtu/mOJy/X3SFyqYyOSt/ZV/fsHTraTj0
LV74f5d1mTfl7Cu4asp0+08Stw5tcKvypLRmqwb/eUGmUxtxv9WpAnMSu6oN/VIFnINvn5jJMSij
ukuRcUmAUXGC4MoAdoEKKa0doXe8wVdA3KrcArp9b7k4lQLQNdRZ68H/kGWykYw6cWvy8Aa/TPMZ
lsmnphs0ER1Sn8yv7PyiYvOcQDo30lVY13c8fbnNv1RKI2E+xAuEpw+1dwhq8D01XqpchTYAdTA3
wJlBAfX+tydk9rq5TkO9AOUSSuFNrJZ4Zf1oxr462e3VBicNtSzkunmhL8Q7DpAKtCu6EwufJMPs
TQwRSbCE0v71XuBPR7pEM8NvmXo/EdSNnwoE8m7/uNzPfH+V8J1oloUePWkI46vanuYLua84mPnV
VEiRHfSYLyCStc0ZLSJVHJUDRY+CFvewOidGdb2oioMQV1pn4VzrFnOg4BxIhD7kcpwvPCp+dFO+
fvFZFGw3E5dj6qQJOWptFAW11FjiZXrb/IDRLja3bY4lSWdVuKWsHjkLn9t9xsYffm4rM7wX4IQ0
iVCTRxPOwws2IgN9BdBKhwMR1Ny2Q4ES1vcBBuPvHK4/NFE+GTJBaIA9rO/eJKMSGKcdXCDfSm9o
oHxAaNwneBSuoLHn474CfrANF1aLsoWbD3p9n87jJhR/uMuCrukcql9wLmMdPzraj21B93q9y6cX
Yl2OSAsJ32f/4tiqDCozeC8eUPq5ijovYCar7JiweLS+jJVBWJFdUkUxkCtSsILX66qLlvhSQfe9
+B2MdX8ovIbcTdqovnriD62mMFfhWQJhyotT1wYZq+oii3rHeYZXnsPvvEPn3rlyWSh/MzHfkw4e
SYxd40iAltVx8sEl6Jm/I1yPYhCFANrMV1iIEDE5cKTZnoUAW3BESmvge/nN1wjNd8IcZrsDb0Pd
uM35bXQQC+i/5iJ1pZiD4C1ALAdEndgYUuRQc93xJ01sam9cOQofRcKbUTEH+DDcvd1Y1Ap0QUIe
RNNPrFyeBFF59kLtfktrT2gfbgJ8x2iAvZh9aWlQoYgjWGmLrkAff/ByznZYv7G68bhEPjfFxPOF
bYa2EFxqBSl9zZd4RSNSeUBjVq+F8GEho3JOttLcrQmGRmDOB8j6+EC37GH1KRn5xMJUznwaLL3s
2NewPbW59VhXPFqUEhmFN7mwbSy9LsDODrlqV/YkWuoCcdyqwT1gw53rjKMMgjYSWV9WuGIgDwHN
Z3bUXmHTjY/lnDVVv7XKS76TyYdHCGNQvQapdwntFbjF02qhc5DhGrtBbsjoKPjP5dFFH74ZAkDo
KlqpdAafZfaNrmvLamOP9EBYA0Nfz4ovftDyy02hNTxPRsLIf02786Od5TOMdEkX21mvfyYngVFP
Pkn0PPZFCkAumzANanlzn3tSzeBDGzBHQhCNq0/QUyA30ueSaoVJ6XyLs07WIqW3PBB6zlnKifkw
1sj+k1gD6aF0rLfev8ZOhOvJR2O0do1f5IOypCoQS+f+jVnoCpsEDVMQDbv7WAZg1lMG2NXwyTMz
+B4Y9O5SMsYMcHozV9NAPhrn8RTuycATZhjxf5cVrbWJBz30WYNlUW4ppGGurCRlfjYq1qOZqMAw
v+IGvgV0ToM/D59EzZ8qjDs1EmH0zcg4H40QXIZslm2IqNYDLNTQTCDMbHY6blhJHkqAx5IatQtz
J322P+B//ata4sHn6byPnsIFYY87p/8/clrQGUmefHe/NoR3vNVXkG9CRLeuEj2VCI0Z+XjSvftT
LpI1InPa9igA6a8cc3wJqHKoty1tNT0AIawY1QFOM/pshPGQRajZ+PKLqFgTpxa2O+HIJ/Gf5aSg
rg8Fo1nBK43LPCSPqyyfFr+/84YDFPNYfaNcISj2/qaSUOvzxq0N5ShDiJpnZU5m8y8gfzUHgBPe
LcW9PcwSnVxCg/Hpjtkq5jhJlO49Uk6zUbQBDsVKO964GwxvtMIE4fOFG+cNaJYhOLK0Cd9TkdvG
Qlbz+0RNGBINYGzEkxIGUEVP8dxqkWLTIKnemuoJMd5+nWqaSGVLEwHmfLZPrOsf8Wd9N+INdgUj
Y6RemRhwwn1MSsMJ8r1o9OtOkBzXod7WUOcwN9kYxcbq1lbKwftBEO/IhB7cOzOnSl6cztpjGnbn
bC8vGCKvlEY0LqqoE7reiSQ5omw+S44tvQzRFCJCGOkcYtq3zxv3CoCw2yfxXZmkhsxw82W/gxxC
qLLg61Yt9w8h9z03+F0LSFzqK3S3G6UZ7IlNRTp5Sg3si0qkvhR9mpgnWFNaxGsp6mYK823kOWo6
UlynRBb5gScxLsmbdhy312+hoac1tjZpEcrjonk/A83+J3dEFwwzuKD2X3g716KZVFK5cY6H8Cs4
mfwyNkQMkROyjXCdUriOTakTmMvVEx61XZfo0PBQTWijpL2DwXCJAHYZSwQ5kPUZQWIXmblyW3dl
TGV/qqkAl8hJaYxBgghJQNyiqKdIZ85lucKjGjTxuEtrG9xt57ovZfd8npQUkBaMIYnwrKPt6wa/
I8UhpiSiC8dzQIm6P30VQ+3XTtxM9CAFSUgYPa+WJKGnlTtzvsi3jOccd3TmiB8+2SQC8HJzYtQ6
K5BHzLvAaLWBs2xckepsA093sPOZ7Lbs8S16rQ4yyaSVZfxPNdTXwLKObStv+qsmwG4JRkAF0ToZ
TzK72ECO3IT7Qia5R+Het1vJzP3DFRMK81cy+RZh7+gfWkw/HnDAp33xUgIhMkdjy21HM4yi7YOS
ivsnzPdx4H72WzLBhiXTUFZNLVemQ1WJ7eLQazOcZ7RpM/m5FkfOyCyds160WuqI8h8vCXbPOHu4
YSWrYTP5Co8QAQACUVw3lpoG1Qjx7mYMobYFVFQBEEw2D/Ulrlw/KkE5mCFDCcoUlca6QX2FR6Fc
hUntjPUCooZzQCEbaYh5AeSQWqxLGi69Ytq1npt4xQpPKo/YpyrtPFVQjuwzeNrFNwUksj+9ow76
2ZB7BBA7s0vAS6DBkiJhZhAA/A0l2mrjgMD934r7vaKNu33U99tUscnriP4LnyYYvW4XHphDryqC
L8gMN5sFJjLHOuSaVavJ7WQFTsdJKE9mmug931qTUP4rVD7BC0Ci12AdZAngYeH30G9DWj0BZEZc
IgO4ZxbR+VVMUfjUJquiALH/gFJxX3C5aiv5Cd5skpW6astYYwDK8xYBohYxepDCxijZFK5Zn9jq
7Oo01WS2WrKL/SrJWibVJ6ue7+D3wLneFCL5mA+beTwMBFur956t6jLjO8NphFnxlsLE5yTrmqjr
GgrkdyL0UQ9VKcAPeNCkeXoH7icHcJcVWAX2hgZ/28/EpmenCvR7SwtHXs8uvVG+fmaPqG3hNOy8
8q5/o2fYzVedKTL5AQNSfEleB/E906HSkZoX7T3+fQ9g+w2gbDyB/GM0mXRMZOYrvHYcOF/Crpo+
3cqbh1wJEmwH0MNftjfXg6j6vFiRRMnPrG7ZDxY+KcELajIyXM2iEWi/BisZOmGv7JvwK6//16Xt
u3ZGAnWI8L7zdfkgxFsBmTJ9TQ81QOVlrgycEmcuSQPDy+oNEqMz1o5oM2gW6PuRTeSLLSZtbQJX
QdUuJpuVtrxFmtUXBUk8V9FOwAigoDCcb3pa/DozMj72R6+fz3dUM++sNb6AmymkSG8nQYVHNwTC
hMf+5+eJ23eDGMmXDYfBX6no4WFtHHcQjyu2oWEgLI4lT8CstIUdv1mZvcBhoT1Jt+ownXHwbNCU
wI9+ddTGHY49Rbdv2xxQg72cs2PoQ3hCxsp1scqNgyvCtq77YorE2dNPw6OdFgj2uS8rMvvZgF4v
poIa7hveIL8A8u0m2pT1T5DcgX5aQreIJV9GmfjfIyc/CaIfzzCld8HONDk+MGeHBs5hV1e/HmxK
TD2nHyyRo878DOVzveZjikAB8eBfdCN5e0FMRcnij3Q43Zyb40rTNbmN2E/M86QP4JxGlaMxJTv2
qtSAI3pLr3km9f3xGIcnfaySVB0n+IPVmTIixR1peJuy9f8yOG9amNYRWOVRzTTJHaDnlvPhFNtv
sF0gCwI4dxj4thdMr3emRoaqnCl0tDcAkevEWeG937Q5qTW+2/vSWyhf2KawSsqOkTi4nA81FE7o
JtJXSfV7xz/YWcpS2AisIjtrsf9ENQHpWseIVyomXZ4nK2Ro/009eamQvXIDqeWIcyT949EgKCpc
CuUdxjVEjnM4XmEtumPofLwm3WklFqfQV02BWT2ph6/rRWACmbos/ukFI6xV8GJfRcd7EUuX+cI7
5J9vIt3B/0mQJ359D/xrhuuwnhPgx3sB+QfwSnDECWKuYvD67Q2JGh8KSt6uXrliB7YXkaa2ShXS
06KnGBNOAy6kDWU1EhwAVIb1Of+cDyNFXJrAlaXLnQjdm9PKm+C2WfopkHoPDwEI3+JTu3IQfRoZ
cFGIuxzH4/7GAeChfZHVkrXLTpWQfCLZV9sN5a2ECQoVepzgOMIOXaF4U1+whfiF3/BnJIay0tFD
c3s6BATPBpjebt7ltFzqDjk2hhcDE0iwnf94UsftL0JimZ/WytWzBH82psoMMOR5DcR6e9NUNQZw
EUzbHr5l1Ndl7ZkLuhLIaI+PuFM97CqUPveBTY4gTVpOZEbN6ir04SyjZif4pmttB4zk/GgwCCvk
vOhPMpJv8/VkS0Ql3/EnwbgbgpzJzg0fMWf87FaR0tk1qrxhk0y4PBbaa46TZLbOTozXmmr5W2Ae
JChSHmc/d3W/Xs1WnykMgLxjwfjoY+Rza8Xsa96Ftk+3nq+Yf+rJNwpaZqI+dbmaFYEi09Q6hL8z
ET87CyogMS5jcrsJXeRlYTErQxGkge0VM73H8PVteRcZ2Opd48JFLoQXk3M/lXgPPR+RE6SRfd5Q
nk1+UADarDjoHsW1xmbE3HgXMgTgY3qXwGr90MxqkWEwi8agYNYWJ1BFd7+UlIs5iCIWbBx5T2yp
tF1hbP6aNBg/p+6QIXD7Wvoexr7gZ6x/riEbv6ddsbgrlE7ql6AgV999usz02flpAL687Rq/gEj5
C1p6wnygmW1ejuQb7o/LIx0lbGbbP2PML77jEnekzAfQawF7gZuAJG7VroBaFYrl0ZJ3T1ITJRVW
QNIAVR7aIaEBPrnc3lXrePMSO5fkpEfuu/5sfsfQIVOvLfspZZos6O8Z9jO/r3PKQOVK++Xbd0VV
6eHsseTa2hVMj8HA5Acoux2BtjGi05rDt67nye2tHcL80bpum5+L3uXJ2LAnUQL+X7xK7aQfLOtJ
vfLPMxcLNmlM0/vhIC17Vn0SECBqx1M+U9OcBsD32iKhmw26Sxnwz8rwXRO9QMLxEbNmVrbBYBw6
p+QDujZwbQ+3rUwAHhHRw2KdrK0C/081ZwO+F9/e7bzMVkjtDsmjP/QnjATSLgmku1g1ohI+o00R
su+VZMmQqePJP5wxx1hDfMcoMt3hS5VIBtEG5PMz3WxA0kwC9Ei3IHEgo3fcKZMJn7M4QH2ydQbr
g7NdSRWcqP6RM/XqdgRLAFBTBp3DQs2QyPHDYyy0oqFrs/SpPeeWP/JOzPqIJ5Znp8KqBu9dFRY8
gopANB1zjx+hSNt0muu0rW9T5kuKsHiTIw5OCl0sokde8EWA0H8gVaynzBlQInXj+Hpb+bLnG0rm
aJbd5o4bE0nv6ab8GLnOPKpgjB/IYJLbcYIoG5OsWuA2AB6MLdihvelMAZOKgpjHyq66bJczZuyT
b4sQaWHuq1p+aYTf8axZu81IBKA58jUsvVo7okVIkaAH36I5HN5WGwvA+2VDYWO4u8Ikh7bFLtic
ttfkqwfzi+pvkmnQ01bdMv11McMPr4wECRdSwta8Z28fhlqWBqqMk0Q7rj0xS81o2bBXlF40Yflk
BQsvHbCzlUfoNyPVwHpBxkDwIoii6dGBATet4JDjL8hhN4k4Yl6p6cvX2urj/BgNuMxWY6lNinna
1m/BcvZ9Y7nXgoomncA+CO//ouAk2a6Ljd6XEaHItX5FydsEMQU+ToLbYl48BgNZ/zfBy77RIEKP
kigLkTDvl1CwmZ+wt1ozr7x0Jn9e4OJr15NAdExtVDX2YLiADv0tv4e2vmQdC+Q+niw7uIyOr3f1
lgKYZRS/vOvYPbw0+divv3YEaQFhL+KlCu5q5acHeOeCy7qOs1z4JirRd8UcNgtiQzjm/eDsKU5L
pIDHjkOsrQeOgb95DpVxREyhK4n68HHgjGsioh4V6T5ez0ecUpHVGsGQS736eFOeoGhvRbEXks79
nhg0XAFN9Kgro8qU8oifjOp2TizvGSkqDbw4vfv/BpB5U9WcslF2NKLTuV8yNLXuvfjgiAkivQ1v
7PGtV25VvviXc+3qufxRZSUGtJ9Ks+q5PL9+BZcvlvSAN2NLvrspLUT66iwBAQTq3mkMZsDogG0S
Zam5eio3qZWaML7NZ/EWeAa6gFJd58SPZBLODazeq21fnV1qhPXo7y6eg5cwXeWrioOAvtJ5/OCi
xDhDBxlxA5SVYh8DXVvzHxj+krM9O5ygFpmty56UdwhbZXQBMNbr4OayGaJZ4LhldKciK6UNwhTc
1isth7RhDCMjZ1aSLBmKwFqzBn3cT9VP2BC9FjQP36nfrqeDN6o/Nvk6fuB5sXiKERl7DP6CWstz
eCRNPV8wyN25HpGB63leTcLMxzVYPnAVo42WwUPtK2lc/y7tckgd7t03krtAuvLFLBEcm0Ov87m5
7Nuaf/myh/7LP50q4QHLS1pTl3NPj7J9+KhartXr0lKtG34o9w4aIWtn//o+Yt7XyLy7wh90i2Yf
WYPikWu4LczRc3WZblgkMgBWJYalkMGI+DykFhc3cUA8SlFrTm7TWU0GnlrgWGN5PQFUG7hdsl9a
sE33+lkrnFUo4uykgjfG/UFLKqxf9pulR5ae9dIpkPSSgmw9ZCXpuKGrbaLhcN754kPHdo6iJIxC
6YduMm/8ZOb4Sdi6nwso3DKpvQZQMCtle29v0nfWm9N4kdyZKIzVU9HXYisv+KPOMLZ++Ej3+QQr
7XsR79l+BfyLjC4dzqGunU/2EmW3P7ggXkGd5JdWbMKuO1U227VKTxz7dK5ZDjZDkI7KtYAxr2pa
FOCQ206WB+hRV6m31/GWg9Jf+76CcVfGhQqTUwO0DMo/7orlZIY5UVrppRAQ+MB2HQBdeD4/JO/g
r/vRL6j4raMMtIq+2D5GnT3+OBr9PX5Wo6hMUqW7uQ7SXJW22X6nf+WzwFK7RyFnLV7/9mjxe+oF
CBjXaN8dkE3X4WcG7Qdn+OLWP3LQWHJ3KPUC5NeA4bCwIuPhbIVdU1CEbcnjYgvkK2p1aesqeHqi
nF17/6Ite6e0b9s7L9nftHTACN5hxsEgAaVUrYIV+tJYRnFPepV2f46G1OWj5SGNd0d+fCK5a89b
U8Jmq8UyFCUwXWE7yck+KLftlAn2jVFS5o1FU062qBLkMz33/iQpZrrgaRWEPOIl4EiVV/JPQFD7
q3/Xka+/x900eqUV0BRqOoC8cpKewg5IjZCXyAxXxrj65SwmCov8rf2wwokW/6+KC8MG1H2/Dwfh
KrUKjDYvGa1LSehTA6lsaQb6m+rMm/dalh2U0oMknriy20TyHEvAb+fE8iiDCs4sYBImGBldq+9e
M3RCE7gzZyUU1ARGPSWa0KDY66zLH6ERMbPhWAtaa+XYa6uNS0+Il+FnPXYvebaEZW2Z+QZD3M2n
dpU53aP7jPhff8UxQPd32AMzA8KOMLXX+DXHXkUH9alsWRoGL3zEh2XohI4YKzV0EONuUg9vOI/f
jKtbt0JOSL1ie/x3wxd6CPxUCyVHg3jERfeImEttuHoSjKksD4nyrlo56MG3mF97IfVGFr4f0JoR
SgsL5GDqxJSweZ6676FP+9ZhHjXvhWwNTLpNzQxcgthJRn3NkdrXOne1P/d42S9t2YQ7A6MxMfK1
D6n3XTZ2k/2eGvwbsz7XRGi89wXl1OV5OzJiKLClpy+ijcC0cFHTYgx8vLyrNQ91UlhDldfkoct1
+ScSY0op7RSSEPSr1J8guNKYFXOeAWtcJ5BX9a3hkX4pMWQd9NwqsHzLhaDhbLNX/QZ3+cXTmWZq
l5TXUUjzsADUshvrTOqt2KKdp6Vph7v0nHKi8KlbXnXltvt4ZIWk18jx647hy3DZ38umIIK880Mx
bkJ7TUyNXv/1rmwE1LLqCGmTIa/UtbXaGEo5bcT9xqOxatk6YaKCCd2B3uAw64HrxqEERS8bPWxQ
UJBsRjxppGmeY/9RVPKANkbe1yKv0zctDVGo9HyZuBwgxaIVv1xrUvgAL4kgDAjhJhsKbtd4Sjp8
K4a1ft/qY+gvpDAtcGHQw+nrTBkPOnF22m6rtQPhiq8e/V/QEAyRbbn+X5xAuQC5LAY07rjms8zN
ZZ9BJW1r06VAt+Y/4iPH4YZtrPclYow2s9RfBfZa5bYUg/xNISajLDLbKGdYqeFwvKmp3HLCEIob
H55cWaBnpdoHXYeupUjiypBRgmXlVAla6kfgA96Y08JRYF12s2Scptb8rYzTWJ6ZKiPjG3ZOaHxK
kIIlfUDrkCh4Qc6lFhgWBIifenbD3xHvNwBAnhshtSjfuUzj7TqOZsgDkefvKHJ1/PfKbYDBaYKV
ew4S84HHoASBNN5izxTFH+ZPLwIPBwNZf3+C+40A1zKtdhc3S4asjaGrqrJhnutBnNLnJCtvwd51
ZrRhW35X8hhKN5jZhE3BnVqy0MKaiUmTSvh8D1RNJ4e+0e51VOyZj/GgwJjYqhn6fsg1KROEaKCQ
RiRLc5dcHr3fxq1kRAkpVMN7kn+m23fVFvF4utiO9/rk1+C0n7WZ5tZKT62AsRW6uzGMqBUx5Dpm
knosWJQt61YsVehggh8AmpOiz2K0lCRzx7eKR16M97Ta+Ud+CcvcWxw71MxL4iPRw91yTZgLUrBt
u9rI2+C4WW1qaSiwm0ITiQsvxh1Zw/V/M0ST65Pf98Um93K4HRTt7kKmqFIqcDbDdVAbSVqjGsa3
Ut27T87WbdHiiwq8xrNtiYEVkOJW4tnKawrV21moeuYScIYxitSytRPWkT85MQjL8ZnIMC4roGot
ZAn/DRIrLYHXFyIFWlY6U+KkppCyIqEqVDPCpOan1RO7U7wdQvaxHz2zVOYLfERL7zv2OSngxWny
h0PaN6Pg3QJNYG4oGe1vK1DTP2rq+rbiLTgWAgdW1FRd+f8leI8Q/9YH7QTanlCfGoQMHCMZm9+Y
mFADbNfNcc0NXoirZ1+WVPFk+hyJmgpWNUsB+sifI8F5zDuwiuD3O0cWSSJcfLMpdfSpOKf9YeAn
5o6KqgS7HvWVb3l1XVs6YdOScEfQU6W35QCVTEm0Iz/7L7gRrMcNmgXx+CsXkUKBj2jLIP0cc1AW
2JnijAjKb/cRUBMI1qZXK4nA7oM9E/dRdpOca0Ubaq/bqDVfRatU5BmVZxqyk4Afi+hIpolG6x8Y
nfcbj5HsJUF4stM4nYfTgsAfc7XwqXApkx65tEygaoqdYykmN/GI4eqQPOm3pYgLzZ+q1zLQZVxy
aLY1yCaOS1XsEc3TyY8Bsh53nGm40uZ/canO/msuoXc2oqpfsOhK2R0AmQ+TK3zJzZeC+Z8ErgRi
HYYH8+xIT2E7CoTkJN7q2UQHKm4vg6UcTZse2QVx1XHV9ghQELRJwj/abwsxq35zNRWYsEQWjA5H
YYfLDEYjOrTdzd6fq8D+tyqZTabL9ifFalHOR7kfPEWFsp81DpZVoKjNmeyfnG0659ed7oHJ3Qev
t+FdYZbPFOLkEFGvBnzg3+3xzDXxdGCXIF+6CBGWlF1s6rzOjsPw2OpgmrmNgkfkSC9eXXFjZ1yo
uI12t0EtN2CVod47yXFcrD57tMF+UbjT1CqEt1d4ugxo/4BxmPdtOVkUfWKRGvnamuwT14fdWlSS
dKiUm97F1R68xcccxER8Hoy4kObD+RcfKKhnHzPWwpzsWwgN5Q7WN+c84lF0hXZ45N0dhHUEqfBX
/niP5kM0zy9pYb5mp+nC2IJN3xzQY/+/cY6GK8yfLupiGUjrkifgJqrmMnQmnaf/OYiZojvSX2DB
Y/kjSCaG8HjHddaLZBaeoMI7CR7+tQTGmiVnxzuIJvJv3mFN1cFWXYmj+6ikINafldoms0Q2QBSW
ICeAMWlUrvh2EaFLDc1FIxJhludzcyaiCCHCcU3FVY856mCjc23v7ObvTpe+gDQRf2lNpaaxgpdy
Fa/TPYCFIEyt9oq6qBW7lCC4LVRQmEut2IS6D5Oxrk/8ZNc7L+uD3Pbldwvhd8ie8iAb3kuB200T
L5yPjvmfvemzUpU7d2QsWoCoC2rZ0hU6E78Aod3tkdSxR8oLSpNk8Jb3lKFVFVMjHH3Gw+UjOb0l
1XF99vO9ce74stkzU7UjkcFW9mOp7MXs+loYhM6M1LI9OkkP4fwNVSF0i7OkSK7CbzvEWAmlpYM1
KX9+0MHfswwC2JOUIEcLquohJRGMLon/ejObjTW+nZfwl3QkOcSqc2eZoaISIbE75z4KsYX5OBEz
truR69kpGAhXsOGFcXSx7a+/bOb3l9KLEqa41C2LEvZHXVZ8xHMYvPklr/pAMJvhFkGQAlzQD2Bt
Dh9HILeoSoYhpPEiJvBqmViPDhcF0+yz1cM1Dkbup1CixvbtuDy3pe2zUKaEUbZ2C+871JxamljL
nUQOvN2mCMDwY6NdSPGj5uT4bjJDBAfgos6kiwKVspWwI70dWl2C1NfjiLDsehxuqjoX3mABdg+o
Cv6mCoUNAywN+0xayurmnNYub3QhF9C72in7zeuzDPzdTuDPsK3GW9SwXRSCXRB/7Kc2K23VpzMg
2M0jejVqBw8bwgRPGoQA3GJWMUpoSSED7sbmTR46XU4hJW6zt/eov7v173q6X2rWFVVjZWrot2PB
bLT/WAkuwdLbfL6XriOh45uyZyu4fbnUaV0uCC09FjeafC2R6Hu097WTEx4fdrT1k4xY68MVxX1n
NPMfTyh+jfbF2iyQOmrRlHC95jpX9fStN0lCiIEUTeQ8gQ5J6nFHFqijsjm8mpz1rR1imHh/4sco
wqXQwVySABVGH0UVjpaZeER2FV6yTzrgXIUILbFpwp0rjSX1Z4uDpbI7OTIpmS24oCfCcLRvB/Qa
+GbIucPS68zgpVubTmUrhDsJYc0ZaU5S7XJdW22ymMUlDfc3o2Q9NObCIjFeOJHwXU9n4FtqGeBv
HHRvXoKf2Vz6uAk7w+Qh2vEr+1+bVZwsMs27aVIO/eOIBVceoY34SAO4ROchm7GX8CYzYKkULWZn
n57f1xQxPfpcVFbuLxJjNQ8JrL9mVxcRfS7nnjjqIrrA8JaFjech61JwSLpHSb26kG9+ebkLY9+g
+6PjMbKwjki2OfCINuU0KGCTx/42aBELYUYRGd6YvEG33rpPZ5C3mcGlABEXNcz++PnzYo+VVv6p
cvmTDpn9y71a8AVp4a0GfqsPRYwO1d3NTl+jKMWqJPsHyMq9X8Gssqsxr1Weypv3UjsfcQO41sON
yjF2qfhpgVyenxRdO2cEB/M+ZBOs0IPutoxfZoyiVl1AAFGelcvk8ThGv8C5/qftssOtyukesLJJ
H+731aZzOiz04eVRKJsoflRkvWGcYFgdE1Ks6SNNT7A918PUV+rSFTqFz2rVI1fJGcAyp77AUq0V
YU9JHPi3EmOhUpFEpfwMJA9YsBZ71dw+rC1bw0POvd+6LkR+tKOn46T/iVX5EnWxR07TMqbG/USi
gy4Wo8Y6WoEFdBe75UF4fp7h6MEVDHKCEhI2WL9E/29IIAoTS4oI7AqY7yI8cO8G0lCWGkesybkj
DmCKaN2WUS8k2uMiucZpNNxLeu3a/Y6BqMVhQ2w5s9ObnAj81WJFxb+Z/A1Esf5MtrlFCTdREuQP
FR61wxUGEIvsSopf03iMk3FQCunFRYpNvgV7PDZMruTPvYvwKhwVr0SeZyAYhtebknxFVKFzBQU+
Zsa83oX4ljyfG6gbbLOPjGcwc1aYpeYyBzEULpiE9063WPU2RbPl+O7STFrpxI24kz/95wBO38rY
UVuvAKFwEp0cWpFyLgU6AR1UATzOnf/14/nEZ9wZlKG7EgGyEzX+7fY9WC0lRfVtRMvOr0V83IBB
hBj/SplzEHmrZC2LjtrbhXLqkWFtUyXqq6kupx0xE0YoR6LfeLrcw0NovGQRdSq/YmFFdNWGbcg4
psM1DKYT2UDDXTwzNtnT7U7heAyPLYLRhWL0gML9LNMpnGhdUAgTFI50VRH46T5FGGAaUf/EXRuG
MvsiT2eXGTKfjxlWCjHsAgmTrGkmzdXtvGFTWEcX95gEIkTOvy7tv4RKd8+bLmIwNDlNtR3+L21r
nDQ8/Oev7iyq7XehZkp72FtmUgFOhAGdyLLZLjpfboOc0QvVoEvMzJmaRCcWckuMEl8qbFLlMkCP
/jnbTDmwN9GFFnf1TH13Z4UhHzZirpTIYWfzxRnWvWVCirK5+Me+IRwg1kRWQywJXhvHMRb5tp15
5ojhvYuetCLSQ1+IJjC/CxDhx7yi5dlirWEOv/xgf2gHYVXodJxJgSxm/ZvIivD9bM7LqHZjImOX
C/7iXyNhkaSfEo8tk0yIG9Odd8zqjwnka1SM8u2YJY7WKsDktl2YzDVb5Nlo57qpGS06zlvbPqgD
K4fEK311OFsmHbjiB4r5XRczn9vmmIaf9/3+x8QigAWKn7EFu6vmHZt+uvFPH08uDE2oMLjRHCR4
mP9o+8D3iIoMBHbLc0f5tSkyu1GQ4A0yuujDKrk+OI5gJYpOyzk1tMyxSza+UQZh//vjCjZgGzjW
xBfg0xwFs1crcnPa6+epQtOFfTy0tknPs9vBeETT1A2FHn7j869KuvbEOsOqD+lteGTrsVXZ/cM6
EZGQluFv0nUWHCIBiyAjCcTWHXCXSwrfw3AyNex1hpiOostDgrAomf3bkQ6bke0l+Z/RQemd0CPe
Nbp91APN3RB8D7Y315dVa8/OILlmU205p7tFmrr0DYhQWgfxNzkxn1avkydSzwEbdprHHALY4QW4
z4L4jwku317FnA7roZ+F2soR1OyImD0h58DNigG0M5lvqCXXxkPi0u/dlYNNAjh/a2lOFW3SHOr9
eg2qekFaZEthr3XEvHKalDC0LYVUoTdXxSaLh4vd5zu2+ievSsmrp1VXZrKUlOvt6JXcKKiUBMmW
J3crk6X8atevJmSmZs2GjKpuyP9DmO5lbNXp4Xz1nYXQl382/t9TeRLYx4iVPvUYMJdKm8uNbAo4
1nq9onu9Qr2/648ySwznonn7JQ+SQvX79Txu0regr4xVvLpZr0XXlYWCnqAQrmJKBaijoDoqiaXk
CUC92GrfP5071Jnn0PPcsWSKdgzXLKbNlDAjQVmAZ8PqnToEz0NXy4jLjpexQHJg2CZoQ3yz/I7W
eGZYvfrPhiBhZq2xUldwYd6qiF++729MfeDlswvscomliHs/l2jUEMLN7dpHEvjaNsbk4PRb4Xfh
rp4iatO+/csdI4BkAkEwQdQaWCakF38K1SoCBOFfhK4+qEVVJg20NYCo2VTzXoBMPeBe7xGMso2B
mx5CQn1MMRVOkxB4finQtj0hSlgz9M0qPKPmypyVDpnuK29f+sdZwgDFiWqrjg/aR0iNSmbTygtf
sPZol2J/BDZWzkGABihd2ppE4P5h4BRxRfPs3OojpZ0lmJe2T5EbcuZay7ksuHXClCF4amSXTPJz
zf845uvXNRAm1ieJSM1DVtAuWgzzJRdnBQAznaqB4wINY3JwGvYkg4yMtq2CtLz6+H6qKKR+N0G8
8MFWDPpVlU3lrt1bHa1pK0ZIzbh2Mybt8aKVVL/Zs/Y/wUZ9FCWBI60ZjelglZyl6h0edLVzyEwN
b4z+6nrSxrwQoLzLF2dalWtAtm9MG6YoVAJceVeddXnZang2cXsBTqy/yP4i0ghyCdbZxNylWnDm
rjNjzFPZt+pxL7AFJOAE7W4HY4wGPyckp99d2rAKh30pY8xrYzc3QG7IGTzK3Bu2eJaQip2mQsuZ
lguD07rn1oItE8FeyV+WFhIhoTYw4f6djM3XlQ501xC+xXY8+hkUZ4UbLyTA0Jrdtev/rhRso4TS
O6W9p/fnZKDWrsX/rGkzBW10pJCBM1jeyBs8hPhaIPwhkPM455xDAJPqvts2l1VDdTKvv9c1S84G
aIRX8NF+GJju4M/ohdOEJERXs301kN7D2v7IjcxtQ2xkKP5jgH22uqj4hbbx6Y7dqQz9ILQA5bXY
sCjcYhK85MRFD9XTHxqWLaUkjaW9zn0U++DxXhvXZ4gKZ0e+1jX0JGS8BHFmtlQjpyJ3UGgW/78E
zCJZw59SbioHnfwCACOKp0mU3jTRD7o+gDYEQFKRoe37VSxaNUlF3cgoXi7Z8hGhO/1+9Um1URom
B3BXQAGZRAbRi+BtiEqqCmVZfK5Mq++p2fNZVxB/g1Z+xZRfelHXSPYV0URQZTutYR8JSf1e+SD8
y/ofFEeOS2m4y4WloBh8QbnSerxsAKp86xUyiPf1d9hgzsQbAnV14hs8CB0vsHEKPAcFE9kzuUhT
k2iC3GQZFYddJhSd6u1ydkRnUjGVea0UHVKjv9DTS4ztU1XFKpkdeD9Cnq51/9ZFGYJvLUKkxF93
neJnyuXyTjqUg8410h3aO5NOy8E1IBV2Pf/stkM5UHI+Fg7QeBiiauwac6pjKUIWN6WuKb9vrkZI
uy9vi7uGtQwt0MM8D+g7GZ91z84FRfVeZlfGNkJqB3WRczb0p80hxo03A2e7lYcH5NRDAjapG2bw
EAJN/MzYnHyKhV7di8XOCqJ1PJCPe8DIwPD11sczrkIImDPW/uW7MAuYAoV2hEvT1BWTwUqMipLK
S2wIUI3pBAEmmbEAXnDsgFbPZvKr625Xk+5eTa2hZAimEri6jUboz+GHd5ToXp/cxPYSXnWr1+a+
9sRFVfjoRWFi7i3qgjCxiUJBQZKUR3ItWHynZLsV6Sbu4A1puR6XaWnUclC/3a+jmSa2v9PyF4BV
PQoWuulW8dB0jvy2Rb7TYaL4VsaD8pZYUYdICxqOEBR4ae2lfhtwYqdfAWL2yzXWF01FREBrXxkc
HRk56W3zBfcjI9V3p16zOuxvr/LpGkt7vxXt8X97ctYgFFZCPE6Qmf2NRVXzJ8TGao4MmKXO7Y09
E7cw7FF6uaUI8HiFG/5DOsYsSpaCn9iC8hzwIA+2sv6EnU2tRc+EN10QEmSSP5lvq80BjCVM1iDJ
uTyb7u0vUGnFk+mACDTjLcTagyBgdhboy3mitvlYZdyrnouaVxCDIN0+QMQiyP6LoJaoT/wO68xs
f+svXOvcpj4/+7K6xesMwdZTC/0tJoTczdYqzTWyU2OGxWAKdXFwu9jF+2DqhRQxU6da8in3c5/i
A84Atu2L38aHIhLLF3vymrSj7VGZWB6p37gN91bPUoYWAPOz/Gbxfvnh7+GI1105HG5RA97xYMYC
USmtN82xsRgFXsfcvOFSsEYUbbaei5hHmHWBWSE52SVTYMWS8Et1C/nJMxaCftmzKBhd4CX/15h5
vQlPSL1ZMsacEAAco/tjurRHQ1czpaNzDhaxmwZqUWOQvWVOF1pFA94Wu/k8itOjI5HtUPdm3F09
aQRG9HrSX6LfPBSyww6EcYcgWwlGcVrnNG8B26snfXTi1wq3YgNOhAqOQtGPZ3nBeDIyl2mERky8
ELLfWBd4jIaNuoR6mYEmYphlq2Q/OHkhjNSCcuHdq/23SzDCxlGp73mPl8Lx12b+2xnYGCfgCVx/
OtvcoXHxwIdUJwOEzGYvuKCmjjzBMu5t3a5F6H2OMi3PF8UxJiuowqsi7q2mQvVYflirFgldC3RD
WMMdGEEix8aLglMpVUv1lEkiSHG4uq+2CX2JZ/Yrq6rV+lNkNAO7W99Mg1269z6X/5MgLZTaSy3T
0mUIGLr8AqCt3W5ty/5mGms9UpORZVg5EOkfd08iJdt8Mb9MBzH/qBESG5BsSVjLGV481h6U9ZTW
LxLpGITfq7/s5mtny/mt/iapJERZqUn3QmAiPk2VnbbaqumGSUY64qxfeFKuu5Bslx27OgoLgLsH
JVpVxiBS4UG8AAcImZvqlmy+hn4APvaw4BUhkmcxYA8rDYgII8Gt218yp3N1Tos1DYXAhxQ81vIk
9nhaaQEZzwUbVmfY+fddQqV5xnsyF60UG2bqZJ02znlPpVfv/MohY+WaoQbnLd4gbKQF5U4oQLhN
pByBhzpHEdorN6CoyqsKYtA/pkfvxW+1M8QNPD+kQ/lAJGlXqXuscqRGXIMnGoAJ6QBK9KiZSAZ6
hu3aGPcEy1LJYjpRDvuQ26KhVwaT81uzKY0VzGMivzLgqIE8msZQ004tAa0pe8NJcbUSJpPXr5Zp
aa1KnRLm4BXtVcVbxS06beh19T/gGj2J1XAM97URc44A/creRrw0dTseTl14Wfj/O47hlVz4L6ka
cV3CbcoOgKPoSvTyM9gGfLZ4XZ202MMyTlDyqW6wxc3aF1mCh8NJ4U3XZ6Oq/Aa+P3MyljKTZH3U
pAOK8agDcIgHE4lU0uOjqgDYHo6JHM+sAXB3g9lhp8klUd1Zj3ChiQcumdQz1JzbwtHHpL+qbm8F
XI2RMumOGefqcCie0v7y+MmKQISAG0bMtvGJEw+0inp9hsoMoCJcmvd4Bt4L0RGs+/aLbrPP06on
yt6oq3BasGcG/wB7xyadqQcjhRwwHqujBlqLpahLV57V3b1K2LA3kwGVQoBQ/1wNmbW4qOSvXGYy
z4wN/6Qtgoc98JXg7k91gHHb9FSDiR41vK716jo21tGIKRcfFXfaqQL8QKWzmGq1khxzvas5JT73
h1OLsYqaUFLrYh6DjhboPKtEBYsPVles5Liyi+UstwqayzzT0GtrMOlnhyDiCUeZWvR+gaES5yJq
zeKx6tjwtzteECWZUkIl5djcM+Tryh4OeQuHr/LtJhMr0EqNZpXF+lbggSdLMDZ0sJmxwyFXElHO
xe9PhXzlukHkTpue1dRN2f8o/OXAtN0McOZz/klzDuL90/vYGLFrmhgKGFXXUpLy8D4/V1hKdqa9
zI6yGWitcfDdTfRwZ+B4cpVY/v14wCrCk5L24S5cCTNBA/3Yot0l97eG9d4eWHvNiBxmaKEG3NDn
1Wbg44abrK7JaLNUHlm8CT9yYObttwYVKkr/YRTf7bTnP4TJ5IjUa+MdrEZOpZmSMHgjn4mUOv97
yqBhty3ELx+3xQ/HR+lgRWW46FYhNzSiwuFONALAIADTv4a6O82hLwMzT6H6M94jk8DIt25ixv/o
rvFYPOweK5OYaIYprFp0siiwTnBuQebG1lYYNf8naD+srhTeeAuvWrba41o9ln90SDGncgYlyaVs
xOrYMOvA0415JEun2hOcylqdgFfxw5jpJQvnRlmGTfVm9jvZJKj5awXuvmefifUjlnO20+C0FExK
sTTE3X9VdLPnO+wfqKHbiwJ+QZqV249AWwG5xyWvwPfZhCk41odjNsxND4Z+LB2ZAI0z2hbXKl49
sDAwoZ5A2Q4IoW6KfDALcmBZSt27wK0X+wNlrc+iGxXMRCLdgT2Aj4ZTEM6agVqdL0D2r9xQkco0
NWnWvSPr4s/DxQV35eR/lE4CGmZ8kIyoCF+bwnOOzUPB0LqYJzNShh7X3Mcleyhcyd5iCTy4tCxA
vLvkERwOM0e6waEoRtLNpaFG+muQ2w30QUFjARrSFAA1hK4OB60CZfFVYhWPTzM13zPu/7eS9b74
2IosS8ELEu/6u1Cd2A4cRcfnV0zUoi876PLQmYSkOWXoxxSX7bqWzX7vA5yaBkPUOx5nichRHMbR
8Kjc+Z9VbIqbnd+B2CpNyYyA5gpBCeobpvyJGjYt98Iwdo/XMtMEakKruHLCPG+fn//RUOu5pfZ1
PYt8BW6vSNBM3+nVagUbdkJo9+wv+uXuT5UQ1lmKOf5x+hrE5fxpiBFvdRIWtaNBeDOMkW/80iwC
Oojv4ctNm5dH8lFWURDk44nocQtteNMfD0GuUe/lhNhqOER7WJgcPdHJkpGt+vM9iQh5D9GlA5h9
LCQpK181Fr82EvOebQLYYuubGoYQgTAUxQQPR4rmWVA5JCdQAZyAXnMdzJCXGuWtbBPoggMI0S+2
ZRMJAp5DtpFEnSdFA8I2jQgf9Ig4Y7m5GSCBbqHinKmYFsfLdZWIG25qsRKwtehlgdlEvXimBrlT
8mphNGNCosARiZ5Ub5Ee39B5/5HmXDr7oCoSdYtgrThqn39NuKQQRYMuAowlO+rTv8e+U5mqsntC
E4urTP2MglJ1sex7f0MNnpCz6enBsIu+sWkPinAmZbzgbSRza4wq5ss1UvZbzB2mvAOwMPYXjbt1
3Bi68G/tQd5UH/HvOdkq5rnYPS7VODC6xMdG6cpBAt8Q6Z3F5y74cNHXR86hRSaWHI1avbvK9JgB
+PJxuQTsTuQJujfk7ivAiGnJNFy/N7FHbDv071Ei8kGQMS38wHIJ8VmwI6Tbaa2/GE2hkJYVJchI
JVxn2E5G2czaLJcmTcCRm2AKJkzXSejQdRhHP1t1Gdyk+81F3+4hHmgWYZ9kDXuE/2tB8ZcRzjUj
vbx4Jrk9LW0s7+aBQAfNB6+DWWyfZNKrMG2vSuKssTilxt+NUO9CGgwBmsY240eWvRFfX3NzFq7I
bzvqZyKneyDpXjlzkXABXxU9MpNGIaDmBcIKSyD62CPX/EytY+w5g/c0lM+0t2u7ff3YZBp+xECv
ziX2GgMwgtV7gCy5tyZEIQdlRNNBVzTNL7nH3q6e3H+LIvqQYeHXdcFIAiif9DA/t3tuJ1OTaIr/
Xh8bNo05TZFtXpJDpp1C3aD3NGbxpm8otI+MK0BA26hWbW2yNI0EMTLNgrDDVtKEomNTxK9wk5Gu
+utnizjzuznSHO8WFDxy0vX2XvPFgIt/o91AGP2GhZs9Qq9fzOZgy1GvBHt5zKh04fGnvwb44oUq
0KGUSClOD/R2llnr2OxDFVgHccIBRgM3OIWebY1oS+D3ZNWmH8KPASDXzvB3D/O/STaKz2kH8LQ0
qrcg597/LjtQN5B4Gr3U3ZaMo9NicHDkq9AzD5vZgeGdGxo83lokT4uEvESIj3ssmhI8PCyhqo5t
OHeqEVWSNE/xnfOjkikE4xqyD+DLj80ZT5XFX2CwttKVHa5MFirJj0rEQLYJe2z92b6frVaIsKzI
Y5AtImo8jArXyKvZKFWUh2WznPeWjj2aAbndwwROMgMC49sNs618WsMP92n6iR4AyfIRnpAAMjOU
Xi1YWzDtCak7SBaoTLWTWT/2CIgE6j9oGO/XA7dYGBKl5/dMpVhiC/0Y4ESWooe2onb1foHPfKpL
yIfM8V3+B0mjN0xKIkzTFA368z++MY5O1iMmRSJyIeZLWn/I2jKTOF5zttCkK8r2qt9nrHx8uf7X
rz/i5dMzyxdfajhHeDY1C2jOvLM5b5dSfFOUrBYJ2miSmPhF6C5AUspqRm+WPRyjGpCgGT37O57m
3P1V+I2RBcuhav1rTRs1TDHYC2BGlM08+w8nVrod7YGAVEXcWyDKN+z39yupmLchBsswtkmTQWQy
VP3cZ4WmbeENkWXArPYTnls3vzS1qiYssZOPAKJYnr3JYlrRSo2s+OYSk8vWFgWMUPkyvQnFznNm
f2gL9drZIVfpPsQlgq1qWjliWLDg1TBOF9CGuyyDuM2dUOvr/x9XyA6hux/btOJI2Na9xHgL9ULj
v3ScJB57/ypVS2qfkjBVFlH2I1Q+3UTQC4iZROeolOrnHnr2sKMrW2/DIru9eL91hGnLMJxQVlVp
kYAJ4KC6XQuIYkAI8KAzGXrrhiK9mXPX7FebvNLIwvuEOmJMuCms6FRnS5EnVlVI8XAn9P+QfSns
I06tXwMe7qafJ5sIfHY8pK2ok1o3IuEH3Yw+BkogyOVj+VTbQ09SEFd7kZl9Auh1jjRqlVde9ayz
xXzjjbld3OmF+6UHvMyoP2bz4k8YqPLadOpRgVopfF5q+5V4ynm7zT488EoohpoXuJ+3688l4mLN
7sv7VjC7TR/keLf7eqzCpzj2o3bU+g1AiHChTyfyrCIS1ZUphHcW6fMViCRBFISKPjFSYoC7hPwH
nnwS7RL3QTg2ze72hi8EmLeP4sczAjClglwie3pwJIoIs795sujM0+u6GVTAL8CT/Yu2qwAlOMDb
dOE85wXAzVcxda72bMt5uJAv6qWHFtcYHRhCEPUzAMaUyiFxnCvF2CE0l/HfiNHcpE/HDBsbAzfh
jzdfFUO5fYcuHEUOaIZ/oMR2oSgcZvNKhooPRTHsUloiPMqPo/0+els0BP74oXEq9wm9UNDRVKxY
ThprbHF5R2vXIk9KhF5VylNhO2HDOEborF8BP27sMjifAHZ9EQqm58O4tXoB9qE5epOe4uo6r7Tu
SiOkjxnW/YiHF3YuF7fGQRGV8UOnXleS6ovTyYiWlKeYVc6KN7sPuey6F/86AFhFVE8yDAdzm3d3
fGP2byAvWt+F3TRyyegaCA8+KnNwEgNDmPErWfZ6rxMoKFeOXb87nzqY2ksAH+xIEjfpTZV/JWE4
VtjPddLM3YsGIZjhALLJNmXGAQfU+7yrG0kEaQrZtkT7FS9jTGuRD5eMbjfye2smZpH3ERFHWb1V
w+RSCEEAv38nRXMqVcFGGaptJn3ILsFkfwqTwJcf5c5wqFeOyXeFIls5PEIUEw56CVeZF1mjRaUR
NCm5O06+6PqJfY5IxaredPRisggHWtEk/xurr1u6Bsez3vqHZm0UVNAk7pBoTQunGHZ/K3Z0010f
PYb17HsZCTl8f6vS6o/uj8jlmslzxxrzeeUqY/pCfuaLXhfxUE+3WToSU2G1vLwQIFTWzwQ6QXxn
v034h4J2HZ4hZ91QFXiWi6uDQ7D7n5WZwRw1z5w0SG9BiwZR3BfQZ0A6DMyyVHh1JX6cn8tS5ds/
0AQ+VoWqbSByQzM9VrUHzdUIZygCz6cqYMM/OXsARhEACHzdI55SPxD2MfkrGovCmXrDfU1wWcVQ
JlIVzrEHracL6gb8s0VK+CbEKArEi3thZmq1qdjFisjXmJJzKk0IX3fRZyurTFHCUt6D6rdymz32
JP7STwY3WXf41Dm9g5Xyk+GLVxbZAgRi+lp8ifa/ew910V/z2a3uA9ymcwkNCaQiDC2rQQ3vbIFX
u92MulhhgTI2YFRs1KvsXLJj61sieeyvcD3ZFSicZ+b5a9kQolob2kAHu+zgpHB2OyJfuO5WLuYY
FFK5fTc18/Q6Joc1A2Z3w0QubsLsI1EExRMT6BvI7RCu0j4HaN5vVXZWd3XL2JwTvI0JGziKuVxM
kMSK9RgZlL8R1uOCkqxraOshl2xMJGNwxKMLoUzCmDu/7JS4h5XCzdV1TF6r/I0nFmvmPeAILEEp
s5BeIbe7nyFrci2utbEsBALKm35MCJTP7o2LMzOZEPNVnW/LG5MF6Rb0v2gTzFl0McwA9lkL8ZFu
JemWQAp31Q8BHLVhtt1Ife07JETt8MEhHRwFnyYrDNAyjjTWSb161A2sFHFYPj5EFup9fKF7lwOj
72B6Dz5rXsFyMbzZbA/o93a9Dug7hTwK3mqknN8vEqwDybnSt9Nv/TiY/u3HE7SsaU0B4X0Ti6Nf
cKUB8F0KBd8gAedK983jCchqiWaGPDAZUJoNrsepf2ydqWNW9BXAaOJUzK7XTkptAS4XQfmZ5zxK
MEsnAPIEPvamxBGR7i3VBoA2EMzexCPATR5yoLODjIiPHHc9Yrbej48bXPITjFI90VHrgyHrnRJm
HrRj8GXuN6UtlaX4Dvkh0lLTN6eoMrzLLT9JGTNbeB17tWXv9IvKnKO9EzT/PDb3XxHQpbLO37YE
vcj6wQuou3RpJBiYG6ON+fWzsvfNvu08rl+9Nzb+ynYZpS+XKQQOcqMHDwo1zZOYDGwGdAUrg5+4
Dn+OjJdcsbUKjTlmioR4IMKx0Vpsr5rbOOd1g2G517yc8sqBwzJhoRYs505C4VWgs0p9Igt9oA6c
4mgaKFhXInVbs5HlsnFD0Uss5Nh0g+rtM+UrZ/9pqxX9o6mE8KYRqnhx4LzOfc4L5P5q7mxevCrX
4ddBYhtxYyy9/RaSB7+Zex+D0f08uR3NryI0lyVlluFtVAaNlGXq/yOhHQYJS3xu/G78TYCZD60k
k64vr1Nfd1IP/hAxWrOWSHu9zCtAu3OxGT8gvkZEiRZHyReXx9cHarr4FcRWHUwfCr/J0NwGMmcl
pi5r3t4LrzoVHBSOE6BEokPsmj44ttIGSvaKHfXLnlpqV6kPMOLw0rM8XLCSOHxbuw/9y/UeF7to
762JGpJfKw3hJ1nm2BP8xovG6xbO0HbWRzt3BQ6xPAeMLwU+34c/pbUN50tMCUv8CXSNSKjafnbH
GUoBqjOsxVNFQIkOXsAk8HWs5lvq3cI3+UI/1UuBCYjxQTtX97A59dL9OOdUZUH397RS92olhqFO
3NtmXJOesfH10Vj9ELWAFAT/XlBaCD3y2oBjy4aN/15g6GqUyJhCZQQnwp6jx+tb0azVDOnsbgSY
svdCbpyCULHa5Sd4Ps05utLVNBBBYZcQnNhewaJM/3kajbHNUZ6AJ0CSSsrnk+JgiIufP1FEJSPH
TbEEh/PcfVekfYb/V1D73p3C5JB25yGxM/9lKaMFiP6vPhmFa82bZ8gC9/9bhoHStcZTFeJvbLYG
4nqtP1hHMc4ZqDqVFsPA7XquVcxG0sal5yS8LPdDDSGPsnDAEdLqOmydswy6HvJK5AbXt1nNMV/i
hdeGt0VnJ3uPe14JHDH8j5AO8h8rLKoHJ1z/XDAay3rVGCEys9Yxlnb2SerPjKMIDEisqfxTKZ4D
vZdU9y13fR/AxffF+LzXFeewkginvy+/ZB8q/MdrvEKhfiJz1IhpR8W349cika5KfSrpl9C6euWn
tnGrLEwT/9LO1WBq10Oah8S5Dh+Dq+Dbbw1BYBmYiru1BmtaOkj4N7TzsrxKcIvD7psYN+365Snk
QJl7XL1/1kqGH1DiPw13nxZZGeWmkdLY7WYFK9BB/TGmZ04O+Pyahpf7ZyULBopQuOgr53Sgz/or
g3bdnf9LMwdQu4+Soheh0+VSvKPjIX5Z63KBXxsJ08jzzGOqskcExHecurVNtPQs293hjU/FVK2c
1j2CvumNW1DNilKwuE86+zQ1H5+omY0IwoCzttlCdenlx3PTqgUQIqrEQVGZfyQUGhIkNiIDLobV
EotbNYmC4NC4bMo/cUjP09r3/mIhX+H2w1/IwjSOJ9C/5h1DQUdhQwID/jaVnvyRgT6go28TB5PI
lI6dkC+rs7daEvubzk95aohMIqrIktkt/QVdQpLbw55oVJFa/zBNGy6Bug9UWDmnk39lpE/sL8wO
rrnqZIodYmV6arj9Db7TIlKLk5hhwZFq1vrdQd5mo9n0++MEIivehsz6eYgPNgPVT41RLbOvzNjB
bfiO5kNmu5TYEvBXhk4ImZmW3yL/C9Zrhz7zHNxIlu2C9Z2edJfi3I7CGN/3Njsq0mAVTbWfv5UY
Dnio1/lfOaVQc3SFN11e8wuZJksQgwcOfNP6/YcHbDzeHC9AoyQGIjLW3xM6NQHKdlPfoelkyNcb
VAdnsnzizRwgbt/jQ9wGbnRQtlqZg8XZlG4NOwAH7qKKaCpRd3YCmDKIe9LKZhJmoNFXvnnUwruU
f6u+5si1ihgY6j2pXyCtkHVZ7rTXrgmGCjirBDUT+fi+taQUDkGswtyPBTWC5QeyDbJG72bK5UsO
RD6s/pIrBT4JyIeZKJPWNTFYDM6tc7KVdq7cEcnHq7reAKSzHgJJumFmFoFWMdbODb5nk4yL2t2y
EXS6Ld4UBe5yUzRfrQZ86c0DPu5hZxGU/NZ0E1LAIkGO5gfjgnqDpgc9dXE6FBFkFE/PGGfcKTMv
UFOUxmVv2hQf5qdgfJ0QWNNAt/PBJLsh92nWYYv9Xn1mpXRjzUObgfMpYZnSIze4OwSj1xziB1Zr
CD82F+qx/sVcsUb1pjovr5rQ5V9Ksrr6t+gEBUdGL5atWJmPYwWtREqC7oeDxlXOTOyownDcgcIf
FjPd4EMvk2Vc/ylovCZUBzDZDGXv3gyrMZZWd8Q39nfwkNuj3fo2VtNpX/pw7NsUMrmkjztvr+HQ
DBAIVCyBMiQuhEQJ+Y/UI9CdtAX2FC4e+9XOEv+BmS1lwTO42PNoTPiGC3uC0VqKFAL9I+jYA9TQ
8pFHzA0bQuhtQs9pPBtoyavYaZOtpJ0odqtK6FywPxoA6S2Jca/BTCQcUu/IUFLn14wV9idFoCM6
IjkNisOeRQ0RlsF0iybkyWV1TtX3HlqlqP8dEWVnm5gb6I6LInYhY4AyfCgvqMqtsFCt+b9iot2y
tb9O3sruISrRMvCF91CXM2Rwy1ncPfb07+ERD7SQfrflJNGXQpgA0i+yUQAiW628dX++umPzuOlG
f7G72WAAQu/qi8z73VGjyjU8IW6kaBYtuR9ad8zYghFfEAWtdHNxqsnUEk1/7/io4x1lLit0NMpQ
xw/AlBW7YbI0k44pK7huX7FqdlWWieqF800zZX6F3oVNJyCHt6nUoQPWdz5jdOLawB9SYIjASXqP
QdKYtL7KHGPEbWyOV2CkpVAUv4yN8XcpNRxy1PGv6WbUxtmUXirv6lvAqVWVE4HFXaIS9q8Q9vWx
GTJmyaLJGWbV2r8vUuUdMr3muG3BNEgf4aZjJuU+QBzyn6LoQW3giBVHYvk/Yf6+/eDeVJJHI997
ktyPXR9uy8gJs6cb4CnDJDwVv8/rSA7DnNgXDsi2pZSofGUYo/6MTWtMz+ZjZBlgsutvw4WqTc30
PIrPDsoDNE+7szwQc5Z1drvR233wqIGQP78469bM1L42NHfw5mMWwAaz8t4Wfww9hwAZmZaTMIOa
C+fAQdvG6SXBPRCTxoGwzunI3nZwKvHSVa+CR3wGgjmkcckqdSJLDdCMeMOANjv1AbJVE3MGSteT
C8shj80RvVpSS8pP0d/cuNZARJ/8Vcgx8wcI4s1R2eWs91i5erE9EPuk2UkIcADVWfuv6XVMFOIk
KlwHMixEDHIm+obJrd3jrYtaIvz/m+bQMpYypLeWmwIn3bE+4tCUV9tRltO+0DdjuvLkoeHt1iuJ
KBizBrNxi9fHhR1Ey1QPw8eGFuQkeV3SE7bMZx/7XURRZr7ZQi9ynzb/+Be1+y+GtKXyQf0DHjPb
MEk1uqcPFeEIyZ7rHL14AULz430Mq5+GQdDlSfiSweX85mbL1dfIs21lbJIgVdPhnwafLrHAAGP7
9OR2sfwZaytqxiO7Xt7E49BvL+vHl7d33DTtvDgpUI/7mWzhcdiNYlUB0G5RJRjv7ybKO9ej7NaK
KqPYuhVAC4JajAJek7jFaZr5WyrEcEeu9feyXptaXMmCds6zWcFZOH/lLAANkpQvU5PPqwEroR+e
wKqEvB3dGlAQoaRs6IINP8XJHWP63Z2ZlU2Ix0kR5q+a4NQq8LXydzoU3LYjytepedaJiH5KjZU0
dX5vw4N69yiHUkhCW9gV2YzgH3QbACFr2rJ7F7Z/EQTM6VsPfq4HY0Nd3JihoMPDOYnprRReX/Xs
2N16hIrGeQWCp0WDDw74lvCPK4NA1uycddLMW7UvsfK9ZXqzRv5bobbXEBpJAiIAH/BSeKL4dyBE
iKYdcpCcLj6Y1y/HUYWRDB9hROYClkYI3TCEHLfLjxJat5/oJir7RsZadmBTL2cKRlH7nww47xDn
FOytJtHFpSxLfgW+YQ8eF8QiahzGZ8Mhzlf2arOOdX3/REwli26cl47tIskLPKbm9fZzD509uc4x
9k3K2Kglii4NSC0kwgGZPsSzBo6R2aoP9wZ7Te3xzspVR3FGC/HZYbNt6y1qqxCYt7XVVuCGjiwt
/NzyPiNoXX5zHFXG8QtgT/Kc6d4d20UfP+ccAe5Zas+JjKt3fJyY2V+lUVKQfouJsBy2afcVvzj1
FmoSZyfvwY/Zlv1fRk/qSODuxmECtdS2islGTv9+M6NeAq5OOEaikZ0hF19s15IN+X+HAbT+CE1C
4IgGaL8eDbCCkTL9xw4zZfikLoGW20pKezhmf7+wBlNOh8PR6KzBdYr0QlRdkSumlZe/9VvUHL+3
Y/MM+ksET1tZMYtNapyi1P3uIWnr+XBn6M5yZ3BypnjTZWzx/5Q6dxvACb6Km6CdzWAQpzbmrPKZ
EC1EaZ6iaKDmUh7z08knDyXbgzEboQuPgnPXWUBX39pOKpMTcYp/C66IwFjdn/UE2RnOrPO1F/Qh
EQjkHxk0UB4E6zLIRWa35AQr+5AYnT9atj1liTIHhRT9ivHLKwA9xBPNI19tDVjE0GYOzr1ulSTA
qSAu/EZgDAYDSd319eo7wC33pd07P/nTzvRbIzdLWD3N1Xu6YYhNTfA2izp6JTBGkA0Gq40Wjhvy
DB/mAsPyE0Mxkxy8zJGWVp2LgJgonj7tGrl2ZSFi+KsmA5talr2CjcUYd/UTle2CfD/ylGQ+6x3x
MBA93+J+aVFvRZNp9hgJ1Np+FQa/ljIeN5QajUObb966excT97U5NajN5ujCRqY9hvY4EnSj5LLM
c5MOR+TEbX6m7SFCo74GwnlgB/TvYFgPG0sqoq+k6jMkHFPOWHEd6EM2e+LsVKuQw2sISqBk8H/5
LLKBaWvhSBh/0+KAyqdtcTu5iotsPeaXCFpXMcpnkdVvpaEDmXrnpY4UmB2wnrCvEEH2O4WRuudF
+pnEOV4ikgxiNLkiaEJSrMITZG3haJreIwhv4qP1YMVC/lZK5+vtYQUVGuzE2FKliHjMhKBEBXNb
wLUhOfMGUhQChdcC70vPgoWN8gF60/Dh/F3EYjNqHREXRJKaf9x/8aCzIsfq9KScd5yEa9Si2kRw
PixhoQxE+2yxQZwGHP5xQPrLHa+Q6BTN9qtMgXZ5M1DtpgSzUWWnBDrLs1pdwMY3Nbpx+u3hB5IX
ZmtuNQZ9JUqs1DXFoXF57EdSdUXf5uWaChBmYbiSX1lCVW0xNut7j/tnbe42+8ibjusE5kZbtCKP
afx4a3a5lYPXvYegBV0DNKb9kJDA4IhKSti9WBIlbrFyRyrhNGSdMLLV1eklOlnGCEc74dhaTk92
WV9nn0QeaUk9Y1y/ufxoF63RmWPJaxpb8NA2W7U7NQ5rps9eUdM95BBsx8PzmEhp0WqewxnaOUPk
tWXwp3sJ8Fk6yKzvLOQ+IOHhr0jG4l2bvsBY9ehwKcvYO4FMgWcor2Ic+qc3TF7uZB18YinNUGcR
ecWxGxURLj/W86fOYwRUcZPB1z4O8FPIYkLeDr0vT6MRfFrmOJ9nhpOJVjZ30Dib6c2bLU7TrHY7
vDmtLuNBZ/GKUc64moeOZszB7Ib2WwkOwgcOK6Sjz8NOUoUj9VyMr6Ui3ZETfUuPjhk7LdQXazua
RVeQNteQtOFAbYpzlvR09ba0w+jWMt7Ag/X5zg2odiah1KMi6h9Nyfu2l/pIdu4iU3bcD1zYk+rP
9rIgogVvHEhw1c2lgZ9+Ujei+i6u/vRTljZgsuUeu+fJIESFAnehoczVaQNWEcb+sf1RjoyIjVqO
pbNsikb+tth/qMqR79/72AUGihfSxacmB7O0/JoajeP9rMBNZsuyi8GDqGXj2Ut9X/QO0sjBqYxS
W5/6zn/pseh4hQ+0PWRZzr93sNBzJ3+lH5LPmPZsoQZWtLPvKEMDUCncxdfIrngoMEq+BeCHGHUG
uHAySPuA5UWcpjgvjam92PyltdbN2bBuGxenP8HGEoVQV2s7qR0kPgHio7L9zlbCAJrAY7xec4fs
RCTQ8rkTJxD3hUSkvqMXkEz1gi1qR3r8wW+G8X5bxe++qfVhJbrIoctRWrt3wyHRxaMLB7Q+X2e0
ansFg5fv80IHzyzoPdCbx+1Lq9bBmZkeNLEhvbuKwnMZn6e8bNn9m/lPI9AsrjSsoMKp4Q/CxZZQ
4igMOFHD0k7lC1jKa0FlBiKeftSXgGS2vM2zvIasvm6YZCIFDRMkRvHCuajQZVjJJZrsgbN1951C
KdtQPMxmcUiHfJ5upQKrPQOWEZPHew54lVzH4Ro4Ie9KalM+gGFowFzPynIDV38+464QdLHlQD2w
r+pre2LYVKeU3aqtpL8zyo+nf4B/qU+YvpR5/AgKI5sdY+RWwe9ENP+rtnUabIM0WbbDFIkDF2E5
7LO10c7KGsa15JA6jgiC8g56wvEDiYgGDQGIDbXFgrbM4uc/S2u8q/pR2rocwryfYWZQEY1qK5JJ
sHaadJ3eSJyyvowlFC6VTuO0LJ16IeYcvUFd3M87+BkZSmJ8ZfjYIoDhZpoEtWAqXenBWUouLL02
CzzHeReaGcK41WQ3VSOtuEQWEeEwwu2ZfOidddEChe+LvFklbbgXFvFpgxMBrgmRKzzO09n/7fks
A++mr86osiILgc3rgiUscMy+1Bj011PK0yM/qlOc8HpmLD05YoQYbcnT+cU0zAZPs+GEODaEJcIh
j+V+nqAauv+drFPoI78ZDikzvCXoGhlhAxWU8zVwxXsBQz2sdOBctcR7kfyfUG20GbYA1Ffqr61m
5ElSguu/9uEcggitGd7p+dJY3VYskdp9lR8y5m4Xortx+/xcVOl/H9HVm3ftGOzwoBTp58METgFw
MLxZt9KDJrxcgsEd8i3oT1HZXLBwNVmRQ9t2D8Tsv6xSFbWNIY2aBWid20+dznDEW04+KBt9wK3s
KOTo56sCxIZoLrGPk82ZIHYnKqYZqqpNT0gpkxCrlW/vCiufTf9FlY7cBN/CEA2fs7eUmt0JhJKU
CX3r+3u4rxutnxG3eQ5gOUIaGdLBhAMXPMKZUwk+EN0/pIcCjgbi2U3wsQirjqCK3YMCscnCeVJg
c8yvBuOQ/nzrkIRqyl9hVPPGClT3bys/iLClVaaopxsg0Fp8aHzs3nsgKHRpsj6UaSheC2GDRvak
FdgSIM+wk0xiGbOwQCgQ4U8DfHwmgfW8YnuquoxP4mS9mIl3+C5vkXyDS7WLg6fYJ50Zxy9HBwoi
ah5KosLlq106MDdWSHIzvcR0IVqqm/GEysv8acHe3dxBpchHMR4w7YGleT75deGrKkwAkUEp9cMw
Vj6TkTjzRYZSZtcoIoNnWlYvHHcVmfSdSX+kRktzZpgoz2CpPE4NNqQ2ua2aFn9lVzsjtFMWsJ4N
gOJs8cSRxPkoeoDlpGv5DjfkqbpLSnbw0XdAP72r3aOFPraWmhqt4+uZvL3jjo3cXwhpkoYZYbiF
jznyDj75gWNbyv0dRGZGSmWKo8iWUcwQrSuJQEc4Be0KQBaVa+4RJJlG9ofgNPBHMxF7j/pBv9Iu
2GhxfjKntfveCWMv5Ds83O3hhfPtse8trgSxoxLMrzloTzRjcN4wzgTAxy50/X1CZgfZrRgXQP48
AFyewQAaEQsxIyZ84LAXQniClCijIWG3gAUnrIfBybd517Zo7QaxJ793IchAB+kVp6zi3JMZ1IzM
3ZCwBfM7fA8W3nT0LEIKJo/NyE9kjcXsaprQOPbJUXdQEGuKF6zKTTjxp5uawHIP7M5DFIbJzGMH
Vc4O47zhOda/fAqnLnyGfheWKsI84c24C59AbY5u/1WpNR9kmfNPgwE51eBOv7k/DjTBscZkFLtL
nPPGfUFVFyInkUjbj+fWHeUXSYhgsfoyLXx/A+l5vW3yMKX+YRxJZoflXKs6jQtc1ubrpDnWVHFk
0ee4jyu8tSmNEzJ070yjOFMbVAxq7Nn4BDaDaRUL1qUFIIfsgA0EazgO9GK0viRMl3D63rIoWPOq
MZuDdjK9yBVAHmjVk8K2fQA6jKGObIF1hSR+SbZVi9dyde7A2NZQsc6C8J+FZa7522wocaDCmKra
Bo8ZTC6hKMvSiLVztFjZ0oTnJFY1x8mpDvA5MR6U0dKZTuTFKbIN4iiNPm4Db6CyOEUArAEjOgHy
ESM2G0mQf3GKP6C/0/8XA4fHarw+D4sgr8ElKc7TBzYIVYNVxbnxnFKPHQDwKd7BLl85bO+7HMba
8KDrolhaXAjwKkEXNTfv7h1buwLcZZWtOfW+czw2/Q0zpFtL0DcqZOIeuM42Xi+HvUriX8WGDYuX
iwnhdRtW6p9STJRHURBag/KiVkrtAEQB4zCg2aGYFJaCCnNzOJ0iT7p3/LJJmLA4BYA2aB8xzZa3
ol+T/OhjpBHF+v8DsiwMFn1Yj0pMP940EscTzQ0VMXmUEHCfuDbpGYom4KU/IfsTd9/BLoA+OzdE
lyc2mqWRdRb26bU4/5+sm9XzUf/DN3Q5vjx8+9xKkNQPi7sQ/kW+oo0HNlDP8iSQCkm/XtalA/Ln
NWQhbf9RSsGArjZM/Q2wQjnawfoSuZTJXh0WGFuBkj69DlWFxltvr4ey+mO9GIkwZv/5LM4NnFHo
LU8BhYMXbzZh1NAWKn/ZPeAUvtg/VJYw0HVqlao1SWPdxoF5gth/eIdyXksY/S4jBroUx7GKYfVq
ikVSunuRwuMFeP/v+Ao+nT+D45y3is9GSif2BI+CWXar1VeaBDOtO/HFfYzrSzFzLPlILhxbh1lP
CCNHloHNmVJ9uRj0sbNWKgNZNGkdPB7yPo38Yp8OKGwKaeZC94WA4ph6OGd44RpGw2sNLqN4/y9r
dSlW6vUTdJ+MKJZEt3AvP3FtqpP+C7TkszUxTFMF/0uijnIMOV/NDtkmHo06+SnBPOp1RSzCUbe4
mJWAgHlTV+9JEnVuZ9PZIyvrsBayHV7c6St7NqrHs1qYGLV77/Z1WYeT5b3TzULWtX6aAaqoa4Af
Jq33JxNz8rIW2+yYiXJgg8HKaBvV75prbeRrJggWPT51K5aKYiIdwuus6uMEFjzPlcLPXWiyMPcV
P5phwxdPOfJPT63gnz2oDZWfmT+qHLH1KjPMKriAz8WSPyLw9d5j++t6s9O8Zr0FfBC6cCjlIwT/
s9r84yXwO9dwPjoIcB6N4AaoptNUeTjf/TUqxkb0IDT1CaxKFqjzyD9BCBSRHz1Xf9Ms0S/bxEqm
lHx4oXcpvyCS8gh98ejD4EKcjIciOzjfI++pnIOVRSU5MQb6O5AVaGcZY230UIDlofBvpDHGIbyB
BjFIJQBaofYY3MPVjfwidhCyS13+cAL7N6lHViTk7JNNPn3FWtqtrNmyI6HJbXnBp1LUWY5pSMER
GkdZxkl4yWnrWWO3FD6wLz61RKaeem21RnChydOMgYeejsnqU8IoKa4xCBw7zJLcLr261RWlZtSd
LKk6vyxU8lXGKih3cisNXzKI3c7UIbM4yXAssZBuFqYE7eP5h8Q488PAjzp/znZLpR90RtZZpYy8
ejTGTfI+MUxZlekFd099zKgGj/efdNAbj60IOzxYm5nyfp8EtFJZnVIExs0+SmSuVlYBV9JlFcwb
rB0/Xa7DBon2w4wO2YnIbzzkqSxAgPgdg/IgeCwcqnmdI/i4H5ed0iBiWTOVQ21XzU5TQB4OSnUm
x5eySPSpYhLxeDCUFSDuButkxZtiYOLWp9r/QEnfwVAgEUYNSjGJEV1zQoYvTfAw1r/uKHP1Ji0C
zPFQWBzbSPI+lsv0WKHeWYn42mAFFF6074hT18p2ZDHTuSkBsd8jmDPcJxX8wNgXGexo8e/dZqIO
rDZ4gkgHJrr1NrIJaW7SZxftjIV05fZEKAWAOtmCEOybGok4/zDHcLtyuGyMBEI6Vb2NrJ1vn8Ri
RpALR8AvoJMVX64dGhNo8NOZ+2A6Tl4mtpxGr5zwrqpCDtKHEfCGjnMOcS6dwxsGtst5ObT2or6H
zSYQs8LcTdmRIqY02QPEJAckoiEbu94oDe6bfsNDUro428FSmrU39mTXSvpz2TiCgskVeDdJe+OC
WdY1nFaJGkJdNP8jYZzJxFGhZ+UzMVxawqUkX0ciXpCAUQgl1ebkAQlH3hRs1fvE1/K0tayxshe2
qmJCds/q4pKzaWbFPh2yyuhTG4zd7ru8R6UyAKWMYK+uQIy0yi737KRAyjpmhunLOUdiWm2EmjuT
7tPWZaSO/vK7zLvqImpTamz4zSfeFt5CLyatYhBtwOU6sUoofhZm+ReZ1c26XohTNDKQ/Lg7bm69
vprzIu93LCXHO494BrAxqe78KgPcuLgGUfvjTloR4lPeu/1g8nujh3cec2yR8EGtqzThuyGo7iB1
75DaGXEa6v3yRFbUIXM+SEPAu9ATk9wRWOFXAAN5VGuUXrW6jfZgCEvio0bwkktkG3DjVgEFyaXa
0167QJlFylYGejIAONqBiwH4xcbXhKQXPw0Zn/u8oIvHF/Itv0XtLZRyNIIBghZBVs3eUF/f+xTJ
+U1qkn0ixbmfa6e6SdD/1FinHk3WJuNQFZwIIya9K6twcI4LEbHmki1yR57Zw0bfV7NGwkweeff3
ShpXXvNZoWFdNSV94XWxw63GvUQ+0l/B+IcOjB1J3zmol/silnUZxox7TJp8w+c6qagkWh/9QqSH
AY4cbQiyPVkbjVP++3So9rnv6dvCy+oapThL5xEDLDbCU18aiGm3sgl/LRvvqiiqj7+cWVGdMLYG
2gf3qg/D7gaIHzyjIdR5Vd7zqVcqHgDX0M9HheFr8CrSTC4ORnG8M0BVAy05u/FnrdaoqTVbVW+K
fxoQDYeVqO1xN8MX3B/tDUw7Dd3UJLnJuVyjqMIwaAVI/QofTd2FexvHy/gt2vED7M9D898BVjro
w3aopTRA1GYRbdIYyvYopBPDAYEpHVFToChZYftclhzfZRlqnu5SGZbTKkA2Gy6mZ9UUIa4R/AEW
Wm1GeFWCGlxB00+4pytLjURrE4QjWQo4zpBOVFYDlaQZJaPGJepqSCnvnRznsyE/5v2k72ZbsNzk
d59m+lE/SGpP5hA+LqoRlH81UzK7sPYnICnothcTmrxUQrjfwh0Cs77tlqp7jFJOQdIEb1lVgSBq
VWSWWVTAsqJDQXrS5e4ZmZHwMC4iva5GgT5gkkGPVd2sIEXIaMUZ+JSGYTxDos5mrN9A40v7gKAo
1hM1/OeRPx0UnrGo5M0p4G06vyLPPrel2dpVR+0tv6a4QSBHCI/D8T0dNsnV91eI7znFcFAWFWZ5
prtbYHpaqQD2hABLRRjlecOY2bfFUv5DUdjTbFlAqgci0eDLC3IEww83ZlZtjFJgK+2bT6WTcJDA
k3Ol3gIRJWOvt7jVfrRcOUl91Ny5chg+ES0K81J2LjU4R/sBpqmD2/u2du1lJ8EDsFasJfKdMB83
Eu6nQDs2S1Hws+qZh6s09qBdmphNA6BhBkRUatx7UIGNzgDuozYaTdeUrvtCV4ihxCX7ba4sB2ER
lleE+4pCwlf7iDyKiqLd7wYQ1bMhfY+yzqc7rZlbrsJUZ12KrTCCM1/LMOjYWEnU9IJR/vd53Mwn
EmJN/wL6BELvDdU6zFOTaDO5arQaA6KXxUctmYyeYf355KhRYQkdf3uuv6gmTD+GAgmodroJYUMh
OCJTYEC34OD1PJtJDPWW2Rh2hXdPank02dsZVTV/HOh9jSMqdtNOg0x4nnmyVLJ/bChkq9lHwCBL
5seFfFEbuXkMaotVrvoZvjaA39MmGtbwuTffknynfpJCNw3dgMm3SzPahoem7Kxp2w0Sca7p03Vs
2t3YqG5xGb6Kkx4d3sIQUAUW1gwz/ng2qPY1iyQ/xcYPqSWNckuCNQ2zaQswzty3tgRGmY9wcxFz
ub0U8D3Al9IIX08C9FSEDg8T++oVUd3AMsaIdYxiPntoq2xqCXw2LptnjrXmbuZRX/3qottIK+N5
NXbuW3P3k9KzVrIiRvgrMqKYGJCVcQ5YH4r6rU0EZ7c5X+WBG60xWVkLID208g3pDVC+3/zwUvRH
2Fc0qq3tFXzAVq99LWT+X6ahy1mpuIuKVMZ1WLtvjr4rvuah7eyxwGs+1LWtqd7nT/MlKB8xGbNU
c1iiDrxnGAtqAsKbcaaod51CF5AYrnHDbMfeHPHQQCOqsKSq9f8oTjzPZUnzpNgcsw3LwarMu9NI
8ZM5QulO+sc/9bikmxlpgAuHenwve3iOtc3b93mcfxv/ph0udvqhBys+qCGzqTMusE5EN7Vpbmr+
is2BFesk7Clbr1ECYWxi9gjmza70vQfVNDf89JaX4ZSjLm/mAQyuf97Sa30HFWlHxGz+ryuszivm
nggxyzSDEIgVAwm7077Z0NFtYKNie+69BuONKn6Z2pAvsaPIUmJdJ2UE7H+gCTH7CsstiMUdCxH/
/v05G4bGQqFnZuk0AqoSNtrgrLbvAMJYcf8uePj+MQmc9t6j9g9tpjNeSYA8oW+l/pq7jQ9eIISk
cozWtWg7Qo+4zuDXrg0rNZWDSy4m4yyPZ/6zUqhfwQ1y+wQvRgjAnYlxsXNsfxPgKALIdKHreEa2
wBTbV/jOj7gJlFjGsOMUzdmdnejI9hhbwz6TfPAKHf+7s8oYmpq1l97CLhK7sMlGrpqrV2w5Bnhh
admHvEhSqgSLhWO68ctKlRflyDcSQmUq2BJ65M+f2Dt8C/CBBpyJp+LIdL6DtYvblTalpLkSWFSJ
24l61SSVZwZIYqqZHZRleImR6uFg4ueSPuF4YtefsasTZzoR08G72D3D0208wEskH0Af7dymlwiR
ILY3VSqWtTSJDahQZgXRvwV4EyZ4VnEfUrdnVyR/m6BCzk7ZggjkgKcbID2PnrRgXMXOvmhdr7/3
HjCDGoz57zfapk4BpZXUdvr+gMSrCAF4BYwtdOFPxC8Qlh85525aRqKzUngnrXaY9UOX1dsE2xji
hLuKtPnK7oIGT0LMxHFFF1pnWXkKiPLrBVztg6iFfy5A7pxrvi2edE9BIg06o2o92IVPPECinU9E
9GQL3fclHH7Wbqe94Cwe6LXtyFYQeYLLuoO1fNSpSX2QnuVXTnyv+1s+VpsKmE9+dCi8xYjQMI0K
xe/xXhVVoQhwHT8aNmaE7SsghqS8NvdmGdw8FNFXzps9Dr2BJ4LHl2Aj2sCTsjmugZ9EveVd16cM
lU1SQ3F3NRsjvTtAfrS4EenZSQFDmKtGL2o3TQWOKsXmroEhUg/RjX1ywZ647UoVD4uCUQbuS1Lo
uqNMspZPFri/vUZ4RUHFXy8aZAWAkbkzYaCWUtUZsy756gz6Rj6agIyZaqjm0zTzXMPi75+3oXyP
NTsyOu+HFmEDli+KkbWtVebXWkv1mfIVaWWglo7cxxuCUYUFmZrMsYUaqbSQoq3DhyhdlXZmoGrT
nrwk+yPTqEYiZc+mBUeUqbEUuneMdU9aPFWQl7e60kjDG3Kkd6xf4HGIKj2qZgSjBWWX4Wl2TBI+
dPn0RLinzoxZjzAxH2wxMD+6olB5w5P5ETtHNtSMveXIEl9om4ul3G26fGruvY9/3HU58yaYvaMT
2dBwQhJTbJ/gNBEamOLkvVwlPH69dPc4RcDcruD3yeLpZ+SsQXZCoZR/TdIciRudnvzZkonGzSIH
zrVbPdclnnV9Xw5i39GUTgdcSk26SmM3ZDS3Y5iOmuGyplxex1b19R1fLVqdj3iHDmSmijxqcDvN
IQg1mRNCLodtTrypUOCagPGWH+Y33DoLR0NUQaH/+WwnsWXXb6LDtof/zq4FtoI9n5Wfr8Mi6zWu
62o/Is5HOMKezJlchxqYqsJMygBeqg4jAX1oujweUN8iZV9jwHeZzgZwIptGctM1+DzmGBbmWnG+
q9YC0b+o1RjLirgrtXy/MKdhmzvA2cOy3Chd1VHxFFEZQ3bX+VswOoob3eYp+NTRC85ZQ/iSDYrC
LzeeKkWaRxtZ+5TL8cSkcH4onlrav5o3rhzamdTxRqnt1vJUyrjuXSaQirg4YNBjG+4T4zP+U1H5
nrjKaiVkvaRCk7V1DwXlWZK/KJICIlloUfH+UYrrQFnMvT7z03ZFG3bSlwjzahDNegnZ+xcMKvhT
Jbd7hZad/JaZdvnAng5Jl0q2/v7F4pZJu9ZBXvJjsS4VhkdixYpcsI9D0LzypvKpV/7vtOTtcgzb
+nAXZAjgF7hwz0h06KjPNYhsxpbRVdNY5YNkNsaMX9KV7c76j0VRpyOy8FJdR1i2NE62zYrz9I3N
UKR7fR/xkvX8hbAm0V/oj7d/n0Hj3l14cJSUpJ6WyQikvM/RwnLp1vJDohxf3cS+Ctw97qjl41CG
qWiGF1AH+gpb5GfZM3X/hFmGKxgTpWiamyc3i/mNkcHLS6etOvWG1Nd+MawaeAWue7Nzdnxedh8t
m4SkIE0rQClxXJ6a8oMAicrSAm1XeloC//9VRKRkswinJ5Om2KAOv3Lg6dy81iEOFQBl5Q46Qtd2
lvPLLQxMCnRvTXuioRrcFtVmA7pbFRuv2ZycQL46FquxUyAAD8/SZPdAalglNwK+J/AoYovpHE5u
n0pS5aoXEcU60eqIvbVgoZtTKn3MBfVsaaYGWX4weaOonZom+t5PZBIXYjVBlRSNAKF5hXALB+iV
N8h9oUNTS/ndt8GTD658Hof7daG2pokD7iCNYN+uG9aPaNKEUSFk/bjnHXcWZtDGMRaftMUTyXY0
id/MWIdSCFAVgEf5wXjzA1r8ELTcfjjnSkta78S/lPVztGernraUYzI51AmLH9FKpGxO3oKf5tmI
/62xJ3Tir4fH0ZsKWLUPCfbPX9DrPWyRWqzMjCC9aKZwojB7wnUT0Pyv3maxwz5MZIngub4t14RS
ATokTRMylywhXX93UrpYhwOzQ8mhFSYQ5Sj3YJdbr4NzajUaHO6D5J8vcrvpd2a7eH2dzImfV99x
rUPVXs9/sSqdeN6V8WWWMjaULTgk2pMmNXGgjiZ8hhhzG7KZ5PDPnZgKv6j/j2MIKC7LTUEsqAUK
ZlT7bSw34y+lY37zY9b0frErXOsngOQ3TVAnSYkJ5J7gQdRJl4AzqUyQQHAXRq856kh+i2rNvvA6
s6GBjNTcEBeq0zBtAH3Y3qvYYtRlubo3GAxNaAZG800RVWGTZH3acfAXC45ohwR+9N2VAwVWCgse
9nAasfonEy6R18MdJdwQtKoLbKil3jkp6m62hJwMzYkvk8lMONh0xkT+IcIm7x4oAjf+NDEp5s24
JRjvokt/JMvYQavFU859BT4bsyR16r8mjnYOP6m7/IX7uF4DstgZyr2qpVLJf0huWApl2br/cCTP
QEoKnc/abmBHMvqacm8CurmxuX324Eslpdf4ONcMqBIXDvGyD9imJZ629BoB++hP9rCkmCTlf6cv
UJh2ZOUaKdysLxBvEYRgupaCww/C87Ny9Twwr/GF76m3o0SZkWxfq7+PyWJDy5tUP9aigBryxZz/
nHWESSCbnn068aMH7Jpkqui3vfrkfxG/XLM6+VFeCux5eq1sysw8/T7k7P0ZuhDMw2i2+4K63cBj
TDt1dp0KsBYAd7oerMZFj1cZqNg5KhSsI2dOo45TNx18F7HBzJQ6SaAoVCPNIDY+tkMtt+LvJQhb
L8hZLlJcNwhpq4U3yFCxeo4ZFSM/AJ7rD7qncqSh2kxMg/sMtnjGoI77216LhdlVvBWR7E6fsOC9
iKRmEzx4ErOXHzGADxRGMsntcIzmwbfZEDRVyu5o8gkCXp+S2T2rQzyey+qm1uqFCyEb7tvsEMPZ
jVSvl9uTiwA1F0ppyo2Eij4aaJUbjKmc3Zq3f9R1fkKUWOKgvfWkA/y9Tm9D4d3+PgXuxTVKZB4X
qnLRx6soSkl+0jn3muKU3KdcuyTwEhl0KidzTN/Y0mG7ZuVHyXHxDbUGsAGXpbpLFiYkwbLVI0YD
SPTC1UQAzhZ+AiMUAz3UO2l/Of3Ki3W8Wb/g6MTmardtlotFAuxHhW8YTQbRx/D6IwIN/HB5Lril
R2ijDl9CJjgvgyxDSZy8UlAJpLZSWSSVFA+CdnmEw946AiIr7kvqKXzVQy9ZsxAhguFFzDMR/a1O
mXNxZDrkkHwV1IUNJ+CTABMtz3kn0oEE60I7s9bLz2L1ozBPYB8TeiXljsIkv5NYR9CrpvcYjswg
3ReYkaU3toOczRCArkq2hZ38XV00HcXIi5ItzDCU1qxKTbcurpNz24Z3fVPbfj+zGHmGVkKPvofc
grcG3b+ZMIK7JmDI4fZhEZuO2PAYkY62K4kxSA3sSUeaPXrdzV3EFuMJFg5S0EzYRSIKpf7cJ1Zp
SKlN3WQap4n8rM4z9eTPcSBvexYekc9cjLpi4BdRiExCzafl+mcIi0l8etM+CIa3PsQrQNQQWO7R
vTuBbmIsKN2mgCH5xNQBqsQVuAlLo/7YBRd4cCMFsuRZ8AVBzrMyLqrM3oSyK2aLH31aDmP1FMRC
Aqotoz3qbTXKdYFvR6PaeqkKloC3kMw/KRQY3Mhf0XWdAL1rXCFbHbvd/lfKaB8wTVesYKeDtgPt
Eff3qD+ONa8NMFPq5uvvRWWurcFB3KcbjwchhBUZHakxsZxuz9NlgmbLQa6ATzVnjsIMFAqXefG1
6OpMirt6lry4PrVksJD1n+POLJ2FSANeNMBmWCJKo4+ksfZq7c9MyOMiYpV0fPVaj5Dg7TvypAv+
NkFR5lruR/t0KqKxvzdkAkXYXivnRbdnUD1h2n0IqF2VOX7ocNWbNiYqxwNzoPwuAN3E1rAcY+iJ
l7TA2Wht8Bwt2uDpSg8UqEbDl+10Oml6YP5rTunGJrSoaKBNW47EtAy+17Yi0d2JAzcw0brSdj9T
olTT3yUJD2YGimpNw4BUV1mZLYkAdM89uCdG5p8r9HpE8dDkUF2Bl7Tm9Tbr7DzYpKdoEZ1jPfLP
uQEzwqzDX0OAi+GzGF4ncUonYAk99psgUyxDuIxSLjKflJO7Y+Db9qIE4JRJBkCqB7zYxa1yMcwh
I6ZfQ9xrDhO0zCCgN9Ty1ICDrXDrn5l1Cwh/UaEh799trnwVdgzPNj8qLMQV+fYaIG0QBgIoDlSz
jYzaAOGfH3DiWdZhIClzV5iXY7juPdg7UpmQyVnQ2ZgbOffgsdDPVAeCwI0sSglXDNFh5TePCel6
CtqptaLZY87wh1J4sBKm6rrgS7euTDv+hBqGq51qkQvyKXoghz3KImX52QjNJ/nO5MP4CJZJdQwa
wbPUa/uND0dfW8JSRpYwk4k9sCoGIkVnNaawBZFeKN4L4zvYxleaB4MO4WmKhVak/4DPnScTqfzT
mE9skmvptz2bnYKLml1jSj6YfsUCZXPRm5waGhHV2iIRv6o6DYRtvL37mctRnSFfKPMOjIQ4dcpx
KeoQ86eOO4JpLdmVQMOL/H4KpiG7g/kYsmW/lQGm1WuJ32yey/OC5uWEdMGK945t/Z82hfm9aGEK
UyV2ZX06MjWv7p6R7PtKTLwB1/62RIwHxo75wilarDYgvAhDKscl6MB4I4wOLIakQx7Y8VhmKXDE
c5AOJKIzSQ6ok90SFv9+CNauo4NWmZ7UMf/cxQrcVeCPcGs1ySqZL42bTdwp1gLhOkxteTLmkNcm
pCWASNWTV3oi3bE0U7hlKejVj5UkQg6aAJluSbLx6fJnbYYLCvnadMBZog7NVnSRzNjFyaSvdKxe
ntAsXWPKSN1VoL17zujjTYQFXfXhPVw1rAinb2fo5+d9cKBx2MjU7TCOgN94k0fBWChOmaZDY+wV
aDVG/52bvk2uGCYV75yO2tNlU3VBZkzsIg671JEXliW0JgZuz2Mmv9nGpUHaXqmUvYVeqxyBbIdn
b/+iY2+DwnV+7oD6GyVCM7qF/8Z6vwB2BzondVcBrtF/CL1fEwer2UpzVCX+Abvo9LxMGCrvV6Sf
OMaA5rWg7nqCEqJzaTptYpewvX1dmESHV1PZeN/AYe1aCw8tlItZq3kYny2VW0LTsNZ6XAoULQt9
JoE2ofWyL8nVVHqMbNgbszbS8HJsDBbCYmfkZoNw6H3uCfTSmiOpsNjhwbn7Er/CEctUuMOvkEmF
3Y2KHEWwzvt8i6M7tyNC5ME77LJIg2c9cTBI0aHGmdo2qkhFYCTQZmI7FvcpgqBw8d6ZfbsatIF6
xYcWy5rQUHNv+U1n8yd8fpkDSG01AqKdjyysOrBlsNoNYCVAb8odIzDhYsR0hNtwIAW3uvvB+nsR
GHLxDI/CRcH1vHiOk26sUqV9G4yGJ2us5t7hlCvmbZmnRXp/IY8rc/+Y92mQQoYYtb/LGMGGFuuK
9sz+viizY0EULv6fROXANBfPWWkHXfhv+0bQwYPbPpRMwwPFuEpZpuVUuKPesQal04CszwVv5gxL
V2xD5YtuR5SPebk3rFIyhXz7Xjz2lD2EGDyqmJB85HhDLAJDuVwoes1ggZ5/cNEcAEZjq9EfVgBa
kWwxZx0yZ1PKK5/9kdClr5nu3VOtMXoQv80edXbMKT/cGHOEwDprfM7fsAl9fFgduytzdBg9I9U2
ADuHcmnvP/TBEf5BLJ3rutC2fj1ZPDjcqygf/nhytW+Ah+KSi1prJHj88F2xWaTrSXJ1tEQj7jh8
UAocSqt+jM9I4N2JBFAqEWOxSJpO8QyRb7ca07gjNep+SvOT6v9aUegsFpzC1V5GLPVa5riuGCSW
KBqh0mSD98iYc32i4GCPpxvKQx/V/qqIGVMrShpne3/0gxXZumHivzvjhdYzxa2Oa7RaIUpAuUxu
K3PCINtLoAIm9NULqZB0/sHn88LobOJKFLuGDzHrmjRbudRZHvXITTyeWpj2trGkeAIwDtVh3EBv
xprFHEFxxPFIrPnQW4har7pzMrOB6JWrxl8X/4HdzuAYfx5SZy34lvvIqy3i7Gx8biXQ8DBPtqso
TAXuaSLZaIRRbBV40YOQGT1r6CXWz/rWt7JLbcsruThBIjaxsYoULBqlhBaXjPzvUboawuoW3yuY
IYlmYadwiiBrp1MHcV0cOe7zqmlZkj3/5L5RMFGVP/crm1BF6vc/IzCYfOkC8FxvLjvOubFPUC8g
gF0GLSdip3z31gHLT6XHRymIc6Rm3vIOAMKcMcTNCpBTV99nO8+lUVST3xx0Q6IFwZU8DPKaBbIk
fODaGPbpTDJVe1HXg6HZeTv1jO5pO9dL5STQVyv1x83i5Z2P+bc7yElJz13bSMwLnZxNUgrkUBiv
JugFvzSUbETi/Kg5P3ES+NyIdkAyLgeFBmhmrIQht5RvBgAGw8RNZpNsJ8lfhV6aXUukIOgzi3Y+
Vg8dAHX1f5UKY1vfaBFedWSMrZM6O2o20k7prYXmhlxo6vvS5lAMerR39+QXUT+E06qaEfie2CBB
3G9ZboJo2IE+PqRuhW/+ms9d7tq46PXcpo7qcPvWUfZrAgkd1oRWNOSWsrADG/6Injbm6I5h7QjF
dOb7nSpqQWpGvwYRHH1+JJIOAi49EoZZFxGskLOKpg2cHYuTG1tOXyAQCiw/eA+GHh0j+YvNZLfi
Kj1i6xD7k26q9VYtOcrLisYVXRzBGoRLfhQ9qVr8i/xiS84qMAfjjDLsVo5bi8Fm4dAiEsc8fTcZ
DJ+lTcYyjo+x3tMwIZwgIQoY1dKj95f/WZ+CHueIuDPcFm8FleOiPzrVh8Fg/Ju08FRjiCAEAF1y
33E9JSlaoa1O1KK10RXuWWXBPvRAj2Q2rPta95uOY2y7So/U+iTgFoqNW0kmyOwNwE7crXj9MKHJ
xXlan0SEZSIi0Qgn77XHKRLM7DWz1qsM81i8Uq09WiPR47Myf7EjHHUSd8AnV39IiBsqHKXzVFNM
ZL9PzptjvSHH3hAPPjmVuzN8By1d7RUfjrbQRhJQ6EucCsgbrR7Yq8GesFk56PYi+PUidXkMX4JK
pl0l1yPJaLrgSjeWysWkh+eHw+89h0LnJosEfhZm4Z7iY6kKDg4qhgyq595wXFh0SUe8nq5VEvdx
raYS485RiwpwVl8SmvOAgKoLIX3N5FHlQ72e8bPWwHdTtk3nures4It1YF+yIDI20CHGSV3xIFTk
UbKuxx5RxDdhxsdnIjg6gwQbsf7QjD7c/V2W8DJ9Cw8Se1UrxUNDnh16Wed6WXSeZb3F0aDSpoKp
UB8JlUYj40beMszlHXyv/jixaV90cAuWhC0IO1ck32tA1Ndi8RL3dtb3T0Mt+jMkEKqn9UGPrxxc
RPy3PZoWW7uyktw1jNsJAU+iJoOjW1E7UU6eHe87Fg66p7SMstkAjbr71qEIyouNOh3OCIMRWP7R
gqO0eOYQ50fu1VpqsySDlAPhtDXs6YxFWF2FIGc7Sg5Wf68rPfePn32aAOycpOCpoXNo91/BzMSs
28EOFzwzULE23usEvl/WMYtibBYUtvdM7rIFXuImP2K8yVv4oGt76dlDzAGnt/+TAoxs+caHEGsA
cPh5mdsPdLiTjsWALqHdOM0tkpii0dx61TYFIThmW2s2s08GoJA7ideN5F0NSdi3pgpbZGP/q07F
U3v02SjJS/1xXZ8R8UHfBZqIxG2UbI/VMvfXga29JvrC9zmtdvlgMMoSIIQbv/+4OUXTDPfBDi37
oIsT/GdJijUzdBCXLGtKDipm9k+1mY8JMQCDiVqFqYVVO9BfUKSN/HZ8I6ViWmKowUTHU+pV/izt
gzSLyejF00Gy2/X+5o4XP58cJuhL1cWa9AMqRCpEj50pQg3rX+hoFLkdIP4g3JmtLgl8JFwywEPe
C/vsS3EUNC8Nad6vhcvHdCjdmL5htxc3oasnkZVqWie6TmIjZ7yyjVbcg6B7hW7R21lSnr+/ewlI
s1RK2IHxYwBQTZmOXKgTVMFLzhAsQO7vFTqf80yHn+w8YHhmQ2xJ3ShcjfvXBOAec6txpZwJAxO3
Qest8+VOXZviF5RKKuZ9SFiVXYql8n3ozxpKg/sVApJDhtaoEmpO5WvT0409T+yvaUDfKssKfxDy
EfvB8BQWqqiiq8Q4Eh+LHeN1BjUDHo1rWEzuXZgwNhkD9B4xe+51Wl1TOIWvbwNH9cwy4QiCDs84
ZzNgq04hoqs68fHEUxV3yUFMCNDWIfo37sfReSsUvTXPtS8hkndIRWQ1IFx9wl16y4oexFrFJCJb
LXlLUm1VKQNOALYhHOL6xDabDmw5VCM4I6XAZUQqDRBLDjmTYaXdzTu2UDn0CgJ48DS7A+xqw88X
fxe9xMggDtuWs+pVEkUUCiLl0wJhZFSVcsbNCGTxDNaQ9EA9M2+x2kwvkU+QEQeTrkIfCrGgfcAh
w+gpB6ULtU7b5qmk5trg4d6apVRebKjeb0n4cSyBszpN0fK4WXzPvcd38OJVfAlQRQMiT9DuOjaK
2MqAa8shvJLAtC/n3Fdu0ITQWFtqhF5s9WKbHvlrTjjlsffuLC6UfWf3f/TGQq9AhAEdTW3l1GJQ
rTACI97+v7nT71r9rPYLkPBXcLaX3dAMKLOufHcYTLMXc/Jds4HnPK9Xq+kDI732SHdR7Mq2p6Cc
UNnJNkDTbT7/noE0Thf9VtTfb1QHFLGr9HKZ7iXCHr12FZuoaRmjYW7ux8J2UTcIzerinnAPcHqc
260Hg3We/8tgBwAWZO2AyEOzZNWG5qjL8kn0NuDtdnYYm+Mc/EKyKeYJzSP7N1yhZijxY770gA/R
6aH3nbqaS9nKzDuk98uYUeRPqa3WCvsTPy/3CAv+K3ElyWRRVuHgfYG1mF+sfTUXOKFrmAMPB2c1
9WLvb19bgdDfIS1vRzejXwck/X7r0qLfo0oOg7plL9kxxRwNUX8ikPMj55JO6BWc50p4w1Af1FXF
z92TMUBlflJlJYa7sZiCkRhcylqiqs8Pwygq4IyeVQrgXvVSEvS6sbiufnQ6CQegt4qnxcXL0SlS
e3rA8pu2RP+8GTPjPE+kGyOPlvpBo7+YTDkDdbj+V8f9oMGUoC1OJx9KDukIKYpIpLL9FSu4LIBa
MDqobnyCarim0IN9+tfyD4YgdEewASLi4FblASYR6GzhK/tJB8Mj3n0TY2DUR7h0itdjogS3shcr
nH4GZ+f7wiYQQBihYwxtJNjImq8BBMgK7Dk3EmpA1SBwEV7IXYbwZj7/SDKydEBdp0uU6wy6Md6D
yeG+5SWCWIMGLlun5OFQjF6sI27Obj3PCObagnS+MeIqKLx88BufzwaIPmbCQkgBFO7NvE3PhPYG
LVUr5R+YDL+Bt/UDE4Tq3kvfkOUXCzXDBQMTXqCs4FjaDHpZYFxBreqO7SpNOiiV1h7870YlQE7a
OB1xAS2IYjy2tJWVqDnNfNdHEOAXPlYpC/ihqTE1Irp061LgP/Ibn6eCj2UqOqkuTjKq6er0yFwM
UwxUn1A5IcZqgoaQGOxXxkqXOogAf3PNgCHI5Pfk6Ei+MAG2v95e5RJvwW7c+2WnPfCsts1cV0kY
SJ/zS6rUd1MeLYvWQVeQnb46Gcwl1O6mkKqsHTWI/w2xTv6j4IVEXhPvzgDZQGiyH1oDzrt0pu+3
Ek/9e5ptSKr1bYaj8oGXygV++H8oin3X87OW8B0gq0sLj6ifjNZTkwpTI91ZObrQzQPLaZByC7Ko
HLVK1d+vpGFiMI4WOkzCYtfKeYZHGWk9fyekxxZ1zg9LYz/rr8P9+L2zZGrA06vYVyKqrvXJRwqD
Jsb/iKOcmkM7DEX3P3amTTDswy/m/nh1LYA/aX+g+6U2cfKpqvGNaeBJsWQRrNnosihbIlfuPDHF
GxfMjW3UvsvRBQkvIb7JYpqti/I6oa/C1+hKS85awpjaxi5ok02bmO1DKT7D/8pJC537e99e2yM7
V1EhmEFBTU82dCrrKlMSdnXAxdIWyyanNevgM6FdUKEgIVPyqowaz3q5fptdlpw7gtNJP9IIliO1
E8H7/aXzzmYOGWnebeeSP5+jDkOnjgooBg/FLMbad/5XUFFj+1fMsTqkYEYrAvxEpkJjKjR6TG2c
YXNNZln7fFHaX/GALE85i1+5BwFeShX72fdxewav7vOCc70G6zLqQ23lLHnXGOhA8BRLFNzWExfa
Xq93bgq89qBO5Zrr+T8nMqkTltz2bD/CicOTfgx8XQWnGd3dnx0N9O6r0ngIRhpzevVR2b1vq0YL
/cD5oDM6aRX1Cdw/3IF/2b05ZC34j1/0ljD++easDMpmyMLUFgEWfbuoqBHoiBmjnU/Oxn3Sy6zn
T4dLQ8tE5fu3qPauEwRAMRbZ9dBV2hN+fh/dR0+rLx90H5zkJw1UC9eOk59HDTM8YPDE72pHD0yi
TbC5QTw7hkzEE7oY5CdcdZW7csAF92h1yuK2TslgPFqGSZdWsoWfHXE/+A2Ix7wOVkjU06/ioFKl
TpmTVScQ30xMnnW4Estu9TtjyMKS62qATH9NnuHflODmMdV2j+QvxotDTZCblYg74Ws9aO/5ttIF
B9rYBJatyiHh1Ak80GBXbiFp/kwnq/5w9r2ddcJdMrWAYpYyP7vDS8Igijc/k4BIGt/NZXggSubp
HXbY69uAB8/iTtk953X1zL6p/8GRSiK2tjUBxE2/qOvaC8iMcVOorDcgxkEppQbnLetujwMm+qBC
5bjn0ZtqAPnq7IyQAffXi05Rs/bBCOIGTsVQ8juwo5o9sD1AbC5PrGqKJYGi15dlaPjJpunYza4O
uR6xOS2g14J5diV942b+gDxfOLALSMSNd/6VdZJdmUYXzucWVYu/hhpG5Jx3b/m9Jcs+HVx6BMg6
C+GlKy7gZgF0F11uxD+p9BQi/+a3lNK5xo+Njgdd2isxu9zA73cFxZRm5Fjp5CkUeyEbgeB8r0zD
uPl7uAwNrnovfViia1eMCKp3QUWpf3vNdkolx3EV/TCxFKeVXz1S6iNTrXreHhPn6q0Pk2YBHuhf
EPkpjt77EFxud0TSndKsJLP/FbYsJZT0qmzl+njB5TfEN88vta5MPJZhWQ5sOVInbOGYGsLrkzu1
xbb1vUzCct2q8T192KR1A495lO7a1kGlUKubuwp2u1Bvgc9J2WnvJnYmpRF4upAl8HeBHiFUM18o
f79jeh+BquhUPaJ8f84MRJHyYVv20GPOJyHiCyitMubCtu0Uwkv2hGOiQumDTEZZKVv33l77BUvl
MFwHbhe0QFC3yIf5RcQG1f7Tr4807L7M6V+AYbAaCwh48lEdbiVFrHJP8A5ieaj2s2QpqEspjyqJ
Vq2fipJfOfmKNjdvwofUxs8agDzEY387OToeVsOGtaBSYROcaT1SxFHgzSzKCGoCGEbn6Hb6VP65
1KxqIpoU9h+X3lDnVSFI0ZfISFihqp5bo3+HlYpm9i+RPLxKKb/HpAz+jV0MX6TnZ94LPs+/543o
QYdRgh3wQJHRswbosXmhzddA5AfPydvOgoM7pZRpJYACU6S+gg6jOqZ7IN3u+eKmQhPwbTR96rxT
LsWzfvER9cCYSlyEhldDa8VOwuxzo419tlZZHIiWzpzIbUig4DAWhUtMFpbuGEsFoGJt0KPvaNal
J/nVue+yLekbtBdz2oRGrn2ybasvGuJt2n0KAHuPuW7CwgSmMg8MwAUh+MzHAJydcRo2/dC8QukP
NNW2JKmuejBTyYQOrJMtrjyN+kCqqHW//G4oVNqiudUpvOOcQvAp8IrSvJFwwvPYDW8WJBqd0aQS
3hU8Qg38ZPFQn0K2ezeGPoJccE05xV6WAob+p0Lc2urQ92B5l0MYfhueb+AiAsMMeUk77w+/ZLgR
hsyBRXNjY5OhEpGUe8gEm+ihZzQbhRL6S2JFlfyPX3pc75ghnXG/i/J9E/4yYAlfL3ifl0rqKB3Q
zR3+XRVoH238d+hRw+HAx4IBjmUa9N6rblQR6A9c7GX5biwwR4Fwr3X/Eeq5b9avllpAz62fU7wQ
bdWT2hHQGXrJOSYdljpvZBiaCw3uWlQbyNYF2bH//9/NxuLBV+Y6XDGwWWfjbdBxCZW4EtpmV5gH
dMhgJdEbelsZRTmSpkq82SkVhFf8/p2vWwz6mow3zZev4pdS2lVo+nMtQeNMDE0Wr02THKSRp4fR
Q6LdsKeOmKbO5Jt/NRJGVWMZIC+Ppvo5sqIvfKQ55+T4G7J8Kuhol3XhWCcyvnDt4LMotU423xdC
ZwO2sIAxR2VcPpVvfX+OAb9jeA+8HataxwIEDBppSzfAWDVmo9/EFC40u2XSh7dvP/fczUcSOMhu
YykyEzZOB5pwZ16Ftt6whxRRbJ+7qsjSqv03MuhtRDoNDp5xlte1btC/ejRXH/gsX2Rwcwod9prr
10EEvzpcuztxze+xbvEXmIVdfl+pCZDAmDHdAB0BpSuCxM4gMmNmzKm6oXC5CqwPvPNc7IJxAFnY
QG1ctCMx97RuFcnH/JlRwSO6g/Jp6kjDgFrLnxpbrnAmN2lIjNd3ib3HslWoELep65IkewV+VrG6
kGZ37ZiBUtFvixiuEeuf+3P/Y/WceJRsCTKM7ePQyYE7CguqxOzR6ThQR2Y+eF9+qUc2tWUriIbn
kcIknGTH2A4pI4/01cViDSEHuP/0O1s+Qbsw04OXvtHW328Nr/0U6Nb8y0DAZEDcfg7tmGpglJP8
Tq+YfuP/rOqBBiITxku9/5iL8ZDTGUE81UyXDTAUxG+nraFHLG151ltK7+kGGIsM+y8q9DEaytFi
lTTvxzcBzBht71MZOyrpb3IlcBHlxhl0cJzRcsnboK4FhJUH0bsLj4T12nRlXTltkdwC8sxy7+xo
0oqJyg+ki94rwSjU7U9extE6M+KDqHbD/kT8yBTNz8TLinlSm7rq8z1yc12suwBXIXDe430yuLLO
azwzb11Cu2Qd8zerPxxqY/tPCOhL7bn96ZuTZ4cEMWlcOg2nzfkegjXdjRaG+929C1qHGtEe+u34
r1jsMelapQKLq/fyRyHZrpZg6tBkOCzkkHSmUj6Ij4nf/0V1M6XwbMsl/8tXcrCvWaxlHQCPGmsl
fCmjO0UIMyNkugqSZBX2QdHsgPpMWlyh6R/vK/7h+gzsVpyiyS+/3UA6igvqXYWOjosDihSnK72K
rklHK/LgIxRseCC46MhEVnTClG2W0XAnAUKV4o51p7EsQblHcTTqYmphsadem3KpvwJKiC6SYWTl
OFWCcB2FCR7YwJMvhhsvhFudXIseXWojP0qLsiR0jkWTZS4FwBwE7/B5AFnW7p321d6VXgm3QDs0
vJ8rE6f+ARen1ErAG3KBxqt14nPmLBz4A36nh9C4SpSp3BcdaxkbPhYBS72WvFmKLNluMC09AJb0
+cfXaNKB5fpmIN7SEKRJXXGmYxdGYh/L69kRl+lQILJ5+BkZzChpd3sjl6iUzKJ3v51pX33dXx/l
wM33sZxlHctscqi58QQVkAqwMIctBqTem0r5wvxLwfhVIbXw/rDxS+KX2afavcgOr6X5QbDJxo0N
tLy3hYxhRMEQAXGB+ZRbLaiQgzwM7Kafb3IVFyS2MCykmjmRp/m75ZcVW36o5E8j05zF7SsHWYqs
wvu1sqgsEgKttXqm/HJndo+lq4wlckNk6xJCa1INDAyKeH1DALFSRr7mIazonFWahtIDDm8Qe2CF
ppT3WbgRrlJ//N9IzOvChMUYJ7AZv++qBRUy6DuJIFPkfowgm3Tv6FRAoGkAyYdAVm3UmWxRd+PY
1N/ntnY/YnL6L6DykdPgtDDy5+dgJsm0brP2+PvmyYu8VLuPqqU1WCnvOUi0bg2J0fMAHkDuyOWN
D9GB2jt0Ol8K+3GxGLmFDGalTjCfQ9yInluZMpabOdOVwz/RsjxZQWPxc6OA07193eDxemBuJH6+
blNB2EZWkDG4GNFxkgXSGKflEqUgS25Q2FtAlvxQUlHqUN6HGGDSAD8ExmBcDFPyYS7Yo6Fs94cB
4Hh43XqYRE67XB8Ie3M27yYZFABol6xN3wOn48sl4nAAj+1CwF8tS/hX1DEGXryV3nqNApSvlZwJ
iHW1DCFydYyybs9KgRb823Buy1aniaStBBEd83C9DRb9JJOKZNEmdP1JovxDlcSMRfN7+2O1SVcw
RNIixe/HavowP42PEw5Ncom5a1/iwIoH1AWc3fCsMo9+kV7I3XyXZKP6eTWssS7IJMbp8kBqkrmu
loRGWw7r2Mk+GwigA+BiJBdA0ARwSeLvMG/LqELN94jUIzR4Igc51U71ufOlbiMSXpHtUAhTt3+F
F3pAsRoBtBNTboiXSkpMvLOoLD0cTq6KnJpt+wvuyk98+tYL7t7ftTOnLb0ZG9NW9U/rR8xXFdda
G+F94z4loCsohTMFREkgUz/f8TA7W/mliKENE6wNbAjqFtIJR9mlEX035wBzgeOtMj1f7OqNqEOA
UKixPhGkr4qjt9/sQCWVe+5Ro0RSNteBUFDzzQAy5W5/2ZpBb5rK7q77HZ26r1eYMbnua8nLcYiS
sotdluSnryLmd1ffZQCXbi2itJJbo1mJGT2rpNeALhu8Z4js4a8D1Rnv/mKKJWZRz54Mx9ja86Eg
NfOnh3UTe+83e1JIhPHPFK80PvRAvpAwELXlr5O4+tDXdGXFkoUvQwQTLVkEGaqXPbb3QPoR0Kr+
b+oxbtrUcNCbll3YBXQe2d4ErTiNKus/MQ0UHCQTZTatLuoifJ/RYh4AvcwQME7V/36/X4w4WUOR
jyaFTaPzLgHUNlCyDEN+9exaSiBEEUE50qCOAertYPK3fxoGGhT5jujHRkB5BqTq6mqqYrtBRg+Z
2AxN08l/S4bRAtLd9H4lsKCd/rI7YqvUlpQeFuYDQMIMHrcnixQN8hgjQfOKK9XaBoykJ0yWswum
xxyTnTbIS/YSrRKdywvrm0icgTgN12lQm8vsiVebCEAO+BJs4aH4NDyuDS80MQbgcvEhvPfVnPmp
0wI8eGJgpDUF8Ojg+zGhpq/kzZsjlB5zAsLnRZVx4J69njBgJUHYK4EZVz5Ja08SV5Ky0uPWz/+W
Z+O+wEUmlXSbZE6iJiu9T+2xqg37OQrjXLtqi4jWXZVf5y5Lj9RB/AE7yNLwpcGedExyLAV1KSQb
ETX5+09MHQYrYmVyQPUAFpk4txkkIr2bfBmHoIi7Xva3gu/qeP4gxuqXfpuxqdz7+NfDGcjDdXq2
cfVyGKDiChTlQqTXq0C5Ov0eGYQ5sm0HkxZ1no6uRLrKvaxQTRChfWsMVT3/JUWF97bKB5pY00Cb
cW/kil07epbTHtcsb8/GEPlhv0RmcNvEcEdkxGDgomNCxrIKzR2ETLxAwB6BxKnUcw2a7RxtXj1h
cZtYEcz5bwFoRVbNh6AADqNka73Hvne9GXMxDx156/UIZeH0tWXrxCJP7+Z3s/BTlVHfZjC7SpqZ
j5NnfaSvDfZiT7uRD9uloy8jP4bZJFltYaynHhMiUbJRz/vm7Eih6l96iYTMTGM3tlcC80W590we
LBxHEcxYhXVbmwM3G8ZwHYvZpcb4fOs6OVPz94IhrrA6P9pzrhwzj++5g9zUqYv8plMI922E0pfT
aAQ/BQ6L10Tobh8HaTcjMyuUAsrjmre6zx55cxbQr9P5Xq+lk1JXVHPpvRSjVIuVCRD5c0rhFhUi
/lPR8aD/ZZU2ljV3/7y4WjUU9rEb4hauipRUJzb/7Fk+hLRU2ppTrXgK2XSPC9D47l4qZAsY96MQ
MbDfBFYzUVhMT5Z9yfcg7Zuy+NKxQG/iHxVT8ov4mY44j/3mjTLSZwIEP4UJ2ksoitO3gT8Dpv5H
TXfxUhTTG073yVvLSECq2o9KfT6c7JAFAy6GIyd0iUOWd9NHzyZQxdbcM/h92C0Ho6AumZyvB1yi
K8WmHRAoh9HpqGwsGqJ4I3mTj7T8WrhE6Od9LJgKqs2GA76Kjvc9Wu2y4TqsNMKjjhWYJr2vEvCo
3x7HZXr+pbPXwlkthIgAQaveY12JPXT+nu8d9z3Jye8uFSMWt5qm0Z6g++HXQp4v20CYt8l5XnSJ
014qvgVNUNQSm1ZODoYSZhl8LJWm1LCjKVh71tSjO2y/+0ATJF+00xPOe+SknGCy1YGJe6zU1oCS
5GKHNgvBSx/z/U01GYazXX2PT2WW5Ez/d0OLCRO9XCBZjpa+ns0oP2QEmn86ntmp/SZWwPICbBCH
liuoW02JZDVsf1a5tmAwLHof3k+k/yuMKLh10q6gAEQpOvVSVUBjTcFP57IcKPit9erBufoc3IFU
N4VvY4Lz8qu6bTTrdMkHzYqq4yHpoGYfAZN+IwStqzs1bu5fHJwy6UA3QkWR+wsOR5CGL0EHdJfw
dIgQK9f9m/f6rJpNKwqalt1OBEYOjQCg3sYM8xehpCGOtyV7YXQ2aNjT86hQ2OWsHjFs/8yezlcf
RZ6FvGDZybkSIhQbHjSsnccjerEW5S1aTdZwB3MtsVi+VkKMf0xNHLn1T9fyWpl9h4Wtr0l4lBET
y9UG5WNAyXrv/am/cN4oep/83datX0S5Qp4H3YUlxcAnvwWmXo+rOY00Wx33HfhAVooTwnIEz2Ag
Xklj/z0usdu6v5WvuIs+1fbh01Mtko1jz+s+JQk/f25ZeNqnjIWDID1bY8zOVx7YytEFGHmfZ31a
oKRggwSGHMoWXUYLZNodtH2x8asA8Vi74iEKNSYDuJGmCx6QIfzCTas3bh6hFFDVdk8K7qf1EUv7
vJen1jXO3RI3yGC2xMSsErv7i6Zq9if8FUVl4dQ/UNAzVW+6gqJIsHIJgltGCt5uwaBPfjJMV1XZ
MYxG8VW8dNv3x2V5ceq8vHpcBC+fHuypVuIMbOH0+rtzXTmBkzJ82Jb4BU/EtDQiMWqAC2FegmF1
Gu6mChWQBZ5VyHH8AAVeRlvU0pQMbojo5wQyfgq7O5jmir/QDEd0iZZlx76rjKdJ3/iaZ3vt0txX
QhCEd5AnDM7ysX6kaaHR62z48XjYBR8i5kd1r3V3SqbU5dBXpaFlA+2d7q3ErT7cX1wU74RQ1iZG
xhUXqOfgfREPlnHz1D763Fq489no7jTnOe6kH1mI8y1JGoVGVdI69W9irSPmQ/hffH19feyZGGxH
m9dPgaYJE2P4opwIn/rLqbuIHGoyMTzEZXMopErRcN4/fPfW/7ADvv/VPi+bh+l9EJLZm6a7BCjV
piaeZIWjawNE7CUZH0LT2KoR9QG4d2xZNaSNpiNhOaYI6gvKUp5hAJfhz1Ihm/1Bqlgs1N1RYgSH
xSn8FkLE71arHWpY4T0CwqYg0RFzHdmX5r7mGtuA6MTSe+6PJF6zNQX0rNOCuzf7OP82vpxbNzu5
EwE83GEvW/+hZH4nO/g2r5bYn5oTT3jBwCOu7FXX1ZAQMvYXc8vRxCvVZzER3tx2TwYaqt6X+FUx
90ZaIjiQQQUp21okxjDZStVcBdWBPlxVrjNXyL8GW52NnhOMki3zUeeOlw6SGcj1r+Z5XoyLvhFz
K4Aa/U6g/vaZDzo7YIO+Iq9qYdSb8LiQfwgTqpu0lRaycEq/uzvhjxv2hkBKDlW/CUVVXVhS96BB
CwU2HAlbp+JsOl2CZepH3UWPCUNaoo2Sh5Ui0Gttc7kKvyWitVDVA53xS+EEk4DIHjSDKKFWciLN
BjtNKqTTdl7XDAW54AUmvnaoSgGxbqdHwpSbqRWwYpjyChT8H3scKcJA1cSFMZFDESDTrdbNeaGI
gx0YIDGKChVZRCBXEQUDRLc7jbAX0RXQ0Ir9TOLpsU3Up75MhahlEy0qmAwQR3dJdU5BN4584CJW
RmJcIXOhm4SwiWov/04s7XNPt5Vlta296TJqSmbiZTjj7V+wyDqnAfRg2ZxlwCDUzv3e+J6Kkuvc
KyT7S4gzo82jXZdJo7V7Su2uck9kRfKbYGQGvZ6ImAkLPUpPeHTfhLQRFPr3PhTtPv/QBBYmS7fa
NIaYbA7w/C1A+jKxhVjsNjXkiDnctL6aR/nvqpkdlWkvQPD75XIBx/ZmM2mVPnZNjxs6VQuMJH9P
GIvYzYiq1iTGiY9dn9q7/+Sp6MpeKO6Ljo9bFzc3Vv8+rT8qFPNhN0FSOTufDAuP5QJpIdnweSqB
ST29os0CmsHJuiFPoJX9+gE8NYhOIm5VwjQCEKcwveI0DyDsxURwhd/vwnZcR442CFmgYLZ4QY7o
Cv4rjm/JBgiBxFQ+WINon6lCYLqVCaaaJFDZm44l0XF65wzO7V1XBGXQdRzGTiMnwrWs1krU23P3
ddYOmkW7xK250goam+HSd6VZcqoygHhVHvd2lbRx8WzUsq1RSmFNBpkhHibuT6nHw3sbIm/f4vDW
/SxTO8aPEs/XUQCK2b2iJB6zWfFnt0bdgyyEuq7WU5L6CaTAXc+CjDbplJSG6UlSVM44yKtoIYsn
fTpn1t77Hq2Jw2tNx4b0yhwpGpME+dgepqTLYj3w3wsXG0phFV8GfyF8Qgsp5cxYHkQYcbgSTpS/
ivRGCtEnRScUy9wl04JNhmMPAhGNc/MBvHShloNInSYiPHyfeM/YcnhBlGkZsVJoEuc4m6Gv/vsD
Y+VSohKI8wy6QrHctagrsRve5ptt8+14ZMgE/2KYqRcGfC8cA+jW7kGW6CHGXh+jUcjnnDd0d4VR
58GHwCrr40rGixGSU0cckRUdyD0NsIHcpPDYVlr+C5l3JEiLv3f0pJ8QFKBehHvobGZF7xL29xbL
tHmmz518ktLm0JlIWaD2YM3LgtoLtavVclVBnuL/glOwshs9U8uIorb86lyBKY2Yn3N82nzIagTu
RC1A8dFwix7paaiexHeErbPbol55wE9i30FUSD5i9PNC4CjfBlpu4jHOwvi6ZF32rPgjSR2Of155
fMIwl/9+oy9YcL+oxhH22D1XsdZ3AI9l53EFE6P19RtKlHlbwtYz4N0wD8melKmWaiEgFkOuv3lg
M9LPGxGSRHdkzo9QdMu/h6kWxutE9xqkiWkQMmvnqUD5kUPdbdK7m74t3EFjp23e3rZD9gzKfHkq
Mq1uPNIUa3I5LtanwKX0JPxVF65yfsfRc5TrszJZceFCFoT3q7Cc1ma+AJwsXwWQJGTejlVmE+nK
TGbxVTsbcjSC1p0pM1IiNB8xe+6nwr5I/IKvSx+/QSaT9RpA+DlwtMhgmyUCpSozlcHcCUNzaF87
dYuUPdvxXrMCgjK6CguxNuRnQtxj6tseAlpl1ugT79CqNTTyjTlbEZcSFBmjKnj6M3Rts/dgFBcX
571/yuFa53hs1Wthph6LUqi2krskGcG2Bi7UBR3I0mehTFWcxuqbJ7COdwlh5y1Aee42/6EZh/Ii
KdmfiZFMjmzEvP3xf2s2fK76mNvXzFo5MytCybNTTCtj+wZhB1PKQVA/2kbiWC0LF/+S0LjNmrs4
02rN3CByqfzAyDYzqOA42+ydQFR9uJbuLUxeIAYXyo3mdaGQowpX4ttoubSZ+ZDuHoO+JPfAO2yG
II9FsFiq5myG7e85mbjZiUyj99LfcVT8K9iCRLzeeiH07Zk7nDfoeKqtO35QqkhQvbY2zI2J0xMh
wwKAwaYPRCBwYokd/HHSxXhsRk4f7V73KZdRWgb2sjZN4jscms+0Q8r1hiTrSj9rXsEIaBEoAPJr
Ssd5duhOvBlt9ae9OKvQAjOX1lvIiMYzdTy90sfED9EogeD0GeXyViESg6BhvO09jDB6XbEeg3De
DBHb39swM6vVzuAH0AiOAEEWVXmOmNSOzQhZ2EdNvVRnx5nDbscc4SERwLRYHtGgTKwtfNdf32xP
cxS8BgmYTcjNjTRg/HbU6ENreYXUGS70PwtZWEiNQMBXZr4P8WgqIg/9XcYJAbZmRycG9nbPiq9e
qbqv90FhiAXfzQo9NS/FfSXDlsUtfjlwy9CGgpuYRPybiTU+N14EdkWgZuJfuZn+XijiK9+9+Arf
1qrOPW/Qvbo/UXHnbrtd5yvUyMGwd4U8S72rIM6IUJjAho169olQS/NDDuEH/wXDTR0mlHfJD9py
4Ke9wynBZTBMbIpolvEqZeS5zOIL+yXZ4xE7hlsco0Lwys8JChcAvGTMqOshBTeLlE45x3Z7HLLv
CTgf1vi1XWhdrCdzFdnj0wOlZSc5NCn+aZMgB/W6xRN5ydrYfH2KLwTJk6XOTiAXIW/IoP/Op9wg
AIEKwXhdZuXbBvhhjKgDeavMzN9e4MaZ6fHHDQRDWEhSOClHlLAMijKkP/w4o1vJnewiv9+Rbiw7
GzS3EdityId5UNqZ1U7oAPSmcpiDFtFqUlqLp8Qurliy6O1fr4+JSh2qJhZId3Wxn7WmBOYGrBwF
wlPuUun3KlDm/GTtyazTBBVZQROdZN15CdRhO2Eo8vxG0pGLAfsbJLwnyLtXVi0BfpcqwHQ72TJZ
J21u59sU1mNZyjxxuetCmGTYgYjIiOe7BNR93v5utvGd9zNrYAS7rnA1j+3ptjai/dooAYOk27nm
tX5Ro13CrltNDRG7veAVAATfiQThZthiYeJo5RRonY/lcWtQGyORZBswaEPEiKO/HJB9ZWMqLl3t
FqD2pU38Inqurcr1OiSC/t1a3CwBRh1n9/Zmtk+lWAAbIiCreKhDdR3y6CKRhiVgfuePhc15sJMT
QGGJ3yGEowGP5uTV5xmu5z89hXYJsVXJLKBhUi4UjbKdfkmxsNLseDIMA0qnNe17SiuxH3ABN3fc
+2zhZCK3chz+ku8HxN4+s8qW8JxW5Ip4B7YR4tCcB4Nh4X0Wvp+ef5w9307VQ9DrlCbjHzQchwkQ
YhpDNZM0+jgee8tOsINZX0+wXvbRFaWAURqpX4TpZ8qym62vU682N6BdebKtc+2fIQcsSbwSfXrj
tOQEv5EYDUlxR+QEN/Tmppr9CRdVeL0WCXwFNSpngY/amUC5EP8RXy1ONdFwcusJolfV/G2Rp/Vh
ZYrFwFT0kULNrLTcnOsSbTMxXJFQwvnr3Rc+7Y1M+4Va3pbzRwLl9UTlNg6liBSWvgIOwAQFoHuc
R11GPw2MrtZfx9po5hCSzO9a3snUBTnXSn9DbK/pD7ADVbWNZpV7va35iFlf7tnip4kqrSuZLy2d
tjCN692m7oW6sep0xh0oROsdqWmfY9m4sbdblLOW8DidIBlybBEEnRubD76Ya91lwHqwauycwnt/
MdjMginkLcJNG/SyFwObJbbbYp2x7yqu0FL4L2rN/6ZyHAis2RASaBV1plGnTW3khLP+jChzyRon
cLLg61sG+21ZixiZ5KqWzIqQvkaWocI7YQ5G7vzJro9hLH3AziL1Nmg2vKSbAAmOiTy+yhMToKV5
TCqCgU1m5TemZ6ODFPNjLdjctCEft3sU07AMiuLSgrbewxdG/g80jNxrCT2cfEYY29+4fmN7xtR3
8wPPdKPhKJgNhBRYGtxm3P4rlJn6ewErLAO8ZmIDVrz+0wgYtElQ2BXmsGAtyixC9mP8Tf8z7Px0
xhLAiek1hiOu3c361q0ArSqPr+A0JiNCaHwJbjIgMEwq5iqelNHh0Xxj8lkH+icAlhSZAA3giwdc
9dEWvRcF4rfvczy1QxdZiKxzBfcDD0hB8cp0jd46BLglo4LfyBeMe2DHGSoH9Opa+Nf92BPuM47p
jLs+GT6uSoVY3qxXS3OYPwgJcxROE3dGax75XFI+jD75BccLY8KK9Cd4IwzXOY4x90zLfAZ6siJt
CQ0RzekVAdr8cIVgY0Nxl4Qz8UHyB1cUqqYrusczNwdLjZFNlyIUraWdQTYXQ0viSnrJJathJGgI
V4uAxobTotBt8xluG8mdSbuB67YJwq87mtFGeZeMLqVm/8LqvCzCBXtR7BVnlL+4J1wUYhkoJUsr
58FtQQms1jhh4D42urDoQN0YDbnzB53+RLYqobV0viVvgZtP3E/m3RQhKv6xbL3xyXGV/Bnt/afB
jrdHCOaHFyGCNl4/giqYkG2twlfl8oLDtUSKbMtXhCwXnvGnE27bNkn+FZCkc+VaL5nqRwtO5SVW
T9q2GI3kuS51NQuIb+SnEtuQ1Jv2hvD+hCZyZbc9tjfl/6agEKa29vaPfAZqZ6vDOBtDPwmfa28e
5vQLKFVuHNNNiYnsedkLKaKriHh3ywqbTLOBKIkjFF9JNmYmPbLVdXc4bLo5j8te4a7POAUqwTWr
4mX2NP/xqwCoIce7t6us/G5SfrSEtWs1L1/TKnvQJcuZoXcQ4sq1Y5WbChbEhntsE5WvsJWqP+ik
nEqDywDF6+V0uLFwKaNiUgvyayWMRNhg9MfB9OIUB1mOHgd/7iR+p/lVwLhK1uFMRgcEdCLKxwCo
U5dq0wdyYSMRolcikYyy91svLsR5QcHDUPhZ9D9GQOl8lzitt97WGFhCQZNMmXMhrbDEW+HhREoI
1eqdiXBMoXhHvhZv9rjgZ809Q+uRzoNZ9FBUqMBZ8Q2S1OXkE2ANpSVKHG811MXOMOg64N1u4Yf4
kPVEIXb8lHKEuf+1e2zTwvhKc/FZU64J+PHmQx3B8Jfq3NM9XuhqrtbHMZAn0L2Ja3JC1BTSJ0w/
/5rdZlD4sJw926/BxUIdMEBglk0yeMbwqOzjt+iGzKmHr29TahBWZwIpUisj4j+qdzL2BS4uinBs
wi2JQFacktBV9esfnkyVQTfa0oXEAAcUpZW6fVqqr11P5045zzRpvxIMgK7xcphMboWptFgoMgBy
Ul6XjpQAKqykuNfjdzC08225BzMgw0sR57ajm0qaSqFIqM5Gkbj8J1VUvycaL72YptwUrGT4AOnu
1YruOSi8DCl01fcME/+Jyb+AgtaG3a9SIhamnW3ur2lpG64+WYjheEk1j/tumFah7mRL+Bs2OOGX
6xIErmllKQLrsMn+IkU0d87SOUjAICz0kKSwtZW2h2+JYLQGRKX0Z5eFoLPgEbNp/yhps9dJXfbD
Qf4QFHEfkv5oRvakM558ndE4Ql0KrNjxeOoJlR+YGNvdK/134ukoYVQiJyS2ctkByiHZXLyhh0Bz
OBOMcq4As+V87IhwURzJmiJq41L0AeAOB6MZRxXyL6g60P63VEKWJsSsIeQP2HULQvXAzJEusWup
321D/GXr1st9blZBNrAZD1GmmJKhd8THg7XHZNZ1loDw22uyw2WlZatwfbOiMVaKsRRznqXOGrCg
MZ7Bir+fCKQqsvl41XinpOECkiXESOWG49OaQWXHJKzA2hnvyFFMHWOiKuWFrytrnS9JobfZiPsW
bRpQLjRxZbcbzkK0sCbrYhe2JVJhRxTjH8/g3wvhfNdTXO3t+hu8DE0TIh0YEJ6llkvMhGimwdDx
KYzgcdGILzGKg71HMVw78+muNsJAxNyKniPPlEa+HgzimE2nQQciw8u5xY8JxmN5WgLEsLkiqzJd
Udy18EHS5e2Pv3A8NlwHPHGv/mEVDDya9Oz/WdI2ih4JOfymHDSLy/pkE4HzOi35DvWfpfZHOwlo
M/Pcw9Vi5G+faur3TL7q3ckXJM7l6HBeedX8dKsWiyWnJ01Ekoh/Lg1jMhpqsC7BCSbrUJJR4sSe
X/NvDQ/aZyB8LGKrw1Q3b8VZSz2T07rWCx7fvgIh1GvoHSEu2cuTcXNqVdNbGdRs0V3GbrX1zZFF
XfIthmk+qCSL0cUbXJO2vARXO9G+L5AM7KbcSdpYakd4Ox25am7Xs/JyGSgkrSaQ+OAYGa1ZsdDL
YsZ9F1+KwV24ZTtiOK0Jugau6gTfpFQUy1FdLZxYyVaX115xHrKMSz2HPnoVyyanlLm4kPCqwCuU
Lhs4N4+PZfaW9oa5OLbKNJwLj7clrhJsoc4V4NmGP7BRb/i9aIOYHyR+kPzzmyxMkPqpXpJM16Ft
G9ncQ2xDvUs9SKgCT9gNTXNxfad1Ybr7C5/m23M9pLlJsA8rm3aihnuNiW0H2PnC3MFIYHZUKcGB
5Mcx8CB8Xez8YFZov+yjeOTONLKkAvDHBRcoD9lUDOlO/vV7AAWqR34l58wBM4bDEZiFA9cKIIhg
eJjFN++l4hxTYw/JD4Ftukit2kkUGMvXeuEIpPwhTm67trjc6qNDPUNoS24dvG1P11pkI9zQLgdd
ZI9KultwyxbNGGYBBxNwm+CLka17siw2/BlWJU5RWQbKV0Qr/v807twMS8OEZtZW0ZUrFOqvKLfL
VdBqtgGcDdn5K03hNLh94MiOQtjTHUA3sTxWpkmeTvmZNNJihvA4vncOfxfCk7At09rRqT+cvTz4
yhq/iUCwts1RqRPDhr1QnA+QjoQFx6V1DMHQ0Y6h+6FZQoiCcbmYL3iT/OjYYXazmicA04nmBfgh
CbHeHS0MxO0LreZW9jkaC6rpjPElcbRoqNaxKkCEsUBDCrSyOfjZXo0MH7uzK4JFSmZuLbR8p+if
dHf45FUMBdQgP8fzRo3bL1SH7EPG9GOjWTr7c7ZhyIXiYMemXusSfB9prFZrBT1rvyWjVjdmMVuQ
VR/axwAONe1d6VofWEgDtLWlp8Tj2xjahVOtTTMgnvqxmsnyeVVVS2TTlxf3eMuLA/N1sEWMfdR5
AUYXVX7FmaJrWtVaQhiMz3kS4q+TgXqrr9bJ9MTWRI5k8508hy/MqcpWkHOKJteHyJvqTf7mJ4HC
DYBJLn4ot0kRY1JU880gE7AUxFoBkhzAj+qs8cpK1rr5HCsi5Hw3tY7v9lESB++4PFJqUj9OZ/mQ
iy2sZw1ACjTRhXJnectypby/4CM0HnYhADltwIt5eEIaOsIwpVTPyvTNEt5H3VnwvRylna8lI8wh
vegpGDcyv6g9VbaGQWkGGWucHG43+oy7pNr0jhTD1+R7R68S7UiQI1VeCTdfFKk50ljJKXqMlfKe
Ak+xRziQ65S4TfPc3zj9j7xlToZVWeAByZAcXi5pRGJmLvIl6dAKyx96raXpmjJWSDZPOCvbiaph
YqQr1Q97tZuPl4cQQPS7LPp+7LmoxBBs4fxShNhRU/OUB1/6bZbAC92kDd1CHt+vWA6sWhiJYN3B
vbpykrWjoP4fXJjpC5OcQ0a7N3/+rW36KJG8740r9b+Tg/1xXv5iuAkzojD8uzDZb/JUE7DmcFmQ
REWGLiPxLcWGITNK1bb4Py38F/mUEybsIzi629f6nOYQ91dKU8ez9sczfz30yskSVQLAr5zflET4
aKv4sM87YD8gpdPN9d6Ri+1fZ3As4qrHwytkrvtGNxQAGoTVckEWKwzZzHG3NwtMP4a/DBVRFrdf
lli/Alj7BdUpeM8kgQL1gsQOkxMQfUWtOLoEokj09eXbIlJWyJRda4cgHZav48ejLKpwUdk+3Zkq
Bw4qUzyQcmbtyXa2JR1Hh3TfCEhZSP2AAPI4xX2itK7x0JdB6qH8pEOViaFXE66Qr5KokrCWZ8HB
ewV8QjEsHULOrsBx0Gy1LeYDhbGI6SoZe3Ctc91Co78TgnaiCWRuWH4lx55rMFKwqgc977bNfgpD
qtonIirGeZyXKi8YOv91bsmzRtK+uBHZsTrJLrlFQQrJE+5csPDpL2/U/qk7JVCs7q3ij4dUyhtH
gMQxjzvaEot56KCFocfPzk5VFhoxrUnW2rHeYbv0A+7sPhCTLQOKOkHYrSYtp/kI6LM+C9J6hYHJ
gqlkQYyjXZWeK5kcGcaiYbdxXj+ub+oHpDrBD6hL+KNzj9A7sUHmFYIMlC01j/03pniIIF7Nn8xY
cJvnDqejzIjEURVWT6fIXt7L449q+8uOVMNmpX5CbVN04g6F3Qpt1esBel2BWaLy53rK49eXKAg2
iv/3TVoeA1bz4E210Z3T8YY0hna8kZQixYITWMD6q94rFwXOqcK3CDCUPnaotDjODH9IELkqYeD1
kNc7NHqL+IlEYL5BGoyfPrVzxjGas5Q3IjQzg4Wj8T+SEFa1c8MADwCbEuGvp7VzVRQRfWJzDRjW
JrgQPAQv/19wXvqn1ewUFSm8sxmdGBLyxzy6YsKR2QThnAOdotNMkid61lNvjisEJGd0qSDyPEcD
9SBVtfbAWEKQPvKZ2qGnIDL072crA3Pm/GBDT7x6En1Rph+v15vx4hsHz+oOwC3Q9fZeurkxL8LL
BKm0zSoXie6pOV+EZiloB0U8+haC7U/C8EoG0h7wqvAAuIMu1Td/xWOS2O/ZrrpUc2Y1SV9uKAya
L1h7DwoK8UeiWIeQwPzvD/UUAl5yTpdhK/fDpiZhFmN3Ad4VsvalCIuMHaPax6MATApNYpGaRohd
3mPlPnzg+nWkp1BlUDju7tFhPWTWtmsTnFN7+k8zaNtyqNtwtIdAOjchBvy0N1dMWk3O4w0/fRPG
o4nO/LBM3Uy0fY8rGZNuIak4+1UIYklhUHpV2135uJ7mbOjrQ1DFgl0v1S27QWSWqSTNQ8mYmOkj
BEJIJMG+wl+Xf0b/CPcG2UicnA9SYaPTRbIC/APUOUOhAY30ARzj1lGPB4aCATSQeY2ugoXTKZ/T
Jkon9CeeCDZOXn2XQkl4Ie9BtZdhuYG1Jmnxd4sDHcS2Pvo5X6yhnZzCijq+neiYXORL3eP/gzDO
nIpIZIw2+tJaOlv9EA9QxE7agdztxizjYW+5xkUTV1UJ6G2bqEaTA+xiYvu7hvqm+Rnz1z6rDqc5
ExDb8d4A6jo/36UCJ+sSMyTaDDwVtzfynJJsNjlBc83PFY3T/9QoiiPogU42WxDsLqTAyg87fTML
CwBf/0Xr5fYVJzGSqnNw2jk29CJbVkI5dKEFJFkM4AI87AzcOsJMxdxhc/AIe/sFf0N812g1hMbV
uAi3STeT3TG5PftmUHjjmjV/1MaZmEqjU7qBtrkwVBC7BuKedmnE3dzit4zRNUr754aYc1lcWuO/
Ft5dPWVV17fH2TWC00pGxzf2zNXjTQXMYRZhu/V7OJpBuVOxrn7htEbKazXyZLXgcRFycaw4iaPg
VJr50e5AKT9jIuqbJIfyBm0AVQ3OgIyujKIjCbfC2HMJE+PV/Rcto4HRf1vIYYHweu27IFOnpHE4
WE7VnuKdHtMciKdXwyly652lCmHk2HIG8lxAxRvn7fxx935ck6XA803FYQQDObAmlu4nV60loZk2
BSW+v0MRQ1qPcCpWYk748qlAepWf6bG/91GdigIwDZZaZjZhJJ6rVhKFg4fSz8gjyuHbNiPdcp85
XCQYVvVqJc768qhhiGF1gbDAbvHVZXJSYnvNmded1OyekFE2NraLYQpErjBRKcK+hyO4dK1ALAF0
SJGyvpf70Nh9Srcd0JIc4vJSzKxNGx4ROij/NjXIYIUme8V/nzoY5rJ2SBr7NyfLqEjoGHSRciUV
qhT4IdCYthHsvZsXX84svlG6UTTD776I9tpfaQjI+ScT0tHc/tEKjcY4a0pN0kbgdevXGJGTZtLO
oyTlBJMjL2C/4pWtQ4t5yt2iAIfJc2TjubrdQpc2PwaLhCrA/G/4lKGtKQjISE+PjNqOPisvV8x7
SUczkqOxb/8y9CcYyepG8FCLQvr2KcbyLcW+GriL3MILoc87LAUkV6HOdvvLe7U/wkdbucrPfLcR
OwTQ4IQI4AsL65VcyY1HiGIlY1QeQV+Kr1BOvpUpP6MFyXKpVi5DFMMB/c6XZLQaIUD5JdABKCYi
Wr7gaUZYKMwq1cppZxFiNjqiu3YrYdzBDKkctoM6tUIyGReeooTHo1V+srKMo9EpkYw8gdLcMuJ1
OTiwmVr3pcX58Zxry9f4CFqkYBnLjTGk3TbsZoAqyXYR1uh1e2MTrYJ4nNJ1E/bYu77rZ7BZXhkZ
jKLUJo5Jkir3a8dwH+eZHy0/gdy3qPAelfaBX1g4JMezZ7CwL5Xee60FnPseUMHMo3vsf/e7ZBCH
h/Yj2P+DkTvBbjLaY+DC1GZ43/pxmCg5MqMt1rM0Jns+C0ovPDI+OrM+vYr4XhB5D2An3Tp6E8qY
Rt01T7SPR6B/Y2ruysAow1SwoPOcxG34ZAX+/qcKaUYkWbPW+h40ULwzR/o1ZpQhSniQmgcuiS0J
8SgFvNxT1DSnjXAu3OgjL5cUlDJQdSXIWEdQ1KbE25nvTdPKu60YrfQArGF+rD6lJgjcBfS5GDPV
nHPe5Kef6DfIwgybnxBntXC0tCl8uk9yHUYkHTqetIAO+xf9C4yLqmgo9jzp/Hg1VtFZIabfavqF
ILT+bRJdwSHmDK2KvXYgrTueMCz0gHxg03+KO8LvYhHYKOIQzg0gimgCGe7aewDJrg92Foa4PfaV
RuuGaleN3P94B33awzCJh/3hLW50doq4H0ngNIgHK4DzAwULQjNp5F5f0Eatu4SalCslVlotvg+n
+rqF3VVyiLjENvwdpRUBrpVpu82ksRo6m+AWwRth4jwZruWP+sCQKCtgSIQD1T9E93T2n3gLjm93
s2wEduvmV9XnTqdiJMwVv8vafdZpk5vn5X4u20ty0huGhX+HOEoF45IsOU0LP2VfOe6+hxBkYajC
CzugNC/ccCqhA5nggryg+xKN+lRY+CPoTZNTwm+9uPm3zLWZmHxujn3Xr3ry6s62+iI07bfQ8JnY
KtGg4FY7gl6TdggZPUdZKg0gLzW61lZy+qgfjcZCON6BVVvDFtm9gRl92zaX+c8mHJ3Y/1CHxpwp
Z+bRtDI3mZsJdqY0AgwlusmrQuK0rM5MTqSjWc/6/7MUko7tLE01GuX5HSV9Gqq9Q3TYjq7AceT8
Jlo1X8PnCcUuqTm3CdZY7huJ5Qhbvnw5cLECFsGrQRELN/zc90hLlcx4MjmXBWO2xrucKeL5LCMc
1UvrLS3hBvQ2Hdf11BauQy5ZnsKDCTJzX9lrVMQeakIrJintUSDnFsrxfxhdy855fxwnP/FktfhZ
2qxTff5pN2JpUxauENtUeZMXf6wSbjb+fWNN1vTmVzbAfc30UiDYVsND6IS+DcI7cmZFRYbPE9vz
xP1TrVIcPUfr+Tyhx2xC5E5vRi+9wjB1WngAWcCK2kwD8IBBKjDzn5ROvazwayXLQbRwomT33xSm
qcxxK5gLkGCyKlCnyf+xo7njg6kDp67Zwc/QULwih+o/LvJCMUgIkKIhf9sIUFcBqrUeuUegOULe
LPSWZLNpCXsT45JhPeLXkPYmpbNU+tg1Pt0x/Iqaf6xmqp4NUWJ+b4RGwz+DwvvAapmf61Rib/ef
kCite2iI4mrwls7SkAbjdUDd0n0XbCKKQyD/FYMCdkredIMVRP1uhIA8IU6iyPt1b9qXoHBGfcWJ
wyKHdoq0Cv2D1v4DbJ9qLa/AAshaNtjdxpuNntAwnYR8s0LU+qR/EKnePObQ2iTxDKuhO6Mbbatg
Aopx9jeSwA/ezRFb8ScT05DzfErAQw0J6kld2UadqH+SX4xPcD0jHtagm7IJIbY2tj9C79IQojEd
292Unx5DYtTcQVLv5UZBDS1g759lbVESEJNaNq7DceZE/08um4onyH4XYGHACApKqK6giN8Txduj
Yec8DwD4s/mtW2IlbIRaRk+sT93cpywb5AXbyl0ghBBkMbxD/B52CBy1WlB+uOIdl/advKfSfLuI
LvrjghYBGRWQp42oHd2lRCmkF5VHm6H6Bq1S2pbYLKZOnZ+8BJoBcNcVr0Ubg9BNby8yMCEzDFB+
GP73m+/Jg5DaQd8sEADwQyJTwLgqsNveffkztyYBeMfzf1H7+3Ui1kk7YR0/WGJ91PMPYuZUC3TK
bz32uqVhKgTR5praeIzFMy0EffA+/is+TuGkhPkGba69/yQjPVd2/KMJMHvjkrS8+wrs0Og6AbgX
5+W28Qn9pVuYJkk/B4ZOlNZk6lF/OfNOw7rEUhG8bM1qyLeKiF245tBqSXtxGmmQzAUG/UOPO7Wo
QezqAnIWLHjNNb8C20ohV9i1TUeKccZwv6xYZqZjIzcpGRWIYeS7qBQo+7lpeVN+RZejm2OetV8Q
0etUXZIp9rIv9czqsetXqze0IboKUZJS7tMxsK92+ChZDM5Z48vogvBqc8ufUWOZFAJ0k6diZx9U
Ocin/niTFXVNoUEkVx/icFbt5Du1jdB3t3MG6I//+S0or5jBvYlOJ5m/U7GhZpaNoZkBP+JNP9xv
kku5cVdYcREO8BVQ28xpQbOvLcxSAvUodMi4cUAp1/h91vcdga4miJCR43SGOBWTLDCAI2KVGF/C
zdpItPe4DfMLXjRisLS8Pti5XG1gWNyzRn0N2jWScFaRmulnPlQp1wp6g/vB9ony7yEYVh26+Kbf
MfVzGUqrCMsajWuiV6jScfqvbtwMhGMHAaPG3YJjJtIdxMFDXszDkJZrw/N8UtP5ymXrY3CVU5sp
M4TyInnluPBds6QcUZC1/F2KBf4K2diMwGDnLMyHgEC9AZFVJUt3nNPgNy+12KurtN0y8CF6K3Pe
yk3AHS03v67oHz9KtcBRaIEzdjPV9EHEGb02zs6g8nvASDWRjRg556t22/sI9zdp42NLOlUY6hQJ
kHs3WhKWSy7m/bHztc1wQp0zT6tndExNf8TOHPNLcD4czHwA92Uwb7pvdV+4oeirxowmhhG6PiZn
QgbZcc2p+iIddqUtRe5QFF1YFXiBXIE8UdbZP33hUNoxwvCy2n2kqfWjU/CcE79HnGQVb9IkfWKs
HwbMu7EdVj3cgVvTe9UOfNLwC7YOQIiBApNQzrNJfV69IcJfTHx1g7J18NAn5Xp/qAFxKwiL7Ggy
fm+Wp6jYaYUTo7rLblcYpuVz4ykVHAAr09uKAtLZH8QCC8efp9ekZJ2JeIhvFzV2zyth+QMN19rU
JHVAVUUxg70+2AfPzScA92oopZos8OnlIGbGwE5XyHwKL3220NDx2Juvv8h01qogptIChXbz04rC
m1GywzkLJme+d5b8i8Fi9SMerHQG7cJK68mvoPhBB7WsVfBzJxqZ+4iuXv8aN9OvIouYHom7x/aD
niVMDw1xpSWEeANeUOmAlj9C5kfPuINwFFGgI7F9TiHUhXj9xNrNt+XgxGZblCR1HAuvW4mswlu6
chHGv0f3e7l5Xl43JZccYUSUeFrHCAyeqxNQDiak8HS36DMJjWBi3Zap4/q5XsZjYfSATh7YyKNK
A2TxNOBunVdyWoH2V4iMXpUZYPWWjWkePgN0PsOwrySiIfzIF/EF8crQfDzzvZTz7z3ClN49EWat
nmO1sLedVICI4ysMKzzjDJuEjcGmmP/IzEgVdJURlkwDMxSba/GjJgjCjoNnz2NMm45QwzLJ2YCH
ITmnRJSFf3FnvKRLgr8SZspEhbot816068pmv0hlckpn1dfJ+FmLR75n3H/0Q5knj3n8ZpSGErEv
3cDs8f34rSo/nY/gwVc0C0FxCo234UtdTZ/PqmeeEgSKkbhquXgxRPXkwNJZttCx0IWP5ZzZ4PsG
5e1fpz3Mkgxk5awLYv2ot19jxCpwUidxVwcilHLwrJNlUoAEFlPxP8YolWcKvyPOMBoraiamAJMH
y6XiL8Si4BbCjgB2x8c7m5b1Vcrvm881J9pHqd71D6vQEKawYsyJ0wLdzP3CPhQSvKxG0/MCyCbz
xclB90j6OdndbZkCww9J7SWGLBOMfwcUAgKDQQ37u9eOvfTpjK1BRZ6QJu6gbK+bJa0niEXzSgcf
LTKeLmvQ3WcUMGwfclqVaGC2NiCcgTthb5b6KFJJkte6BZn/kMa5n6Z3mjHK9G1wAmBj+S+bSoRl
kdsjJ2J1mkb5e+pB2xHP/o+Id/eZvZj+Di4wjvAYvxPoDgZbt7T8i8D/y55PE6cE5MHrSNPIy/an
KYuW6u/onBzKJFNN9H+F9mUJriUrpwKDw93M3dAP9U/IjF+SGIhGJvWmmafXZe9iA0SNmtIItlmo
HrruwBtRwBkg2xrZB+DuPg8HJCkTgiPCnkjLY/mIy1zwoMmMcWUqF0CQ2WULkGSJQmpI0rpPb5eh
/RO+J01GR95gDlNPdvb1KkUzxKyjE2YF9SVnsVWizE6UcXbIitZLyGnuPmgk4Gy+DW8xV39BWaT6
en8kLilvfKr+F4TLlc6fqzhY0ujfNpQHLCqVp6b6D05NWKzZP0PFe4SlqBlap/FU7I+gq8B8A1bI
UmqYlgNDz7zNt3x8HL8OmVu85kTXdp68chPh3VVl5f8cbonoKW5vSH9yX4+NQW9Edvq0NvdIqsq2
pFsYsJ086VCvdsdJAVhanIEcO4U61uDvjb33ytvsveLezZQQ1UmNyrDXDeJDZrzG6jn/sv2QQQg7
zH5NXs28Ip/tYHsjXZSbkBvQCWjI4PpwpgxqdoydJmCQ5hpNL0h36wgptCNdyG5hRh47WysIiC9C
w1uzkYmM6PWhLWlpgKda0gxQ/1lp0b6Ffz/0LFwy6DvgMriCpifIjuYZ4Q7eKNp7m30ULEUahhrZ
x2FfprcOCrCM6ca/DjnevwqWW2UgssskadWZETADMvci86gTcAZNmdt1uBYY6XyR3IsPqyqkvzgx
ZgFhsY8GiNX5QetEq+JhMhSQDnXyrAvR0wBiOF/vVFxS7QkKXBHB/rwYDi/wnYOJENVWqJWJw9LN
M2YBUHMY3SQl6nZbGWGbEYSmC1RVPphMFp6vzy5Nmk60KsT6SJq7TuBhQr7spGhcpgMW2jqIsbXq
fEXXOw1XbbQjKDCNoee7A+nOF6KYr+4A6nlsqreU4/fMWj5UQ9Q4ipScOGGaXfEdqkmOwjxVHh94
7SQsR3IULKFrdktKBAWAhx3Dxc3CicmisitPmO1nWL8/5fFULCRPsLsjahTQEEW1DTE7euYXaiIO
ASawodCT3mxanaW2UynFlbU0Jkq9Qpb2VpqcSQDZ3o5wAtM15lwCjBcytYDvBX2LH9MplNPLGaoq
eXV7qnDsGev1jaEW594Jb+PkHxLdXD7TNlkzuN0mJnw8HF8vyk7GflmdbIpKuLzHDJMcEE4VrIi+
Bi8D29h9exUtf6bX8r90KmtcIspBXOtm9uPjOMpPC/UsPoo6nqGg7VaIjL4EYz2tu411x00tXpd+
DdDNHPVWVuzDunUjx8w0wFn57n3XgSQqiaUKSEpdM8ox374692qCIHqsn1MyEPupSgEkHAAs3s2d
xwYCOGNNeKrtpJKNIP0tlfPpH3dy6EFbtGyP6M8XgwnxN7PJqQgMIQ6gRZ1d77J9Bziv30Wl7oMG
iYFGrx07xDbl4Q9bZGiy7pmgK+GbEuR/Unsc2rUhRseS+0NnQQ7rwQpr/ndjAri6mglpJA49QarJ
G0bulil2YiK39thaKeJuKIAZ2uA5PX/XIIzjLh0kxOEAlpUsKcDxcD0an/niuR0W6jNXT8EdoEKS
Om3WzdFE+K4nslxStD/dNz5nA7KaG9CuJUqmH8aajotN2+1PAhAFVOO+q8LKv+0bTu5uN4WEiUj3
Sw4+r+/KGSzkX+Pzi9VrZrganzVpZVau2h+oDvvne/Tz0wpYoGApYmnM71LkBktrIpMQKxiw+GF8
89uZT+cSg7fDnsiLmVFeABVanu63aGN2xDJiI56kamCwM4Jfy5NCgCfRrWJuav9jUJzLHxVRBclZ
OHU+mZtXH9FWcW7yidj4HJoel4B0PF1qus1n0wdhulY9+ybPSs/yqjkv4NtSpo2LnPnCAV6jbIjj
bj0BMeOTxR8LYfg+JLpmQKOrTFzGLuyygaRhwYlHkqQ8uhWUtsjf9M7t/gjIEexzcXXOZ9AeJ0bN
wdaxb+W/V3AXZHOT2iknByily+H3sv3HvTODkqpqziDgVccexEB7Ro2Boe7d3/pDZyv8munkbg5M
tRhxR7uDyvzo1FrSe+qa0goxh/xB/TxoPAWK+j8DCa/8iCa2QvCb+MFM7JoN2VWkz9+rZNVCLqBi
JrvEqJW2mhYfdAwxTsemMo8tR8daLyIpPrXyq1oQcBxZ2iB01S370lTIhH9zNMbGdACORucR5sv9
8EeYAdxZPBqH8t1gwtO1c1zpCP2mpm2t6ZJ5+AbCtb20AQZpkZGO0wY6Wy5fcogzvkqRC2isSEQ5
h4hnIOR2Mv9dE/QhJU/2EO3MfHZ9AZnbUXGqQqzjgi8P1fcJNJhIqaeiJ0wWCNu8QyRWmHhuFOKW
kSL/8hle4XcbHcNvOBL8RXmeK0i2xtvEv7E4Gd5ezUS3tqdrQ6uyIwGBIZGPDENAvwgoxdIK/DKz
l1N2VamxCNgAYDfAQXV66jxMPobQzG8fGpsDPvE0JofHkSBZIUb3TrLHKmHrPJ1qAoyILG0adPem
Z1wsMpawKESmKa32qIucSK8p2yphiNPkGnzZlDCzbB0WjK5gCMrEJGBnmma3jZpFsw6NRTkytFLe
0rYG5FunxgYszJQFe2OkWpLPG/TwaKYsVtUPTRkA4dKTrXB5U3Cto9pdwWNRg2AvzXA8pz0c8Jrm
5L/78kDga0xUnNjroEybDNx5idyAZDb7PjHiYHxIy9Ufo+bRbO9+b9xrPtIZOlOQXtc1QEK5cywC
ZO3PMJJRARLhVmLqi6/FVhUr+QXhglY59IdJ6BkadfOKL4VTxWRL9NFpNV7fg4zf6mj9wXa/0sYI
iIFLVWIU0tfwreIb6rs+cuEtbR7rWgSJUUeoDrdFBg+ggAnhP4zzaE4K1hCpOqGr/aMgAjnLalGN
CY8M245ZO3B3zfkbz8P8dipCbS4ToK1PN8BejNIMryo3otimqeAQYvz76YqfoZvx5EPz9wtpFrsF
8Bj1laF552QgQclxoruw6Prgt1C/yq1F8H8Nrv5sxLqK2en61K6XSAY9BF3GlkFgqks6h3tKWEcb
myyKYh9JeHGnHUKTw1eaisopczjxhRLFxlvkShDxHB0QtoDc22o3snExnejcmBoUwyY7N4DbxPw/
5pUC9oUYsQGkhsMoxYrR1eAIgP6q3q/btW3v7vdMRw3URkQlkyTE3x27k4TH8JgsU2+biRnqimiz
SCj+O4HY10JZufiDnXR49xtzpuV8rcCgF3rJ219ZHwXtiFS5uGjx65rVpZ2K5rGAlrsJgCNArfvo
tN6kN/8gUctU7qViaWUsN4DSvAMf7+8Kp5n0cwXNkfPhPk8JdE04/xB5BZ/9kuQvxqEoGVGMA2HA
b8zFmDkE+xVXqAfTb7+ezwxT4OYGaYrFdKxnfFgfo+3J07YziTerMuJcyWMSgxd2hcPpr473oGoD
4acCyfKTEPF88ABHS/4JlXZezMU+wu6gCdU+8BRxW7tSTeKsMqma+XG3ZZOp2jNVxyYzwKVnGZA/
2mKg7Otk3T34pWuGNZiK/ZsTs+yaN/C93jdhUxP6BuCXA69Gbk4M10FRzhkbmTSAYvFnLBAG2xJk
mJeTjK2yWyC7iAi/xEIQJ5X7XSZyDyFiSSnwA9jjl4xs0Xix5BQWMjLL3OWTBplAv/Xnxem1rc1d
l9yD3PteqMEBLPCp+06owbWPDiNTwiK7vv6P7tr63TttM0Y6pwfU12h3/u7Z+GtE7EEUFXRbiKtD
ZBxYnwrjQoYmXIvD9HC1A2SIAXaoGMkE2Pgws2kHPR/+F8/pYP5OuzcLHZAl2xMPtV9PU3bRM4Xi
HMO/wFhQ3aUBj6Ox9cfjGR9F4GxwkrwZJlsQY05OxP6yNQIZVHmLPrjgZ0TTNYvOweJQ6VCFXH8q
YYV8aPCX4Z8BBzpwDH54rg/pchFTyB+fNT7cie+vQgJQNfRtDBQVIWvTRF6sXG9cvlppa4et6qHt
33XZ75+hJ2CHQ2nJ9BGM/3YEEwIdVK4pkytiq1AlcOS75TUl0esNUGuGMIIX4yu7c9e3yY8vsA3w
TC7+tMMOfgTL2SlMwF2GY+9gnBiERnilsFm4yVpyx4ShA2OaiMp2wQliaJdx22K97a6STP+P+5bn
+miM7AZcP6pP8VUZYtQQJ7gEXLeDkFX4m9vtzz4xNFkRuGcBSRFiDwKDamxXU2oLvBUAWfuHIS2B
G/MdU9BQxVCG37NkulmCG1it0UL+V02tutNa1knfLXOLgAtYVbkQbX16sgn3zWVsrPHdyVf15guQ
G9YzjN/AhUqNtqnClBi9L6vZgItxZtYchrn2/Azz340kX4MuHWE9q9uxCcxnEBRiro+SW977BQSP
51vXWrvOtGrgzlN+olxDlKvkOjEICdK56P/h6mjsEAMMu0D8KmoDnCZEcwIbGABIrFfgRwywRNFJ
vZ46skUN36muCggN/hFmOtveObL23vJAOXXM3Dzv1jcGcZc0GRKE4JuldFAJX7FVWyxkFMYUI3RN
SqtgaCvTRqRVLmvtged4CmZRO9YGPao8eQzvbmMChrYxx0zS8bpVRILTapSxWyiXgDKnIgSEGWxo
6XxDtgGXyHnpg3m6+Ve8maI/Su7n5LjIdqCennxuVHqL6D/0Wcg/A6WuwqOrAHeRBZ2XagjwXfXI
IycQpNb7kc8P6h7vYVUtPXWoelLGYsUz3Xk3TSFnTb/XL5pIXl9yuzV9087fjv5qKieyregfUzjr
EZQhZbvhtoi/+b8kV0BXg8Kzpb351neQBp2AwdZgrwBtONlE/vkyYX6GleA2wSaESVkOTjFd/fqt
Z1IsqIzWtXGjh1KsPIKcLjXFd3R7FbguRR0lrV0FiWqQUvcrn8TdQ+Iwl8r+0HkWWj1IvtFWA+87
8CYER7kihJmjkBDPhb7Dn6jPivlH6/4rxfIbXhc53Zyb/z79dC9i576qsJbtQD2QzYtzB7PQf+P8
W4BlC1nARg00IkFEWicyZMjv/yLJtrbST9OikuaLwHKGRRamvqn6bShPaIJJeFFqS2pJBRbzK/Wu
fbp/+0fseh+klBENq4EfNRYRqboDX9t7oTXjnoMM8IZ1R1mJqpKsvPDwg0QhGWqR4DO5IQHa0N45
O/6rydcYEXY/owVOBxVRbw2I1ay4rNrp0/cz+FuEjuQNMsZ/Ueg3MWMsqoIUYaNVihJ4zFkYme2u
OCAJ1qjNrpJs3sQjcK2ccP5dkIqceWLJj2qmMnKPbETgs4Hcd7J3gCy3/UP2yFH3nD8FarK7h6mR
QeL+6+t8DH/UDxQRRz79JEkW7GePSV2BtDSts/yU237QBQSxT3X0r4eVmXfhNIkjL21Hgq3uvzlD
DrTrJSQSBhP/sm9Y8qBT2XwrYajwXG04lcpC9/t5d0TzXGtVeXoF+FvVQ/MWoK0c87x47pfGvvHX
zzLEIJc4yWEpUy5/sEkJXStbKP2M3rLD0kDRNOxTcDXt7ODGEkbPSrArmXqU4scBvyjQtxh5Wm14
96tXtzcrcmb6A2xMU0f9+5IacAGlQ+FZGYJR+uvad8uoP+VviO+ZPsLUDMSsWE1v2lMRSzJ9DEpB
1yWSjeVoMCdYAadsmb6uN7wcjBFcmcnPidiWEM2GUvBQBt78Ker14eexh/nH8TpnhMjNy+QSXfW/
dNIvSoiCQPDIIgLCg6AIs5vCADAIMP+Cp82Kar383duLAEUSTOYa612WBymfuskZ5V37SLSiewm2
jNuQaAIeF5rEatC8lIIAongl+vcEq2Rotk17phLc8/SLpT236YglriVnOk3eDjLcKS1WCPyRJiFH
LId7uJMaBGdEsFYj5G9eQdfQpETRAJhcgUCBhtLM2z6gzp+XuxbjI6s9h9YD8iwDiYJKJbZAteZs
qZBsxhR40dRB7Wxf3aUFNGHPnLaMpjUd4s/zghr2zLpZ9701A8y9r4CyV1Q/bviF9OBHa9Faww3u
JNFgbeDlfRaEp22now3HZHf8lLlN3WKmjpYRZJNXz6QSZBST+QdZ47ln5cpNEICa3jPRZ51ufmRc
XEACKv+7dS41j796z1ccLgRHOmuJCAr2xZua5ljs18q91RScpuGK1QhvulK9p/a2Hp9chSrF/RJ7
a2EIG7APS171cZsb3X8fo8E0cKAnGd8OijhJdWeAAqfiUx5ecMoumWGTy2x+MMPPNLhXgacmAyRz
KzQehrRfxUfgszpo8ZR9kjWbRrqFksqgA04/B4q/9QPcrf2DUbHZa4jkyjv4zu3p0kDpS6lsLWQy
0yYP5uTr3GVWCLbvQPzbKdBSMm1U4nUhja2I8N+r/nWQgdO5oGQTAZzkf81yhItVrqruby8DWRVR
d3dTs4NOrsX7imQS6D0p1YV+54Kjzib7hdghajNIVl04fGY7VcdCpkYpTs+wmLwXAel8AoED16Ef
PfqXbemqkSAWDlJ8pfeauJY6R0Lr6owO844eRJLyUOt9seorCPo+tghxzFpPPNyCj43a2F2UbBqj
UTbHgaQ8oSwHrL1RMuFV5t6yyVhTVuo8ab7iJxESeHdL7IcYscplRdooQmfnj7ZRGDvuW4fhid0R
/5PC6zn7pARPGujQRvqLR7sXCWf1iMGzCKE0UcNrfaTZ6IwPeLdHaDDZ5I7e5SuQ2OSp4J4zcMOE
blMXV8ESKenHu++LwSc1zkpXHLvq536Hg4lSjejSeJFUT2QbKMH8VuSCreSOKOXz5RMGfWXh0lUt
qJUdBfSKYs5tWnf7TIUeRizSPf2ntnk5xYgmWW6lMBhNi73epGvCnd7E7G22rRUJrNpHTDonSEn9
mStOPlujq3xTlrFZ2M3djmLd9PQ/W/1hrFgBYNbtcQJB8DSmb3IPROfzs0tjrGlstVs+mpqfxjic
F32Znmp3aJ3bf6Dar18UFmaI8DbRhuCm2PCZ8HdvTHBYOIsDtpUn4LtB7Jt7PnKKwIoHm8YicLdA
2fjHRhwDT4/WSdTOcAEzrqYY/PRcKg4Hc8e6Phck7MacL0KEGlDmMFIQ4qfItG8JTTE9ldhSJ23q
Ozh8EhM6FX9hj5NUkf2Cg7YDZhecDvDVq3PK2l3CmBuh1EYxNe9Oj2AVvJanfsHqbi8Lk6/X2Ku+
W3OE1Ct2Y0BCqd+N1WkmnO+NyfVEwM3vFH8aD809wTwgbzNXdrCfcrdDbbzzZCQX4ysnCL/2FYGb
OVI1xp4GmKFQTitBTIfwVZMZebVSApdXHnJc4wQVSIDLWnYLJ+/yGRo7ck6fWHTvIwb02Ku6Qz+0
17HJlxQONGUy6ZhD5Vy1mAyPkoOYR3rPjsiY9Ow45r+hwhKJcZrbMIOyq2W9VhG12beFFzRb1Qfb
WsBVO+0wmDNkO7Bez1yP6lBwNrjFgazcILwOaE/seZnCt5D+MmYqSyfsWtvJbhZTF+EP6VTUPbaG
2+5WJjTCv64OA//IiJCk1vV9jmTQUWjD37x8A/OQSO11MSjqiyjGU65Nz3OkWryC/J/wiS7qrMBG
vn2CFf7KQ0Nq1z+nYrW+qZ3bm3+y+P+ttxsjiormSjEXc9Jm2Hvg0LL19rb/NCAIgFsdtuNFcXyK
FRu8WISWLRlSQzDtn5SwH3s0FVpqwOCBmyczZ8YzV8KIYpnRSyKWsUd5zQza5JfW6QvE2LenKhF7
wR87e8RY4Kg+X37Sc5Kl+36dI2e03q0bI3NcTa/fdMyhVvshrGvEt0ZhP9DuXYiSnpaYa7BU0xFO
AuMl5P2zGWRzVmX5eQpb3xOha/loWJOFPxg/9YWPY2DRbPdG36JmjvuB4S0jVbEyDsW50jeQ0D+R
ui+uVsEACOY+zKDxM9COEKUzTtlaMdzN1mYSJXqPcFYZx4SVfbnuTf/Y7XV+66iMYzUnLrpA0IeC
I42OnP/HL4dtiJ4hPcQOQoljAzMCwbIeDEMbZEzFbJ7Oqsl4mxXx9mDsQAJJDxXiPKleUEIc/Jk7
sUyheOBaqLBPdK3k0K1mWMAeN5cD1UkAJH2EjGD3WretKBFesOJrR/0Jf+7H4P78Gy1nv1m7KWhJ
RHkaCkUj3hwbGw6gMHo85cV94mqC7La2Fqz6xliVyKNWVGbEby+Ef94NwwZvfXXOVzkgQOBtJHBf
z+00eRkK+w+a6CM6H/rOJC7PSsLs3e/cypg1Tk05B5xyF6TcljHGgZS+8mbES6+cpYE5nTwg+aU3
0v8luwwGIvPnHjLDLpqEvKvl5B/bJfsWUOWCb7k5/cxL6vTJKH1jWcBIsB7JsEkCstJaAoIEhpnM
oOMvvaLYihehrmUv7EZfyKvUjrdOh9Fx6KnMlFmRUH2m8wkrcuaTem5e1d0KyyksHZpmY4ouOYMT
0uzsBqsB82ooOF3eZtw8g9/48tm9NEkp+n3S7x/AIhc+J/9VhekwtrcVN2mbRRAJg4HqwpUdyY8i
feDoGnrgzBVt+nTYFViiJ0+fPjOYthdbmUlB18l42C/A8am6rX+Nb1crIbT8rBr1nJw+Xk7FKnaw
dWfQSYLSYQEwbqe20LimyN5glzH0AuXdDgIHwdXJNltNAYLYURi7pCB3OfVRw6cU269s3fQVjPku
fbgg0sC+zZmn6LzYwF4wO/BInqJx8dC21nAWZ/ukG+mm24rTnKugVlZkFVJ2N8JxajWwSLBf8Uib
Ckis15RZbwPjrUFgBc8D6A8C86Nwz4tg40bzHUBLgnPETA7m/z8WMK0ubvAg6sm7O196KAa2Rjw+
Ss/IdzX0EgngesGEUom/Xi2GOflLYFmHThop9sgRgx91t5bApg4sxo6swYv8gL5em+Do4Ck9G9O/
QptQPeuP8r8AV3muCmIhm45Pa0ArDboF4YswcgIO04AYu1+dVFi1MWvoYnf/KKxh2lSFW343sm2d
hn1tUktjAZoLPyMmxkFro4+z0wrL3b/M95J3lLxCrWqCgix2tw8F9I5va9HJt3ltdXOmjFla4u02
3ZkkcdOHLcELQqUXL9GcmXpD/0NgVVhl8TyGmasMfGrI5n90Gd0+d4VdA2YgBRatlfO9bMppm5+o
WHctX4KSzMsPP+XW3XsmqqG0s+4FDtYbAhNpRDHp8lP8to9xcdpcogocp0bCp4YiVFkE4+lyaf2G
3KBhIdRlvee1VP4auIEcAVP+/suyuvmH2T1lkMbEpUTOTrdFgN+PvAdEtN+JygAjOjgRYK9FErgc
TwRZQGfwx1ObzLrQ7hF4ii3oMRUQCQ+CBGRQhugpIFpFd4sWat26QFOL8PVwkTkwkqFj1x+WaqVy
z8VjkCcWWjJSgpEVxvLXfHUTMkoLyBAtub9HhGcJk5DspCxflw/UMFNqJtCm2vezLcMF3rtOlbuE
QijZZap0ViGXgmu99KXUwsIBuzwJ//Bp+JfyASR+1K1Zvt/vHld6Qb90uLFyEVDVdUgzLxV5XNqb
ZOMtdGp9+77GxM8AaCwRQd55M+QF9YMC1rYHjOSWrdwo/NkaeLmGtCsb3MWaCvdTvNhcu8t+cjy1
44s4nhh5JKLqzMuaQlK1TtGUkL3i1FOvZjJy1Vij40qSK6dCvXrD+7IjXVeR5lgyETOtvIatI65U
TcTh0Jf80af1KN1kTnwXqaRZGNv3WrNCPF3RJzIt78vCK/TqzdOQukuyNBxHhP3go91Q3c61FZ1L
ysHVaItv+9TlUULmLOr8Ld+IAkwkgNwHZtrv0iGzGYK/LUVXy7jopZ0TKsXAdzqvgRCHlL4ykxdL
pNG5qB3Xc2hBFGbia/3WcJIg+//zqpkhAUL52rslI5T9bLN+1jJDp2N+RGrv+Gcv1/8IHpRyPHUn
MkjoWYryRi+zl6KNRJKoOqpHyjARRAIO5v0vqssN0ACtkBYWfRpgm31Wznjt9OqNOCsFhGswrYRU
8POjswjI3JW8hYNFXRPOHXvVaM+fnKVwomgmxQJzxGflynaEARuBFiioTGpjxFMecVLdCCnCioOX
Nj3ofLx0Dc87EWD6/ukjXch0sGWjzNPLmEvM5ad15Ve6JxB2ZF+g9SOb+9++SoxgzTO6hOUh/nRl
yKFmVZhdka3c110m/cZkl/AboPyvVCswZBo7CQ47E/fyuH+dQTeHxbv3uDPk65QY1vLajMZ90QZr
bXBPv+NgvXDY2BOiMQNshndBR6D6nr4VxL8/UeA9GrJZpadEk1IBcynvVvgHZpOpzeSmlEvLoueO
WrlXjwS3f96NsNAKpEZef5AGXrLLBL63/V85s+vJ2h1qN6D3xOFrxq019TdTHHygeyyd01jwPDsm
3i/ZCycJFPEZJeG5eRtfhht8yoVKwGRmI1OhWdiH7/+5WYL8K0bvFbTUPJfVqQe691dNpbx62Z+w
BBoWyHeoKJrFDBLwKDdQdaBh32S/sZYbL9xssPgPrv8ad5PD8N9Z1ATpShp1FMKSJYTPiky+FMEq
1YIoovPlpf3XnP9Z06r9MQsLMGCVBTJ5PM+PqQcblWcWlkrUUxKFiPM3CSmCRQ0IwiR9Mno+LEnp
BrmArwc5FnS97roFWtR+RQyqrv9QqvrZv2/FPbMusNrIXe8nv82yAG7aWlDStlkhWUAsiN1sH8y0
m9UUvLjPzmRw/64gLpb1iwlFHAJDbL0DRGXMsvhQsiveH/JorE8sYjUe9PE9AZ5uBcKac/WvHZOa
1E6sNpBaZya/8alGC6F8Q642+oAW4ZOfA7UGJt+jasN8XAh2pF2w7BW2Vnday3GCVULoiqVEuQpo
GX161ZmEoxMVziShhEMliKcqqsyikReWI4ARuksGORa22tGw6Kd2QHGFwGg2d2dhyjI5N1D+ZUDX
z8lDhaaNOS0RPyASSYhoGR/zvsvt+AIrYmDw81UXIQlgEIc2yRdMZlGyhr4+PS8x+A2GiEf922q6
wJEQVCOQozKH/NEL6b8AKxcZvZCEnbXMCXPEu99wjRBGfqB8NPSFYVNXinH6pkhNWW3NHuikhj67
KSRQMzW2NEa2ue24wy6l8olW9O/gg6BbDxM+OclnKIHBjYQVr9CClVHzGqAyw2tEkezKA8pYLqcU
YBtu/Z29Bl17snxoSoSLczgybwDFtJMZdz4A6eIQ/v7h0kTYvHNrLpZQJ+8CfnhGJaIQ0meGz9ri
Jo4rS2VqIb8joFPT94Lj6p8FwslEr/f0YazFowWPKb+WszVIOM8W6yK2AWYzivK7PnOjTdYIDMkj
Jd8HnUX/N/AJXUIbFGQ8kBTpbdVujzIMkgwgP9rQW6xiIcXMUEpPr8jblNh4CXqkUirYjasBmUgt
3weBMyUPudHriwa0Wy+QZ76imwohtkqZPfinK1qiGxBZNn4pS5UiRvOBj9M0X7UWq/mz/FMri7rT
sKgOdecqO1G/1f57JgZWcOBTEt9SKEXAjrhFiCGfX950xXc2/GMl1FAAcoA1p2JKRi/yI5IoTClI
C0pXdFUk5jJCQyfRtzvLxmrm5rt1KgiENbQebnshoq8DUXbK8/gBMzmUwly5Dt4P+xiKjRVhbSyq
2o/qs3IK+zh9gOY2edNGoVlkhp7m/arZ+q7bNF8i80iK0T669A5Eid0AfQn0hP0OBAmgGu9A7Jjc
19jLv7skVHUd4egk6Rj8baUkMKPR7/K6J+xsvGnvs8bUzhK65tiL/AwRSpW4tCMtm28AQmFX4YyN
YiMqmZYq5soxCs+O4Ea74CzLsQyp854KtlJqttP9fFqwwlr0mAuCOaIPCf61/41w5/rlRGvV+meW
c8GNRK3H42MBPZ38YtjvrZWIJwzV2VfAyg7dEloNL65LTz6QCDBipBvjFtPAHXmnEK1sFZvSAIlq
p41oNZceKfu4ZJatGk41e6aM+6NbSguFVclNHNElj9wQcXFQiR8EOhn+TYzgYKENV2YAV5Y0aPMc
e50PHXPZY5EREfuTKiReMG7A9z6KZmCpLk3/tHsotyLKTVcGoXF57aVx2kS+MQ79gHlEeWsi25in
LV00pNo4XbgXzFpvYkBJ7zpNNqG/v8oILXFC7z/nAr19KxCfqTqNTXZ+l9oDSJIomx4KLNyVrP9Q
RkCx+dfGPo4POiHJ00L5MjbsSPXaM+RIKq1L9xo3qMxscwfGUiug/FIOO3aqhY+bD6JL/m4Sy6WX
1QB6dTxnshEk3oxpyh343WVkq5RcOLTOsN3CL8l0cfpEo0hCjQUuXw1ebOmeOvpd7e2nrXQKhR6u
foYhRgfwt/DQTKWP79dI7gKPIJeoynKOv9JNwdhFGXUXPPb6NczoCXZaVwR+FkhNeHhdMjO4OZvE
dvXQdg8XpQXHN3ZpvSk8Fre9yuKN3m4Wn1xrrKDmCJ8GTFUQiChCTzRa9zQszgQuTQAJ2y0bOxI7
1bc2/fGX8p9rryt5Hr25ZSh9zsUV+wnussJ1XqyQQ3X9x9IjJTm7B846d30SHK+Bq48axafc8a0z
ZBr4VKqxEzMHODvEHv35oZZjEngizrz7OqjkkKrBlxuPGyG31Ko/SGFdLGcCKEyTxZoDt/8GZxGv
O+0ebgn3LgChc2k/c2dFtEIcmUOqocmNhb6Tz6pQPzH/vTsdKm7LmVzTiToVjE3yjGdms0mUO7Gw
8TIz2B64emtZfyGWTI5eyjNcMv9iRMRUkZzX7137/di4Z/L4mcYRNX+cuAjE8jpL2cU8c6eveMQ3
+FfYMzokL8tWb8h25+ZsDnz0BVIMJ0LB5HDVzyl/LrEgdf6EUXWTXwbjJ3Wkpt4N+uRERf/KJLtH
3UrJEgSceUEfXMxMjWBJNnkhade/CNBNojEL0r12ZTvJ1QmTpAHNe3RFWzMZqJ1gyt6k5DHIv8MZ
8XwXO8Q+ifnMsUFO18GqK0s6z8tIf7c9FK371v22QenKuQSdmGGF2naK8yOdE+9A38pYJq7unPbQ
woG6W11ygoss0JAsbrjKYecXnXelrrXFjOkvJ1KzeVTLQF4vcW/11JY4wzIOiYud9uFjLmlRO5en
+YmDmuosUGQ0stoJSDdPtfgNKTerGMfy7TQLfY2R1s2b/ic8tcD4L41c7T57UbavNZCxZSRBmmhQ
hKJaYPcSO60aonpgt2lKwH85/sRKk0a2JCTP3MT5esABdDa4S1MBvTBSh0QfcoBem8nDxk/R4jO+
NLzE5zMoHkSjOvnvQ+X/yvQ5b8sG4mvzzQQ65sFkagI3DlTJ9Jky5s6UaCqeky4kgvy8xNdoR0US
PF4q6Ls8F7Vu7/FA3+AtfCRSmhF1RKmlsaSi+Btb76Zap50J52Gp/eCjNCdHxRWMKpGENCCswBT0
OsRtAxQT61Fl5bkbuxCpyYnrhLXuA117BcS5A7r4g8ArDxim655vC72s1cMwSKix8hlnb1T6nsef
kHFPSjxH3MGowdw5ix2vMTgyv5nHRpjjbk2JMcYhT3NTMzIV9C4cpJoCEHokI97EMCK0kOFpf2wa
eyEAQ6pocM6mOqwRmtoQXnTjmOJEU4rtxJjhi1cVGbp0BWxaQ934Vp+ePWKwNdcRUFaGULF9hOq5
sakfCh8bAu9nXwD7GYjga6LRDim8013PNzetIftTlz5di4fQAjad/Jqyd31fU1KoB/2SYdCMoZVL
KvIle9GDtMJdeuNhFyrWcNBpoHqytuS5e8NNPeFkFymkzRQwayxOthFoyq9G0M/9nCHeOTA3zQ9Q
gHMF27jiFn0PWkXiRTQ2HwWHNrEwEKfIXKkmEBaNTe1IaS+QivY0udmqnHF2r4G0J9VyrRFVKa7K
HHyGlPfrATnSaDnNyC1gJNnyU/1Ce8eYlaviRNK4YYDAukVsmlSXIR6cHe449gkAjA2l3/1wlLaI
mhVBY/H1AyP31IiiEblSRkQBN9zShGZXjbezQyLMpEyg8utspeHnWxWmRaZFnSrHLwjk0PHBZt1h
UT6T1AWzUedI4Gm+DDZEoYCqOy5E+aIcq7llgxsCylXw7OAbSa3ZYOxmx0aC9dtpKQE5fy87jjHZ
JABc3KOHpN5sQn/FXd/gvftPK1wvYnWgd/56TWK/N3ZxdhvPzY1TSXKT8rZjyY+qHR56DHZA6aA5
JO7sPycWJ2LeawZN5XptG16ErRL+gRl9WqhgEqqs62QSbzhSD0EDIZYTW/WHlzHkBZdTAHjqn/zB
ArTjXQ0yeSJ3MeOpysdy6c5glcQsrVNuQ55sGYdT/mr4tyquAD9skfepnTj4YJR8XlKBid9LqUDv
yLZQOyB+9FCUcWwnf/lduZvYA1rTZ3UA921kgYu0IrpY3HJx1x4bQd9nGZOE48vyWToeOpP/QNMp
mS0jvW7ThHPVzBu7CYPvAyzBoT1aeYH8haa1S+ICcb3YglsYgY8oOAnPwQ9GUtzutM5T+IvRBkJa
ayYTWHDxMh4AaT0+0xmoxjYbYuOIAcZd3+xqT6Fp5UoPnpoO9nztiUqe6pBlzdN2zSk56zD7ErG3
ojgwTEqa8LajedtS3strA9hiYvIj2OA24V+KnRhg6rTZVcrq5Bqgts5XIu4bI583H4kZ9Cr7wuoB
iZ8XWFqBP4Uu3Fr1dFltWdRFtDj/pYh4E9rql1fLU+Njs+LK1padgVVHCH6EAykSNo1wH6Zt+cko
CQ5WJT4nuGBCCFfP/mlz7GDPmBo0YPagKbZUINhIshxxVp5Brmx5+WOENEHIJglo5GGyWv4MwMwy
pifvA5FBLu/BHkcogR+t1xv4e85t91iH1goQS6G+xa+8PvlIen2JMKQf4ZqjOMWJTbHUdvxJ9+Kt
h1k9NGVl+OxGIUAWlcAPikc6kVBJcabJeGdQ73mnqBSDHM3VLNIjOeZY0/LWukhnFbJ/gLkMh+E/
7caVF0/uyAJIX54EWMiR1vC+qbKxJRU+YB/Gvks4Qj+YmmvWjlvkl5IOMmhuH803xjAfwJG447dj
dsRpxfA7ed0IcXBM9SpDYLYH//HZH3KiMROP57+MzmfdtRZRgUCSnv3S5lQoXS5NTAOY2pX0aHjd
JTwiOMDsYV+CTAju4BmzliEdgH0mm8LEcAb23HCGr5RMz8nlaQPYL3yG+RBe+tBELIuK7MsQ6S1I
3mWgwsOQeWRbDF5B8amo3/Qbof8Uwndkzjl0vi5kOFWwMS2yo3z4zM7splMOCGXyeIkM6q/qqdlR
NU3qH5++xadW1ofP+s5k/z7Z+jRddENsjw+cU1EnBHayZLegdELcBqP+x+tVmB9vMQkMPmopNrHT
kfIS00o3TIGKmlrKpW2Hn6Mhzuc1FbxHL2OZAcQBOZQZjpSD+bgDXiETimRkuurl1hguDZCQXitg
9ojgkFvkJSiR7XWr/1MJaM5/ErAFVwB4iw5IXRDHbuSAFv9xTYreV0Ai+J//m34/hp89x67FZqz/
+f46pxyYOMeHyvLIekSrsK7poi2yreOtouwmDMku0y9kohEAO7IczmwUzjNETwvcms3g0QBAF6Al
ZvZTdrgAZ1K+8UnU6rpJKSkdL7BSYhrdeUx7NsgPtMmGQm1qp0P60M5TWCUjzjsMknFQdqdNjmUW
0zLImDakvqWpODCaHnoNrquEWQQhL2talhTdv0RiZQ//Kgi0p9Y55cvWYrR3d7uTnoL3FRIxqe8P
m0vhLKKZN0zZFIzCtExLsSNE13WVMySHekBt5l5tN2/eBftqlIysKOlDz5DpHbXdXFqZ6BBwJuWg
sSowSo2j52p+AFn6dQaiEAM51FM0BXpGPSAdg2E4dzoJX3HYhSSZNghEQz8FToYJBwcnqy3h58cV
SeymromIt9vxMF+cCjui3ovUMnECczo5L8JhJ+NWbIcKSGWSoAaOPp41YUXRrO5koZKHjdLHJTVe
SNkomnUtY1kB/o+hROIWHehhsdK5xJ9rW+MNQh1uCwwhJ+y7vqmzinul63lyH8NaxS9zb2rS2MR5
4dM9fBUttKicTa6p/f6/OmuER6ZaYCsYNsdks6uqxdK1dx68QYS0ThzeO+E15IzcBkYanaNdr/Wm
Ypqv4yxwk8aKgPZYz5VyVe4BJB6nCVZybVPIrZ4drqr2z6y9iukP3yTS2Im+IL9r6psM0DlFVknA
yXWKrDo+FCwxNgcdU+23SAVOtJwvjMXT0xQWrRoO5LBGKAqzdROrzf44UXNumrrg9zTocCxig5wd
X2ol3JodGIZNvTbaj1Qi1GnYXwjkc3XSN7JfAhgIX+D3qmSlzr7oy4Ab4OeBMX8WTi3/4DlyOkPI
JVe2Vc4mE60JLeDRucUA6LQ/kAR2pGl/CfdINBMQcBsz54BLzK3jkagNvnfXLq5EWxx2lOg+C7wS
fqKMDrxQy2axUroCZIzy2z4xiXghPgAM3veH2Q5lape+QfuiHzuQKX425snEQJuofk7j5TvvOuic
vYUwO8b9nD6iLoWduw9Uk7U71IIC4b4gPBthWFw7UUTfRwDq0HCtxCej68CN0gMPXISgpU1CyDfa
X2iLzQrU5a7qdX5rlfStLacItk5R0+yX4QukiHBl/lu1s7HBg5xqlJfkF1bKExiN0Pgz+JwA0sWE
CHveyWzerOSgD2m6OAzzeprDRiB6cC4M22XxUlC+TCuZD29Wu/Y5NXWNR05pH+KHmhvBOpmmHEYg
AMrfnZI7bLAaJEa16NEk2UAWSkv/VUbcUoOO9psDrZrCgQSVFva7XBhORiiMy02U851vlqhzlC0a
86to6VZTIBZtTxCVLOUcjdk036nh2N7lfA8Avke6r/OWMdAcBJL0JiV/BsFO4s3jmgq8uF78vQ9D
nkr3gzCHt71Fi3F20W7DWRFukRrw3+TBWElnXQITNlGE/IWGsHa/r3ES4+Eqb0yV25Q2dAv95Ybo
ItdpQ0pqjwvZV1tFCcXHQdkR4Z6o1NFgX/YNqMMS0IblX2/468LXMHLDKU2pSWc103JmWp94zMwT
OJ9XxMTnPsi1UrlhdUQtgoBMO8jdnGxCVb0olkObgNDX0yw+d3t5WwFndEcReoqjNdcRdmRt78zM
HGnsnkdt+LkvKsd0qFP5zSTNaaOAog/ULdrDWInqjRmVSW1G4p6hKjcpET0qruX1oAfkQ3pYG0Rc
dQ4Q7KbdHtwBImawuW/wRhBRxwvmpbxL8r74vrHYYmWVbfk1dqfNEUSdd7fpghFHQkORCRwfvUrG
yrhM+ixIJh+ll7QLyRY3WS+1QDCP3F86BzbOKoNgQoFR+QCHXgx3f6M6Se+HPKjsxFT8RNP2gxGv
N1a8OHu30J2HKeBC4KIXoU+65Nltnfi61jzz3K6P6FAmmM4JO3fdAyrY5q69IgrGGm+6gA64V/rL
5W2LVUAfTzBnOYhY9b7mtCZaZF0/SM0Uutwy0Keby9pKOMxmVsERlnPN5ayk9FyAR/bAv1bHj2+6
ce18oiy2mf1wU2pgOV8zzQaI5LO+0pgMGLwprIahvGmaj0P7wTH9gUIksfCWi65tnAgrL5+H2BER
24OEGZqUvk9Q1TWxDxgLayeJoDcGmnSaT6mC4NNrTkdTYTCsA8AiM3tTZWCpZXQVtJFii3HfzfT4
ByBxtZ04f7csbyoKMnUPqYhCIGtJ2PDKUpcJoo32g196N/nFdAXh8xL7MYWnf5n/ZuIciemhAGbJ
MBFxGw6Tk+YWdfz+VkddMgxnfPXy4cbVshW8CD/rdDlTb1jQe4CYJ6hu+gWkv2AAlUGBvqmT4Y3U
7OYxPTR2BKnogD2cPZUGwrHes+OKFW97rAgbMZj/qcVThWqXx75/mZ0pkfube/sjgpUyf09t2VGr
+R5vj5piT9+bsNH2NgpEht2tPIZqWDA2NGX1aY6uoGR6/l9/prDhlxDIvrfMVXyFbxWwZ7WGPr9K
rY2nHFcZ20h5w7Wh/FBoo4XSWYO1/4TRVabdTrDj+q032nDQudMY2AVUnTJKcMfweTpczVOrxg3a
0B6q3lf9cTiY763i1AoQvFBUodL83b2LYMWAqa8iNJnlNxbLNHXM2DM49aoFvmMea5+pkFNqFc2J
6lPuf+vDJnb/vha+lTNL5VPKiA4NhoqLlOsQdxhD4PRmr75P+zxQH7zNQ5LNOQyn1ixraJJaWwbd
mXO3aWSSK0Lym+VzgUsjrSznh7afUnN4iHUb2uzi1WfDBXnr8uUXbWJM4dil6+i6O9bvpU5m5fDT
2Rv45Ar/rABfIm4NH78jtw6DWOJXR3Fba24ojmIDX27YZsbi4okwR5+p+rMNTqxqlXBbH1wJY0Bx
kwwSYsfhuGmJjwtdhKr7akmu/bHlaPLXmZuZKFhHxQbmhqKGZyLk4X2Xz7qHcClD9AMXh+oGUIm5
TTCMcn90bKK4/Br2TzVzye5MOu6OT6chLTuR294E3XyJu/C3n06EFeagk1wJYR7I3koDeS/Y+Iqc
5ChiEB9IAIkzBEWYIN3WXvmIX9FFBXYrX4iVmmaQ0oTRQS8hjwOlmydB9lbi+EIXm5VZ812S+TbZ
QCLJEOAoAFgkCATysb0atHpC7UOuMYmXi0nrVz92kzEMs/RBdkRgU2dVXAmq5tR1PoW456TbfMTT
7b5bgOn67Cn6ttM+HgDpOWAFUHn/WI3QOYGVXPWYf7nTXI8S42ZrlvfdeVUjW5VNO/pDIOVH2qmQ
5BOB3DLDpen0z+dPp9nXMaMV29IsTUPaig1OnQIQ7pqBOUIsUCppnE+1palfJBM6sd51WfbhPwUr
MwGU8yMcz8wMAih62zYJ/PhG0PYNW65wFwzMRdZx2+O9b93wUaV12rGLgWfs+2oixXiUrF2V3jhr
TyfFkSsdc6Y4QtqcL9lOytQktHAKxrueWR6g0wNYy5iyFnigVgQpPqxhLTERtyC47p1e3QRMD8wE
Psp7qxm9P7rENkvvaGBHU0UN/64CMgTq+O7VciP5/2pcIbSJ6ZKszLuvgjl+qMZ7Lyl3wxtYKQGn
DVdGG2cCzBSXCIvTSVt/Q54wWxt6lHxBW+HE3BmFAeKTQYjV2b3nJSxI+OSOL76T/oXsSIyhp0rt
/LBi16h92UlOMHpEg+AvMGBqvkCy9MPJSvFaKXbuak0Wk8nZQUqYyREZAkNucVErXsz891nmoyS7
wwJfMbRV6xb561G3IEnGEKgytuKV07gWubpfKBeql9gGhIFrE0wnxl/tNAbDO00Cz7Pe8BaO+tRZ
nOmKCIRtajtsOMZvtJ1XOF0RQdgWUpLYZA2PaR1DTTKTaXzLao3W65Dc9NupUrMH5t6wh2T1Tiqi
QzyDNncuJBvzeOZOx34TCyeqwTtsXU5I34yM+c7cFrKTsXL2QkFWc46e+orRbOz/v+6+1A4v5Eqs
RwQMgB2XBir1YT7SBkPVmK0xbBwcUjYTd3ffNOHoKObxVOF6i804MG6/ttmqb3lYCnqQMuVb/5PX
wVzEj+0U73HpGqsE4TKZckmhV4o5KJ/3JZEvKTvwa2SNQPhDhPBw+4rIq7m1HFxkCcq1WAQ4xahA
SmxzZ4DQn3ORJgzGnhJ3WZCsZqS1XuxcZ+MPC1qixUIM45mGAdYPdURgnsw9pvssy7K/M4nt5ZG1
m4aWSYdM6XUZhbLSfRSqSH0ZWWzrW1En00w3BUGfgy9XzMAG/HgHrz72I+M7LLrJ/iU6aR4ODZy6
AAxaCqPGViQUwYJOe5pzxE+rzwVWs+t/6S0OU4SjU+hENMyn1EajSFSQPQlHl4BukkXNPeXSVnn8
sYjTDkGtoZgN4OWPMASO+lYFf87HDwQrN7TDDdNiRHnU5bQFH/SiQgOd8y8ASBd+h6XYxJA7q5CT
YNfr/Q3QSHWQ7F5o4Yu9DRB8Dh/wjoEqYht2DIB0hFKYiCm4C19gAuD3ayEV606GwWtz5uO3+Oab
nOHcRI+x12leE1I5jtQI5QFrvO5OhUHNd6tZMx5GHWyHSD+7efImS+MKWSwS2N8Gm+kuk8oNvJ8c
1tCcWqb1WQcCxyLyKHZnR1Ke9yMYdfIQ5ccDliUsIYUzLNP+gUfyio6UakDVIs1nAhOj4SU6MWPJ
vKpN/UH4dWp0m57kck+H/6smobmG51/ESCsoxaRdn3XYKqA+52a6OGmza+uocwHBcaE9DiEM/xQm
ptNRxB3rcoIVuSGjrUSobuAS5wq2uQexOJSNkbBQK2Jrw3buARtGmrhOq0FphDCCmct9CNJWNjoW
1vMA8gxm9dAzUJCSf2SpQAgr8n+1bqCMxLL9CniOL6ngO3+COTpPK1IL3Q9s29JQJ71GkOBaz803
v4YGRpea34V7q0+z648uDrmDOIhUGCFmlOfftNxJazo8cDNNm9lJgUnz/3pnc03MIAk/t72oWCZz
EuBPpkrp7Y2v1HUIoD7KwTUYrQKZghm4uqLiy3XFy7qIkaCGxg9wZFpTbXIRG1NQ+3eQTcEm3pKU
DWswIw5NVsTqJ7XYnNyP6S/lEtdtQMiaVhlEmNk3dI9NdVlHeNc5kxV3jRqoj8lwMfmQWqj2tP1/
r815meYYxW0gYC+VL2W94hjGFSXcbB/BpxK0L9TMRWlyYz/EAqcLByTFf1mrdmc9bVpTSgDltADd
TKUhcSf5KefIARweImNHXeSb/FsxQ/+H7Ie4UsR+jmCjtNTNzpXk1JjGG/AlN6UVl66NRH41DbLh
iSY0g8+OZQXQKiwcNMv6WzVn6/eorb25t/2iHysOxrvCBrsxTmEtDslNRfrWbn2iwEpKBu4urvzx
C5tqdzLX0yTs9UEfAgpgVFgCpPek0T0DVsLvea+nB/0MNZjh87AMmdH5J8upmsHvSOsJldk/GHqS
7vd1rvGo6tgS5hfUrB8rAfIoPtEzcWMuzx3kSO+rAXvZcrNyZbkoGbpD2UNXjH4qa8cyKY1zsCMW
TpBSB8a5mmywUKe03lKzYBzHb22/gEioW1pQZaAS0PDMxkqoPcKIY7vm29JHvEm/qhTxzvQNs97l
r7xyKkktu5OrYc2j0IF+rCrV2dyHHNf2JYxrh7AIF7rSR31FR+RzkSCR6YGymO7YzSNYPOj3ddgD
uE4etHRWCvOtlcNDdxZMuUoEFioGskAD46juZeB/NPMSpTZg8fH+57q+LWlNhWTan2XUlwQjoCLQ
t0futu/raebj7maBUOZRKMci8Ue1FHVPsGfvTY7lCDQ26IdUd34q1uMziYrEaefD4oG/pm5EAuiG
HwLkgjsaiCz7mXlGwvFVIuyLsMI1MKWZ99+Nuf/g4XoL9GlPI+rgHZx9ZwyfwEtjDfLuGShlYAW6
t1+CQOQh+P2uWuf23bCPZoZ9SXHQZIoVygHbHlvDVcNmw1Ee4XUwAX6xdHrvFPK5lMei2LgeIoFP
+qsV1K3meQtjw9UTHTlkdS5RAG6G1L5af9Lp4FGAr49k86UdMhLxtkhqGPUwBFUH2SUhYTR+1Qea
HD+5as1qRWj0IvO/USWSvrCQpSzztiobMXcAB+8if1pnpQYnwbts1CQalOB/8Cl5WxAtciM9U15l
RAFCMg9sqqoHC5/dQFedIoNHYHIyxEog3YCO2IIS0kt0VPz9qpufwhgCcmmMdA/vI1JQjOhcSdcE
pAm3tnJR0ESu7O76R8G+TfE8Ho9ELqFB/M5lE9Nv0iC0AElyCzblX9wTWnJrb3Iqd5FWTpVhhbAL
lSy8qk8hGu9J6Jn6bgCBoJAWPn1wb9Qw2rBM8+JA58Uw8QzNlnxYgwQqXkq8TnUysVXD+JcsqaZS
1yr2KnpN+hFz7SCVh+FmmPaVU05QUCh5rTiSWtTA7muUqqwKxvDt3E8/knfsx3rkoK6DVh5Ce/jp
QuvrdsyZZIYUst91RCQUy/sbGOHkmYOH82HX+Bfi7Z30S1+0mLDLMKwSygKO0af6k737p22bOKX8
3juFJUzAG0YDsovEYFGV2XFk0Suipj8b8k3LCJG7hUuvLlOymATbT6wOOp1m03DWRQcuMuZrX/Qa
gYA0gQXQGAHyC3jBtNU4gPuckmPi0kWr3Cl6fFDeSJ57HifWkkxSSZSgyFnOupmxELfWAqifaH4C
9N9Av0D92BXt/GgJ2zNZg7nMYzNHcsmDBaEsAo2+h3mZxgS1vNV0/ysPoqbrLZCf4TqpGT9+kUFe
pEq3pt8Ihz4syegnAZWNSRv9KFBr4s4a2DKD0MQOfia4l4ksjRL/Qt5Ps7fPZME8mgHoCE0popSH
wwtqlPO6AHrnBEVQI7CkA2CTsmbHduESnYcbuQ+Y/BT2soxigyRHM4WdCDlg3+WVJAvwrkYlwHG5
j7IoiqyAfWsS7jCjylagTyPzQn529iNiZFQole86z/XgMUcIx5s8ppDQ/B/xhiyXEpbhNq5ppvmM
/l7iECi4TjqUyaxb4AKDf82YgOsODfzv+3b4P7vuOQD9F0udCxsacHgh8MvN37Oq8kkeaUgN3sGe
oJdGnMLs1oitjEE9J+dlchNWIoAHckVXQF+keKKQEFI4U32P4ylhcGkeE792yiXZ9eCtyUWeWhgO
3gXARXWP+qQuVIrxSlkEO+iw6+aMizBp9Sz0DzdYcvR+1wXbpu8wmCtCyfxEO1bM+WKbtHAtCAMr
FSh2pVoXoefQ8qrdRh7s0QihaWevfug5UQSTmi3jFxlBNnuLc9rnYEGVzCDaEK/sBXoo1LoDPbYG
FQak0M3y9nDgtNg2kxh5Cw5qiVORuiNMjQgNPWVsDWjE7Cl3jr33fWdL7bXgvwkWQDTOeVu/Q6Rj
LR59ftV2JP4TcHXuSUz5rjspRU8joVoW108AlgEbfhKVeSNEW+MqbPv739aVi4jALTu/kxMBR5qD
HAKVnyKBF6S90StuEgKzG3NST2mUoVu9f/VZaG6pH9ZXYK6xTNeF+lWqYMLY3M1OBXVQPD0R6rPy
qQK77BRky4TlO6MPEIhCBuq3wKSTT0EGEJ5g/KUrad7k0FRVCmeF0Izbpeg7lmCDTWwd5fS2O8sp
lO+nuBgbxA1N57uoGU9DvwOv/QfCtwQCsyfxPDNF7pT2lEBcsgF8leTIDkG+1PhMjdBtuW/QKnz1
Ihars7IhhDrGEyKNoDO+gS3RnqDhnstFY4KRcYXk/jpCQjPOWQnJ+eE0sVdjPcUf7oAHpCcsBVZK
vqevYKpbyNEJdPqhX7yi4GgGE5NV9HggTA7ooi9PgX7sDbjqXQR9Kjqa87rceY+WgjcOHtg+7swl
GSNCy4fhkmFowsCJbF2tyYbRJJzKg4AztNAxrIRD2TpyM11f5XNpdVhZ+1RVqLNEPMjb5fVj0Jh4
lkb3brZZ2BET1PyX5ahrbhPwW1dghp8TtYaQc79BmZSx9JM+kz96F6mQ0QuMVZXdRjAsXcK5ZUWt
KGROk/U+0YM739C6xmVh478bjHlWdN9TzdXc5w9mZ2kAfcN9+f07xd/aG4zP8r6ibc/cUZf/ov4c
ZNcd5DMhdVqMEU2jTJo7Fus9E7M4A8ImeGAXd28pjBRFEFoKAxqKJhwNrztciNMZJVJ/obQZUhKp
VjS7aFe1oxgddmwOpZ/iFnlE1+zMxwIkrkj8co+guUak/IPukxCuA2k/bIZAAi4MrWqWFPH+tbrJ
o141PTLilXJbZC8+YXkWzPna2NL1ODmZXO385r0yrBVAuZnT2AsLz1H+fY6mFg/nw/fnCiWxyU3a
ZpEMqxAoqoX9zfCYo3Kxgl0TRpVllbZYsgKTnlqutPSoWoGj3kbCPInBvTGHbsf2oDlZpoGEbjFj
naSjUkgm4aajfsaK7wZoggLTjQ2eiNWkXAsm/OyFYRDNeWRH+tSyMC1CdYjdPt43UdOL5YgGFMNE
19UjQBs+SC5nW2o98yLs0HNVeSizgCZdxts2XOuD0CKUczluz9COSZDPquHyMEQVdludupFqUHD0
f5VThHg6ZeYCkt8lNJsKmJIwMLN8x33DMqQRuTDe+Tu4AilVOWlmkvKTKr/hLM4Y13ihatBLcue3
WOBMMOUEVP3SQGiVUuEvwwkuYbeBK21JphXRA5QMvtDwt88q9GZg1SZxIDUwLTV29nOr1/2s9J2a
sjcDLMt9j8ewrqZd/MEwZx6FaSMgGgduemMaTTBBs57LpkHw/lHWXBDdAICWK8vT16JdO8N++Z5N
BGB8v+2RWFS86LtoJD1pE+ZIwltyYKaZ4Dz2GPgixFVf3NlsCij6X5a1dCe+3dFplnhHnXXe5b2o
NNNlWypvYvD2gVdRXSjPp04UzThPvO8PNwgIPg1yEGA4OYhKdyz0LYphVVYBayI1Gvae+aEUK3hy
J1LMZUTMHKP36WCwjrSDcPVOPZW9nX7AU9MqPqc41wl1oQZ0fjDx0GRhNCZplMLRKECg+7fHNOo+
LZwiQAf0MMNFEViMeihJ72ZiHvAegVtfw3DO6ndDEZJ+WKXktg0qs8Lm5UR99mRN1HTABtz8p51S
PSN28fCvp7v5OBVs6O8T3dAr8itvaFMFQhw0UJRFanLt/Qkbx/4uBZLhBRA4e5YLWoH3G0TiUT7L
F8ZnaTF7oYkutPwPNETrg3RMsaRMpPwkXbby+ZVTt+AC8Dfjz2Ze9BhRPqR0HfcrnByHrRcxATHw
JZEgmYB3H9dHjAFFWACkcfMOIlJm4QuDsqKueGpqKs09V679XoVfoS8EtfZRi77i38vLfsUfVS7r
FeT8os66T1Mq8tnnxI6CdUV9BKprVj9gwChEgsgrgMklZaLmkSBfP4P6fonLFnal8zIjnFYOfkA8
PEIM3e8ltgjwQafV1TrSwZrt2NzPmQ1AGYlT/lvHQWNH1RfQU7WcD76NKgr4aaxAk6TYtfmSRvf3
fycuvVuX2PF70vRi+qVHHHoM4pLuiGzqq4CYyIKUDAG7gTWK60SzTX5wbWU/kN8b1rfneex47fvo
KcJ4NOl6HjWH+NIpgXJu0odO8OrkJPv7BeyHd5RJKTFGE4CWUFfk13+sdllmmp5X3OXybxP9k2+p
2mYxyoDmgXX5GcRPIE8DtDhwNWWZYl80qgr7AwlkPkCzM5RKKnP428qew+9BDMyAs3T7KpYz5iln
9XdzFPMaGi1zl72Ym1UYqbCiMjo3WcKizkVCYm0Mw4n2Uph8WeAHISWTzaFJtbBVmSYS0RU/lZwO
eVsqyukSsR78rKLNETDScAUAtfTy1fy8v9jGEYi7TYQV4ezHu4RIQe+5PCRWlvQzOf+Fx4N0IeOH
U50Q+i0fHiuoDDI/Nrtj3t9vXrFLACS5AWT+guqPwCAGnd0uR9MIfYxLLLo2rXD6kvmk7J4FvZ2L
H6s1/hqvA3V/GQeZmIH0rVcL0MP6JRh1Ate8AtcXEXD0o6di5dfWbq9Cb15kJO5AoFAMjXNa4F7+
N8fF5HZrJgYf76DRLCUi0959T1lwp/Oodzch2TTuBri64AZ0qZ6HqOjPs6Jr7eHdH9xNUzZBHIVj
8ThDDJ2i0w0sMi2Y6E0gilrieYgl8a9c3ay8svcm6j2rosGGXtgJOOv9DVkGDt9F99Tg7ur1I3p0
u5v6AACW9ip4DGN+WFsS3C1hn5elMrpUi27Z6N6bXcwSib18zj9ZxxiTNcwJk0/73MeEpGX7bwWL
rui0NwVAehM7FUvJbeOWFbQ1qaCyU8r50wAuapRX1b9JNj3k0b4kb5sCQ+J8vvgNlBC7UcDrMz9X
Ur/I99LtxNwLu3WxIqV8aZ0on0fkW1uH5wtUACLSbcQW3vdzPGNARDF1h+3NCXRcrWlBRTAPG/Ij
btPdfCm8wDZ0r8LzVJJzO6CoVnvOHV76Q54QnN6NpqO7Kl3dJn4s01SoIExi+FOmp3k2J51kJT9H
Z1sDfuRBzHonByM/DEGK9SfhgWs/obEU4E9ud3pjk9NXscdhHacK7aWWwcSe942JmN5r4PMmUfO2
uKlw8TGh5urLkGOOvwVt1C9VgmFZadnzhuV356aP0sW7wwtQSK4TyZH0NBC/ofzSCgEye5d5k3M1
Vud3m1RdHhozhiGwIJWs+4NLWS8WTBtfSRBobZA4cyWJ4GE0yDh1sC7nZ/WK48J3+9px+1WbYIlt
6aoXyLI1+K6dh/bqwUE/5u8Uylx7OT8QkgFzx30ST6H0a9Ea1wLNS4xbQzLIPx4v2zGIO3DvDtYP
BVny/p8rAdzgRcTyTYiklC8KPnA5FhoK91MSZaJm2KmLiJ8GMfV3LRrnOYP2rlkejlHnDp/MFB6C
Mj6E97OOOxnOXLdUatL27hJg65slqOCVC+M7PEYjg7JM8vVtfuZdphq6Bx+1Y0DfpHAhDY1g9eAw
CQ7oNCod08SnQPBqYCuyAiE7ved15U/EyF6Rvuh7bZz5lFIAFlmaKoGubAfgjhw40JnK2TAlbQsW
BIqeA7pTnxY0xHs7aPJgYTwGGjmYJL3FFtWkTZW4glzhOmQJdVxq7AkDlwJi1xpQOuf23oAgLLmn
n9juWh4PfhdF+A+jvg+BJWNlyhUgDf0ZklYDVY54b3b08gvAmLZki+rXKgBNBkLUpuER52308ugM
xFTyvL9NqvyZQCLe7HFSPKWqGL4uIhQdfwq07Udx4MtbU+9b9F2KvVqstKedi4gPF6k1Nfin/5On
UBusjoaqIthosR8knlyEx7EtYIfJ6+evRXp60heyjLKmfbkFtvtkNt0iQEYMfVp2HpWPPP9X0u0V
C1H9C9j1x+eLdG5iBydlzl6xSD37klGFrTUny535X4nnZhZrrhcHBoja3RE5Ha4gL9ujDTO7XUtl
2QcRNKER70ACcqrgLM7F2xnSmMFUD/WYAXw+m2MYkfw1RSibXGg9By+BteksYCvm1JDRGI7JsmJq
8hWGYiw5AiB2WrzsR7XMqZC9o8IZwCMEIn+wNhVuHL98Yoq38JVs8qOa1Bu8bZb9aCz76+UGV+Cp
VPcEydamrqmfXNQ7TnYHjFqIx8AHoxPZcGZv0n/CsA9wXdAnm19y28Qdy3VIWZ7kEytdSJULeT0O
ZHGIQZFRTGsrsBR8HCWVakNWSCLN8CPYNm2P4Wuk4L6Wj/4EmU2FK7yVDrt+PbQSlgehqN0iJz3M
d2Yx2vm5O153Wvz/788xz2oyLl2pZ+QbHT1pmQTJ0DVBhvyrfnKUUe05Z5ziN0k1R8h0N3jp6fZh
CLd5D/PZ35QmkRkIVSTbQmEPm3Sz26eS3Twoe3vbbxXUWleRN18CkmcOvl4tY440YreUIhVvmp/0
qyZtzfIy7J6JNj3U3ByosbEhcx7nWJdJCTtRvwv85OcJwUVdT7/bhxc7Utx5NKZEJuyoYXn1zyon
8HZhHKtloCJPo93Qqb0TTAisORH7c0HDGZaotQNIaNn0lI306YI8JwGflEVZEgtCdZRl7uwOoEPS
TNOX+SrMCouIpfs0Pqk2UvWVKK6Tup3ka1tlxAUQEajV/RadnfupRKm/8n7uTqiTYAgrB9xE9Xca
5OvkntTxo3ktwDWKmDe40QN+Z/KXIg26ELcAyXyziVvrEEi9/8Hj97DKLIxJU0RwbW4tHWHnCD/g
SoClJVuxlIcgUwG6O7wQCCiuPDoqTk+79O1DY5uu68Shsoc5dMkyg1l7GcSS6d1NJ9ErPfIRGqhx
9VDOjJ6Ip8XkEmjnzKJpMInxZ4l1Bz/pSF8t0usY89eB60m8HwqO5uWE5A0p8Y6+m+iIB376vdKH
iO3DTBv5R+ZfLZ6SlSjt2L/OrR0J5IoB5CAUqjn8+9imzQ2/4QdCpHqr24JciGQ3XF7+zfZMVWRe
CUYGCGv9P00UzkFhV8tACo7a5kIT3qiylaqPlRHlGz7AjUjN7Cyux3Rvzd0u7xZuzTMM5YJLyZZ1
fKahjooDmSPCO7lSvYo2OQtK/7g/5xDTFLdd+lJ6v4+mI4nJU5AR4kMBeT+R+qEW9HcvjuTbgE1o
lWPgF25KHceoMSwpPy8d6+hRvt39GGrvagfsM+QT3idvjxZ47JMJsbjldmc7gLzso4W82TXvOaFO
CD0oSj8AeBSTXNfrMo013klV5bvnbe7iFvAXkAdp4wTarNmOMy7VdPFuIBuTqu8T6FzSs/3vabWK
nz+6tiKoB6eOWw8afduK/aJstKrPa4buKVA9EbwWhHgsRMxdyUcwNC5TQJwyozdd6XuQSsh039Sc
SfbM2vkoVK4Ide4pZGzxy2dpDz9NXW1SRs+aFB2lRyVvhoi/g172rOFK9KVLTfrZ59/lTasBWyMW
XpM2ufY2T1SyhRrkTdc3AN5kEPM1Vp4LlbQIEH88PRU9225VwHmPiK4drDCqjKBHWocJBaEePtym
ehGvbdup346+V+Q9cB0/FAlFPJsy72PBpfLM+nNeH2kY8WkbEr/N7tODxpl/FkHEiP4R2UC7tXaF
aZ1e99k951qTbXWm614dO2yWbIdxodTFLlQP5+rkI14Tigew/qfFJ+oUqoQNnu6194PKae4cgZMT
pM8nwFFplf3I+rvrV9o9smjueIV/FWIXLVpU9c1LPmVCSg2YmL3Up0ePhc26HytXBADC707kmO+X
277qax4sxn4B8Kb8ChLZmcMLY1XLhG5T2eUTodIe5N+jYIiXnB8moRVRYwvlHfPh8vdNaRY1hnFn
9C2vaG22hRHD5cOBp+TCBr7Ox+XWah65Eu/Z0cQyL6+Yhy/ibPvQ5P/JcDuZxARwxqSOj1rMsGqA
b7FVbV+libe4jvUvpIcv4RMq1tudpu6X3eeJYQABkUwwM611xnKw/Miui9DVqvQdU28XnNLXoins
/ZzoNDID2aJtSYG4H0HlQe0FfF/rrMReHAi68hd2QZJ/mDkUxjbSBhD9LC1s5KOjJvN/H+UWnFR0
DxP00ET4FDGpFvL6dc7MY/ZDcswyqXFn05eW0HQQ2MfporHdx8O02LmjF3rNHTMSgJ/yUIDQwlwc
ZriFAlGU7z0bKFYiJT/6SZ3k6uE90KNs2U7mt39IN9jwBy80eTFkDGuXRxRLdg5gO1FvVEMQgkdp
nbY5bL+4QnoLA7phz8L1GB3gV605w9D4m5lGy2RQ+dYhEWaV0EdlPFOquTOXccOsb8eXRtIZR8Pj
SP3qc5l0ftrOrJ+mRh7wWAVN344Qh6oU1Bp4iHQ/IhWUUGTyVI5+2OMWi2HMVzwXDkjIrDQ3YNeL
vHxHVoc5TZV+2knsdxm2+x3tQ5cS0E3gek1PH1PenCFDPB66c5Rbpm47J2RP45ehq/nxf+hJr3zC
hp+OrKzCts2aR4lBHOtGn6rp3IhC3kY2G0ighy4Wz+Qea+fmsa4VlvR1QR1wTzpSWRWADUBa2ozq
mDmAX0xh/ADGCc/CUsvAtYfyiC76GKws8ioaMKa1milJSXIkoHrS0b1Yla5KWFyouY+Au3tm+JK8
jPEE+0PogMMDwMbxYSnkceTUIA5rfj9Gr9rChtneKczCqopNGmGPHgEV4Fyzy5WYQotIs0O4f1Aj
HdOTOVaufyZQ72ZOt7RMMH7CGvMVkOwc/AUlCrgUHLa7+Zsnl6F5SpI0deP+9OSnjiumQv88BOrW
/3RIImtx6+t18baLDAUq5ZmNr8uHCZfwNKxpUfG4Bb4TWhuYvn3xGRIHQp9l77htjFw2Xnzwd9pf
0OS8x9DSYGnIUu+3Ii0L5K4/gmjIHTLzGVVgMAqlQc36gljYyvg/t4XPnIpSM7o/Qqk6J8xCyLRa
8Wo/P25ys6WKmE5bUB/NYz2O3IXDh/dsmQlx5HRagslBGvrbH2Bo15bsA0+X1byHa19vhHCn46R8
yzic+uvfaBDPIce3EXtGh3c5mHsveOg7yh/Vx5OH1us2wlI/5NsoLhdkNwJ2fzgOhvlm66JFkeml
AAdYJUnKWr8EuHbHj9BvFKyoI2H/LAmyA3RafbjA2ZxEKrcOiJgu/C1JTGL33d2+wp60qulk53kY
hmeib4c+pbIL3DAP4oSXnzQQV/mAuHG3CTCd5WR9nTkLR76Jp/HvEKJIRoH5VCYMgGT1oPJf03tC
WlOX9yaiEGt7TIOua6e1FBeFJ+uHYRpYUDtabREeK2rNO27mCmFoVrRWk/hIOXostHPJu/qsN3Ks
tYHLCz9Au2UN9W2OwZZnxrJYqlfWN6odmcx4ZV2n9fGfOR2IF9qfSRd82Z9S16VReGCQ/kWcwdOW
z4/mWOjpVupHkqPatumsuVyaXhv6d5yWAQa/sfe3dQ0MeLHwRxkmSJQk2+mSNmkOB+zYNLF6PGjo
A+THE2WGhk54Oe5XyyFTRXkiPB6v9Z7Vzgo66EpuFN4Le11eOMBuJODnLUxBRA0BcTtsSZz3F7cK
K2VywgtkhqCUS1baCmCByJElcMdIIwvvf8qzdQ63ddBNuz9PJbcovgz0vW+udn+H19cICg27t84i
LELeprtGQQZOeL9mh3sdmFoMtJAThUFrqOdmXWaRcodlxfcc8L6+/eb1fEPg/AgjAoL4voiYUV56
rAMN+PJZS3lTSlSPAfdOU+Jt+DuWvwKdJaRtCmvrCaJTqOk7KuH1KhPtHCMFXA6reEit2okDf5Vw
YctS2QlCC9BPQ7fJOAs/CPAjTyG2C2FENfRwrP1ONdzaXzE/uwtOZ9+oMxtLK0H8jD+4yUsqLjd6
RgExDVuf1Ki8yZ8dzCq+vzcHtzsxOkx0mwnh9nVkpWBKQWXql+0aiok8vLwl66Jl/nvQpJDdXyYS
r1AW3mU8M6LiGwL3izcsX8D1piPoLwnzy/0ikl6Fgr7AMZcVye1q7zbQVWZ3WUvm8tmI/HXq1zn1
RhF4u36EzfJ/OOrntmcl9frqB3kFzk+MLnLyD0tJeIZMWprnx28wolYyvrwUm5j+yVHSeqWzIUeB
S7ifbTDIIBswv9zqeDzFPHHWlnnl0wLbDtDC9IqtXM4ZQpT2ET34h5v6GFILPxecx9hJyJvy52pU
3eH07SPz9BYJ9x7W0mDi+ZE6Fxyex59+McqUFV6DSbnb3N6lOA4iNvL2kZasB9Kjk6V7c4hsG+rj
w4rLbZskmyk0B1QYVyUB0jTwI9Hw5suNXSvkyJO2ZCdUJk07ue9ruV4krKLumhWOZcChOZrhX/Gx
BQq0rXrafNocDtN8DK7nfiRAD9N8dnOVOpMlfhXTqn/Cl9XEKr/228IaXQ/QfFcsGoAZz9Pb3sqb
0NQunq6p0iTJ1LvqU0XlEgWoBaA00WM4zSd9OLNBwTDpH3fDxdtyB7SHyFmPU8G+dEV0s6ljyCNA
xA4XAAmczM91iZZ6T0DDLKxIJ0gMYJdzU8RbMJGJnDclky4v7cDxF64h/fSaV4mFgxQQkvQltaxX
6aBuf4KTPB7g0THMJeC0Hin4qPbqye8keoyKpvW8H4ZJ3b+xZvZx6JYSC2qKdSDHQbMYx1bYODPz
RR20uwbxgfWbPvK2HgA/mCsd8QAwI64ZQl4jF5BxAF/cXTsLvJUs8kZUK6Z1Y6jZlwSSk4hp+Pa9
JJqmq0haMFE2ZtxmN8IHvmtC2+cUcrezkDgLH0Bl1deWrJqkQL4ocubSQw36YhDcZZB9tm/VRTIV
CWIArlVc2i0Nmn5kTt9mP6izsIos77GcAmiHp+2hkuj5p/yCGwyKG4W+hG+dsPp9d/GCveDhxD/T
Ky/ad8wdXfSY5gQqeDU20I/JbXdeW82Jm81Ja9yFBddC1cbpHZhw+1Hzsah1ZbPdq2xx1xm3c7sd
kc2uziuk3etG9xTEphohj3juGoNOUcK2gOB0gDZfAEfYrnIZWOfyjEVvRR7phZH9htK9/HpGzKED
Erefh++oAh9jlaWdXpOWnTe5ulXLR25PxxgiDBfJwT1xy+4DXk9rWbnZYVPUYU8DtqZ8o7GYwdJy
KU5S1ioi/rBsyWewS66bL0sgPiInNXjtOXwmu8gq3QVlLUbGH4yz+yeDb3XouBM4zujrYIr3WjFX
MJEtBr+tadx9umGP6bWGspckD1KFateqeHYAoM6NIOXzLpSqVEvcMMOAJSUpgTVPxbnaRS2OIglX
9xnu1NYTwMwGJ+K7GeJNwSHyQPFLB3kkbui6hUDtIDixM2/XvbsrJouyczPdKcl67wmmhGM+OLQY
uBHjPrHNw5oaXK+edwQ4cMwVRSEMXRKNiLeigyfzTwpD+/TNKmuzYsDRiqvHaS83ybJmnVM1kMZt
XsWIovGujWdvAjzNi+ZL8z9oRNDQ2JIqOx/N6wVuGhGAYkluK3j2mQutCEFSdY7Sn7azK94ZId4l
6TwwgRbThO1JbraXvPDLaLIFeqMWxN/9feDRgeUpyyeuxGm4lLws3gBpQkQBbEEcXf06MRuveFYB
njdFEcBLJiVVRuFU7zInl621BkR9BYUL3PCkzKHUFtVDfWPQjyTZsrj/4sNvShWO+Fb1m0Z+DFNJ
8C7l9uXuj1hCOpif/OhgAKC64JfQNBZSbvJK1FYSmhS17Vm11yD/8WBk9zZiP8XvlpgxpzMSXdf6
K9vDxApO32zztgvxhPBKbFypqgP+H3fNVoSVnAryfgLRxVT9nac+WrjASMsMrHpgBqjoSudEthiC
kmkz6qEAas2u5vtX85VNcvU8iCr3WB/mtm5zLZrWIzy6vRmZJTDKK2NDgLA4YPntQVgCCVnbTd+g
GFaGsxDAac/NV4pqS3VPX4TKxCZ6ZgMUDZyWFmNqUz5MCs1QtegwuWSZvJ08yckOJqwdQDH0Q00m
8bim1hbrrX1pN8ubLhd49FNBnzRTdhmI+si8swAiWhJyuI1gAzwjBiNBORdGwgH7aWWZvgNhjwfV
i8YRIszWwqOGpEEEh8a/hcH1wx41yDdonD+eKeD0cYqNA6t7qV2jusOUt3W5X5TE6/adlvvYqrHx
eRhj8D85OR0Khl37ptXwhxaoo9ugESk+4vEjGk+mk6+SS7kSr3ySn9MJDbLKlFTQ5aBb7rSPZwab
Ufu33DSxOAe32GGPFUru5ODQ4kAT7ci2fnPjREi3LLRghO4ZXVTKKzXxNSywDahKljzUtOj8FWrZ
qEPwZKYKkT+gs/MqZKTReZoohrxhjDhQgV0Z/HAgSNS4lEIxQTguSMcEY3DDH25YgPA3i0lHG8Wh
oPNdXeKCdP6Gic5JhCZ9+/AOTfpZ9QDzaBKJ8dHFJAbIl7H9WGvsroyUNfcAdEi/FnW/CLPQPjOv
crKX7Kw2DCFVO8YWAnWm5axgCbbOZ3fBnm8ut44yO6/tcfTuXwDAFslBiKiAM/k5S7W83tVp5qoc
/3D18DLpKPMhPlVPlmT8mZGMA+MILKqh1tCNtgyqmqNfxSroGE8kdKh2HgKkLq4wJdPV1wCtWKjH
Zdp71Mj38ktEpnHs/dNScEbpMl8dPhIuwSqFep+ljDkKvRBkPAvA3CFxFR7uk7pOEGFXPbq41Zvg
014yU0wizxjI8xDvm9rWfSo8zv0heP6h88E03XWlykSUgf1CDy5NX/R/0lgk16J7qgdmuk8akCMS
/GDt8XVpAA6eP+nApvgQC7h9Xn+KAW7+CUG03tCH3MB65mY7XXcTV4hrgF/jm8SVD/LFofP7+qqh
SnZ9C7KGOl5V+dX/edBDu59r/ZgRNV5kw9/adjQueJFthMk/0aGFU5bU2o2W5ijTybJUdV3xxjm/
h+vmkVLRZMH5WEy4aYcucI+dsrZv8NRqh4BHlP5CPn5WV71XfKOThYS1ryh/kKF4MT8i38KWpZAX
6UKiJzQZ+tNbAgOwVNLY9KJ16hy45mOv9InkYZgrffITNn9y7CnoOJp8rYgBSeFTy+abp0pkKCsr
2sbdU5dOP3jGtKagFj3tZXb6TlJCE6YWLJzzkLH0egdUNp+g8Syb/NrKfPRa1n6ntthX8yLV/bMx
Xcv863Y1sy+XdkvRpVms2aMkYVNkSE+vw/c8URnGRxPNwwFzLMkv9cvmkvCPTIj4zqM6pNcdENs9
oiyYnx6ZDTLk507/YhonEBcypSVRZ+Cffm4DABjDDz8mvodoIunr+atXLzcs3fiS1FsR7GHD8W0a
rTLcv+9auePr4MCvidxUFr4DVmaUPDVk7Z6CW7gRvsCpC+hTPZwl8IMxcNOLbhpyWODVmDMRzJh+
QoaY+DQUP75lNTKR//hCLVAX6NsfGkk059Tv4A/Tl1zkk7B/Bxdg9qZdf6hAQ4WuIkCLdH8N/us7
vGBSMvcA8vK2mz/pge4tHHmgy+5EjM1gO+SS6zy/2e0g7yj5+hALAjZ6EBiy+foVyo/LLkqvz54v
1GDfYXY+r8yJHQmGeLlq1uiNhMcnKDS2qUeeRErHbz/o2Sgaig8FvcDcNh3+8AjyFUxyfkY3N91g
RKFV+cSn/r6+IDqM9TMgIDn69PGizcncKYbgpKTKTqWe/L14vD00dl6obckA6R/Oyyns7eFBkJV9
zafkPssNdv+7d0OXqAtebaLuScNFgiFdztRT7ZS7xYg4f5D6rvJNT5TgvHtFw0uJqIePIPfzS9fI
wkx6l/aM+iyOPGo6U+7fdegNcxg7wpZs8TIdL7OyURZi82Pb7MiJBOMXN11zjVTy5prysxcoBV9J
C7KGWU0fN0VYiVR7uyG7c1M8kF9klg3Uo3uqlqe15Zi9f77n21XXvAuKYllK6Pg3sYzRCHrQjiED
+7zHid/7iOINQiPKXdJ5+0kBxOCKlmc63YqVpg/DMnbuZ0O1sixasGlOaPHRzTg0CA7MhVFT1uz4
1dcNQpjb18EDZD/AoqcQXC4BU8w8ueF4d2mpVlOP8/iTv5N7yPnHLuRMpRQ6/C0M/6P4e0cphLnw
c3VVbN/k5f/F4YdxbIVaINz/c7lSgCsIq0ldZq9AijrLQbhzEJM+plF9X7fbLGs0s2vX2XCVUOVI
ZN9aVIX4aojvaduptjP4k2IqrU4B52QPTHlyIF8M9OE50dyNc5j8EcgAcdf0ARiYdhNzMmeMxSa3
kyT9L9wbtmU3ONu+IfFPl7HV4dMLhwRCLeE9TEHQ+qjFc/rlJaLxfhf+vRH6xdO0Ib0dN9N1FipJ
lgJSSYpWcmU4XPwsqEQwxWSE1VN/zAGns3BlFa98vzCisoZxfCJIydvGp1T5BtwYWut2hVEJFZt3
G6tUhJ0HeWDrjI7n7g7BDVNk6mitgNFDMc6lOhUxjlhlgSa7I1DjLalh0Ywol57FMCRwleOqxgE2
aFrASCBcyYXHa04hEU0w/1x6wV3JjkA03Cz0iHNyDl9Xl5tgAWEzWkxF/Mpj5AHTv3o61/6ialjs
O9XAYQSL2V5o/xHjVjP5Ix6qNaP/pqUigLn+6xwURJMAQ9wOYmdkQDXp4D6T9l2GAop6cDjG9tyz
6GYF8fRC2otZCFoZLF+NU1Hplg7ROQyCjX0WUmlASvhbo9jwFYsSARGGVP2d1ORLSM34XRoeID9n
gIquWMEv03bvao8XiDF7HZPLTn4mNcZ3e7iFsmmDTxMqEVyDHwfc0qAspjcEws6PIgCw+ZfyZyQq
FjmILQ0PL9G75t3hUvBIf96s6b213A6I+YJmuAW4Obh5CC0V/oxVLcm3TMjd8s0jtxUeas4cqo4D
Fo3+WMaYlOeROwx+Vc7FqIKdzmxQxEC8OCOE9ELKS1M8mc+4Lsxx26FN+4o4Pnl7aScSbvdbI2Yq
tlQ0GqBKybJg/3AjWu7Vtppx+yiVt1pCPPibJYrD4qV9+vX2SnXXkHQb8v53Ofbbmnh2Yf5Bi71v
xkH4+7ZKLUrNnpOeQD8+Z3XZuvVYBWC2O/mZDYoa5QIq56mAWmx0Qfiq365N5oPacIeSFD5ru0ih
f+lQ8e2zmcZqu59Gl/swivsbyeWETVwlkCPgxrZ6umw19QwDkPlvH3rKb+qydBxbYe0bH5J0b4vi
H1nr3MuA1gGSQ6ZlsJTMlEYtrRdXkV1Q6EIG771d8VnO/MEz/0sEvhN8O7d4wWa4FP/abl5TXUbW
WiIlRFQBfSuEcugWhCeW7qghqDuk2qsxm9Qzi7ctZfQeMkMWFw6SQGIdNCmxH8wAIQaS/T7c/IPj
QvxZk2ZAgHRFp0QGEI/YeIg+IpiVfWTEHP42wySeLh/OFD/Lz/D02Qygak7vSA5LeBt5q9IK0B/V
GMsA5Oe1JOrLkkiVltFZqYdMcRxyCoKKX6EiDqGoojgWUuh9Kb23+vdL9jKG5dqEAmXgp51e2rUD
mywMvbawYCa2VL+ZiT7mC2DHpfbhskS0xJqq0V1I/6OkdVRaSSm9raykZMHzLaOB0BFkoRH1tVhL
5svL2w0hCShDJKNwP6dlrMy09NqqXC7cfXG4NME/fCGhpP7pbEiCTRttTvdFUnmZr/Ttgbfsojdv
7mh6x2Nskn7ncr3ZqAdiwb4jUr1+ew3BOIYOUw/YGqHSKhKg15GQolygn6IlT/xTPc9HksnFa/2/
+1E5IilwDOIZEADTKj8uClTRjytNsKeQZJtmTmYjKp6EDlJicWG1Wohu210YtfugqggaC1+u8e6g
nAhTcK6+4mkjneKs9qH2U9qpqHE4ZOxuV7vwEyq5BhiWReJWvE43jeq4EFaswc6YOdHKD1jRHq0S
aKXlq4gu7E9X/pCScQ9Dxs1c0l1+Wn3zpom4iJVEqNbFM1Lm8L7mSIaEGvDspA21D5ju/NeftFgE
lm2PNA1UWG61duFqlUYfar52nI5LJHOJCx2LN1+dK6FgF6PDJJYS2rgC/oZdPFVA6ip+3qJsLfzx
wyKzmvYb+nZ1aj5R8s7n0OOscrPGXZV++9XBgXkOtZ+b0GsGUgTyUlRzOS8eWBngjoJae+8VHrGs
jSlZ1h8jtWst1Lh25FMFePY+dLyTbbqrUnO4pBB3SSGnUafu+AU1H49eCzyTQCogBXsh9E8SHxZ4
CE8BfIQZGkdn6qPNSc7iRNrdRjw8Po/+6i12BJATRHH5fuZv42EAj9Fdn+JRoAAUbTFHRPyfGjsK
FISvWsiWMIku3aMSf5gthlNHvQtII8S2PVRnIauGC6AVsto9jIvOZZ1A0QjbpwP9lRMUXvdPVhK4
fBDOSBDLLRf8o5Za+/+bK8y7NWUOAo9Ov/uC83pAJWM96sB03FvT+wx/XnKPTZDl74gbgenlucsW
fnoP6uMuSDkgvQnrc28kae/g8Ope2+whrLziRdHVyGqBVlQSfQg0LOqrOJ+uPFtj2476LSKsD6De
IrHp+m32jqimYeLzhmDqjnofw9ruSAx/x1rjbM5sl61HgR8TPcEE5RalmSenAlLXFbx8KWkY3usm
qGVdBx+IqQpBK6iLvHlmNcewab0e0Ey4BWQDZJigggiasCZ1BvnatNqGnlJp0YOBzFlxSbjanEto
8+OivNQPMECzstbSy7SKCSxYTVJbTyL2eSfWoOCCn6Z0ekUR7dPGBXpx0Uyen1Azvr1du9nO49Bz
QBkde/InyKEP8E6cpLxQKVg/clVrSAcJF8BQ3BRmoFnBMLdXInT+X6qpujBBLIPrcKCBBJSsdFMz
LoaU4AkbDi3VOhaUdQlw0KlBY+zFzDb5sNqbnzgc55vig/vV73tu3fQvGcziBf06oUZm8WbPkcUj
XMkHWhuwWf72MCwO2yHGknwpeRZtqGFRZVwxTr8knPb8sHHCiKVLNVOmesa3IgsCGN43epG8DASj
w1IuShPTmtvBQeRNUphbguFVWoU2NeZisXXJ+E7316kaUo+gaLqGkvSxJyatMTMRhWy1XAPcrWlu
AFjtz9FUu5JQ1UwumS1ZulEJvY4uM4sJ9nWUQ49PRwwDOg5bsb3uRISJ0JPW8EWwjeEcgU5bulPb
w8Dw1Ia6BTk+BZPErs8GYcSa4VUgYidPfE8kkkQVEStt0wfy3HmcoEa6s7i+p4DPhj0MbeIX+7g8
GgBl7f058+0kiMLkFqn/qz3ZoY+ckT/3GBrDgul0zQl4h0uGG7ZXsId5KM3DZ/NkKRN1Qe++z2Lw
82wwyaFGopSe8CNfpd6zaE/DuD4vb+uNYRg8nAL40BtmgoqM9hSfzRsR/ZkAS4DWmaLVLf7hhzmO
a5mydRcOqUiPjYBxbmmJeFaTbzhoRKCZPAjiLerr9AomK8dak0/X8H3Up9FdH3WlkBPStsE39S4d
PBRQzKrHtDVtGPH1drt4cyLQlyskoIVzHEqOlink2aF7RbJyckoTTQajUpd3M0Z5vOiR3gcmICFZ
gUvWdEC3JF5WM11X+ygj6PNUuukiM7j6G3Il/e0DubqLjIr88WK8WeOCB2ODqArsLObK1INJhACH
MkTOpbm8uWk57S1M9FFVZSf0SKys91X+YzQjzbkTyAb1uUc2SZjUe4VAooIvuunLPPh1q/EeEmHe
C8AZKASXOJR8GRpA5X7M0f4EJyMZYqxaf8VDkzO8QNJKiKLi9mWOJysRfPb8W6X/GpdTQW36r09d
9tge9VKFJ9g9bUcgpMaq6NTi0ZyruRLS0Ia1QNTyySO4SFXgKjD+CbKMIlStl4qlzacQyURKvpcO
bHIHdhs5KRaCYEM56rVV3XwBTL5y7PX0JFSS+wSjT3F3a/eLOd8NQ4e+A3ySBTnriWfoJqq0OtMs
tgqbweQ35ghQGyOhdFrCXDCrF6nQXxREd8Rgd6gogQiUauLO0oSS1G+p2eXWRXEltnpE6kWriAoX
/JXLgngDv1Ind4vQCOjib4HBvJ/8L+yh1UC2CrkgDInAHLFXjzIgPVg1rzW1Vfm5XpM/L3Kocg76
DG92lwZGGpFJcy7MMYX6xAlkJ2LhbMLi1zX2r9SJUzpMa/xHOzwqzVWo1Uj8U7v7iuLAlDOzoEmI
Aov9GP80MnjlPZeYuWgIuwR8QCJRsHLlMm48jeJAVMZY7ga20WZWYHc3i2rbOLV81+opQaf2Y7ov
Y/nGUU7OEdT4QwEiIHlVCjKDH2EI/RnTv3mbRWuKSmTkeZsNLPVrYL4kxiQgzfPgWPsQwh4nifx6
2V0RSDGJGqweuXl3p0Wtk1s+MZ+nEpKHaIAuhFqK6IaoMAkhLEjZn6FFif7qMHa723wfFkNt/BCL
j2JSxpk+td2rKpw1owaCe+G8gOLZiCHqRQiYiIeSudYl7T4YekBhH2M8dJc54csN1HyvvrNyjFWt
vl1doiJu03a+bwdKu5Ml6DqOpFRb4n6VyvnJvLBqi9M8eKkIU0SLtLP6BazvGUKF5e7Y6aZDYsWU
VInEjFGMEBxqGmwl+bQrbXRI5NOrZCnuEDTldO6i+R0ScFmpNa7ii08T2/ePMVlBq8L35SaY4jRL
I1znusU9Ne+3RXq532gmbNQ+gxgumY6TzRRsUHaD73xMWm+KQObB/RmTIrpssIPuXhXldRUq3+VG
rHtsN7M175zPMDKisiO2Fdxq3JiYXO3sMlF7KNiWxvwYpEN7gXWQuCPZW3m9KXIJScLcvE9liaOC
GH3LUHoCB2aFAEgHT+X5NI+QhU8cbdhuUK0Ajty33aj2HplGgUgGz5vKpS8aWsAGpNkj1tl5MrXq
tbYd3C3iffDb+aq/WMk2oghyZjinkBwLY9ltQd8HLgn5dP/j4On+LJ/ttOvmc546FLZb4cbv6b+g
mxId161nXG1zCGYvG4+9hdR8gBRfqzXT8V2Fzi6/Gp4m7WvwpmKvN9BDy8QL1iS7hQLB0ruVjgZ2
ke0ugCOfoPiiQxo+LXVhGNuN6aZNToTaOEJVulsvGfiiSwiTKMUSvOs86NIzLHz2QytQi5Hp3duS
8EUO5y2aFe1bldx3yHB7H4K834QbALFGDzrYY3mFKK0TItHJf8SKwfxQBBFswRBAJdAOWIAkvIWo
RdFtAoutbwO4nv6TK/EZUVN6XJQ2hFMnbPV3XQQtPP5hQ9UREkRUxo4iD4Ksqj+uDI55WD7H5w/m
6/zAmb23qJIQu8u1Qnv/j+jVixBq9tqO2s+Mpj8EXfMOTaKOFTMrkFMKl+ErsV3TlcCSvEGpFtnl
D6srMjKqRXMcuFs/fUvqwLu5U5geoHXpie4zDXIZuO0iULLiCFPJUN7LCPE1flkDQ4uD4l7JDyad
ldDzXDT4lSiN3kCF2TqXmP5W5WtcpMKSffqL9/UC/aZPiR2SOPrwtdBn4ZSocA8QhPyZSGzBpC9Y
eXmKXUQAG39vn1yh8HH/Su7LGydcx4h1pay6MDEmrsGSCNuiC1GW/V2zWW8iR0OTmkL2eSZN3iuA
4el+tl3Y25VZrhRAna4ZdxafVvw4CkE11YZtEN791yiCezWQ+tOpM8496pFm8zC9a28zfr5hPSXJ
7PJbfQcZjPUm6Ae0t1v3G9LMk8owSBxA1Gj8pr3+jitLKKlUN5rd0r7ooO7QMpUWcUoarauD1mw0
lWqiVgyRiI+G1dqXwwBdK7e71UueuIlKRXvMo2BTTnAAi37jcGTMq5DZp3i0KVmXsL8GAf+Odzdr
gi7SCOe9BklB1ZnSY0+oOHjO6BQE/v8mdMpq8bFN2+rwXarR8Eq42wqL6AKpP+aIlyHL9pLLG5Ml
8FdJWOsnbjZnMEBVYNqYCvKLOFyUgy8aIclJVGNeNSPX+OC3egOqpnkONZDGXsoNC3edZ3ecXEKQ
J34kxEmoNyN/T2mDYlvesexzIDOwRfOfHnMLIjDYQ/MfjN3Dym+voTzPBqrcm9Dkm5CJaclsT2Bp
CHicQtakYvtDPbqpp4rZ0xfI/5xCn+KOtXmLGx8dJHoRTFqeJG6eQZXX6ymonPLUv7tu1bFzcPVI
dq3OK7VRKTW/ymWFydZr1PyYK4TGaKMJdMMPXbcIx+/NT4Z7pZc3Tk2/uIxL/gE17dz9xXBQ33WM
9Qke4QIxSb4WcdYt3a8dOvMvpKfmePAjjB+aEgVP3WUtkQuupXYSiYI7opvvsbpSqDu7Ai0adLPF
DFkTQWeISqJMhDOq1ya7K0uCYXXkRGcvoIUOdvjbrKY0J5NDamu8PMT8VQtd3tlCuASgSBzcyJA4
jJiripiMTHz+A6bhYX6Dzi0thLC7W3P04HmoeweLWtTPXgSyd8L4/OA1n5+7t7X15Ws/QSfmtWat
T8B6+vYz06SIaaH0+UC2ILY9nydRJ/KwRje3pQlQpUxs0GD3eAlFBfO1g906BYXUjdeajZhZ3kuo
BJnBTtxVQF2Zbuve13GrPp6ruz3A/dofDZHISc169ffz8M6/oZ8FB1TTHrsXn0vd8+AI18w8ejH1
LFlNeL4IQcwUpIYRgPTwAXrwvtr0AbddWI4fHiceUp99csES4zH6MpSfk6XhXdPvb5OWNwAcDELC
OWkhrO7Sg+bx7zh03+mWbhXGQCYA3WRr7sn9G65EKXq1wvx5KCQPBdCZ33qKIrh+EFsZCgZwgbxK
wcSXsY60BL6U6Q6fZZw8xaj03aEllKdaKLNiCdkN8ccHSKYM4xUu1n/5LdhTGhrBggiv9M7vTblt
GEW4TJJoMvaB9BpTqOxwEX72TXctbqkj7wmzoksIdMVIxOsEqq0aFnvs7mMBham2Q4HafsvXPOrm
ffOq2rZPGb63K8y5BFHdLY6xwln7D5QPcSVW8RztBPoN2niAfRX/c5tEjxELzRlSxC57YY1W0M+C
uY0OPRXg2NMln2y0BA9i+94bnjSxJ0f8BN2ROE8FwB4le/ILN8VRtJ0LwHyrom3Gy0+gCjdgQrin
IsicoZJOI40q6PQ9AmGWWA747/XNi5uSyxl+gEcR4MbLfZvsh8wcBDJTUTx9GSETjxs/sxeJzXWE
f3HETzR8zcK7LQeTpxvwQkaASsIhLuT9DeXH+8bqUH/v+nAZgC093CSbZzGGysVN3CZIlQFATSua
afhEnXBIPltwbQ/hhftItHFSmU8/SRIhEO7lDKl85H5UUNKKu+zhxZnSpaH1RpgFP5LUlOAXiL4G
8nfDgagXSGBGTdjenLSBnOIeble1RQtHbNzX5B23IvIhGwdVQ4VIe0xWz+0y8g8TZatrgdZ8hQIr
GL2+zOexDWP/YDUUKIxbSVqvuGRogw/w59fS9NkmlRhBfnORhBMURP6JE/GruU3Whl9LO95FLIg5
70aXihV6WSldP6FAItuDpBR3r/cveECFFdTCgKXREra4ZXBFWNBAECBmIRN1S3VZPaCMAmT24Zyl
lMo2bFeWw1CARHRlbKzi5f29zmmowBQ/nKiyqq4IM4+VsSCTpwEMb58JgoLbvG3nQRp1suoqX5Ys
/lRUCoPKvhiQjgGNjaDCzGO9DWI/K9ZwX/k17O7OEK+O369LIWcRMCTlBk6n79Mg1ZOi7vU9QYtC
8uRdlbB+pk0SZphKdvTPEeV9qTlSp5jTQGd55QA623Ar9wqWLfIqwoq3CmhosCp/qxwCzeNfdu+o
04Kq4pU20nay9RscKTewZr5qBUBKcYuYFbpp0n7p/Ys493VGthBgQ7V+jvoVt0SxDkW6/6v0m9h+
vpD2f+doTLtETnTyHF6fLjHZioH1DRcnQ+HTRpn4hzI2pEX2mypaMKrRnU70JcrcoC6mZnj4qYm1
0tFKoZQ6GCCacpjqUvTB/VT7hsony4xB4p4ZdznEbOcO/gY8JIIjwXNcwtRfHQcc4fUnZovV10Vq
7sywEeXVM8+KdXuQj/vmcMn0wtc0T/WTbJ+cTJFybLZ136ViJn5n/D5HvM3Ws2wKeOnBPTw/x8eQ
FcoiihLEsOOBoPx4FKYGz1fMA1VAvkx9DhwtaZWMCp6G0Yzx5LkAVjat9CNZHeOn+XYDvX437uTk
XgGG2DPE6h96DFI5ZNHMALEUyWeKf9yOt6HMmAGCtkRwAy2QB8vI+G6ym0Ri7XEECIM7mEVTsr+8
fo7bzd0D6/0gRcSIgJRlN2vOYvnXG1HtjvU+FAfCYkuMHHDNDY+JwxGT5dUr+wpYFCR7XhHZYWZ8
8XGPhXuQuPB07W3G/SjUTih/7+MiRNAfIsTYpYL+Njr3by3RRNAY16WHPqOd/uKGcf/n+AvQC90c
mnr7zxWLrXXRhL6+1P5USaCdcbfF8M0luWy92IWNgz295rwg5QmIkY0QonhbS2o4sxDs+mEmqLAh
dlUC2hpTX48WT19p4+w4utXi0/fIilyaA0PxIz3/Ub7UBUHN+p3Wyp6Ttxx36t5HZveaRlmxfWRQ
iOAexHSKhppXUWcZDgPVL6oeXH2Vp+utCXruB03ZXneydeQMO+1r4jcE8o2nEUH7FLI5meeTL9im
s15oLPFVKKpR5SiPE067PLeiJwngaFTJpgALvUhA6OZIb0XRV8uexxtLKeuCfiiguU1tVTyNHKqh
qk+RZtXkeuZaq6gd8VqP2qFqINzNBCy8WTCDQWZXBmA6CFokwnCgubu5b8nTwmahsA2NuRATdx+T
G/DGuc1BRJWrPZGRBzzGeQxi8uwPTtLrPReVFcxbppnQKgRUcgxBtaFxma3rBueBzMzN2UgeoMqf
cCxUBAgWOYuv5nmBgdid8jvM+l285Ez6h/wQ/lBslWqztuUWHrLNRqdyecm4NTW3PAR6205NGock
sVTqh+M2DBMabWi8psdsmttDumwuxGxVjJ/HXFz0ULPIxvNCb/eNXGLhlgPIYHIfMvo0Odrcp+Ft
ENjpIUs2yK8bPGD2OGayx06mU6OAGetdZWz9kJ3ziykqHCwoKUUOu5ocRIszh3TP2E71eainB+bT
Rgf/rH8ZQ55tHsy3YaSFxekUTZBD0XNVj+l27lUdGCzjGAlEda72XA+sxTYmsygyWTkHVkLs5O5p
eG3pBggePhKkbLj2vIObD5PvDKFQr5gL0fB3Y+WwaHHWjLHuxvIIpwMSe+9crDwGycqTOYB83t3r
IxR0fVQMF1k7nJ08xXC9B8xCGK70dN3Nt7LWnEcXuihnw5Av01xP6PSIZoxwgDxNEmAIWHh5J/+s
TV+EwRLbGs2fmQ2mGBfD+yRB7p9ZAlVo5H7IbQH7UMbriL58/nRJIvCc1O9q3RlV+S3arKxQozmG
+uQCQIVlpD5Rf1YZVfBip5AeD/2OnwGQ+519KhTH1SEKpANmGuvTwiyih0DvDyg/lIOmHgVAmG4Y
pzMweNALBcRXycK1xPO7oLUXyz9y86OpXRQMOpYwy7fqFAx0uQAC1QV4NCGumrFW6kmahemTqqyB
py8/0G1rlBruSePA2lxqAbKgfJtgl5caNE8I2Wb2g5A3pWes+hZKMTRj83vR8vEhusZdVlggH+5s
yNiJsnW7LINMWgKYXFEhJyV+jAlYDhBa+n4YsrBaXe0TX4NB03s3urmLA2oj4WwQ8+FJkDhlnedm
UoKRPLh8mcjhkvstC/kRs6DhU/egrcg2NsA7YhTBXjBFh92Yqzo4AKyvnLVCHwkncR7osypnS67s
c3nlwuSf7lSWVPr18YTrrWhJy4+5DlTvvLfD3jUMoYtLK209FIexzqw7XLZa8Zn7Ed5yqgk+G0m+
bL0l67k8OTvxgPR555p1svdyAjeFdTbtD26D1h5B+HPOZgrZusaCNM2Awj3fOy1KqwvG3MlFZsAC
hVbbB2ezOTu9R+1pUvPAKI+1RR/c1ZwlF2ZauSKGKj1X9VytJUtRQFz5fy/oVpJyka94UUz9CqtW
/KLu3kSbouBFsf9SzRKxuuEeD959Hamp3p9KjRw3HwGhtpzeSRYHdtkHSj1JtMROdXWvX3fCDWlJ
TuUMNfjP1Fy56A7J3ClKq8/WF3fuZRQLnY6HInpA8HBsjfvKdEidRtpn1+21+B8oP5H4k49Blhyv
9WE1JHXOC+gHj0Hg8lANZ36cWACt7HNtGXYNgnHhclfHqJ6DjyXdbaIr5r3rSOFo0YcVX/8De2rk
WuiMK6E7uj/M2DAZE0OwNlML9LtP+3pEeXOTMQu4pA55qUkhQFn39wKb5Nh2ZDnbHiPNfO/TV3dS
dksyPXtUQrVFAebePCwB+feKjvDciDvt36ubWGLRXCr2sXZNmWF8Qz+PzRL98Q2z2ICMQ0bMWQYA
nkCikAGacTYa0iu475uY3zZVnDRedVy0A2qmjMmOQPRiA6E9luA6wCL8Dqi4TQF5uTHajbWxthpE
Hx0SX1Lp0K/Gc3+gbv/IDK/DAyvYutK0vrC7R1bRQvXm8ueOJoGeXShSP3RT1BBPymIGU9eG3Dmk
lLBPD0cc4iM/c7GrinkajKiwAkfkAqWjpxyRRE/ZAFB6YeVsACVVY9pmv1YQ9p3Q6RJoMamIOkXn
p1wzLrMvxJtFNJdyI3xksMMroLmv4BMJijJLUsRlO5ttXYS8JeG2UrSGSX5fYYyUvIJqU51JzIEB
ZgMGBolIguNc7hED9j9CJy5drcplXT9YkVbywnG69vUgSUSBne8WsmOz5tlM8UFpFiVrSVQLddJ/
i0zOjDVWI8Cnq4W6BTGs7ltm/S7Oty5nBu/i19qfI61SnkHftNJDsPDlM8uzByDNzb7bcMlvIBGc
GiHFVaIU9Y6Q1YYJQrNawtOz++mE3DnvmmpHIF9gBHMkc4Lt3t6SvTz/DsEQ+xd5glyzCWNG/jDg
TwSwQ8S3VLq4v9W4MiCOqhlZKIPYnXJtY0ObFM8LVjZNrGE829l5zJ5xmSaxzKMlR5HXHNForrTL
jkyRB1KiDv24STceIB7bnSY+Ai7IjdxtZx0MXFgbNP8ia+lsdATAhc4vAUy1Rl55/WVcHM4LC0Ll
VMdIMlBfmdLuyazFELHh6l2IXRXn96aLm+MRV5H+X6ssenc+IIBsP4ZrxbHX/UsRTu22ba8Be18R
hbObtAp8IzWYybQT45r5euHLUGCCu4MGrtQkD0c31U3jd84BMltFhF17ysj0+lVrM5kZJCnNIUvl
VqdZH0QLwBw27HnIUQwtr+65I2fqa2WilhEtlkwF7OAWGjYwNnVOqhPCHFFjJLwGBm1eNzG+FcNM
5oiYIl/tnx5PyxjHKzpWdFKC9iYyUoGdrfcUnSz4MNseGcCnBdQ37GWwvAYYsDWA7NDQF9JtboMf
eowSGma6Vwu2qAK+/XPNaGQyaWokQboyDXdjjcAYqYsBDU/JvJQ+qnKyhpFsJYPV6D+gbwhGeb2H
yuE4tNSQVcVwDPdJBYGcugDZUNTiPR4n1vBQYcBSN1NRk/DYR304d34eQyjakWWaMmdnhEIszZuT
HP1asV2/ZDTH9YIFa2DsndRgPjsk2WWhEYFbXY5GGa8dSEQxBtnrV1vlY5zQsKbKomA9UMFiG7xE
auw628nPTXB2l8Cx9BYbSQznByvVTg1ui2IvS2vMBB3d7bjEjMLDMZ2sDW/kA8qTqq4SuFET/tDN
Xw4aGXkGwbG1L/U/dafnltaU9/EvoAnEHl5huzN51T6D/LYe1xeWmcO/bjP0JryV1V3s1giwcA4l
31/Pz/LFCsY4TFSyXSDCFAUjoEjDOj5+VGTWj+L8IHA2BDxOyVNFZjhfdEbK9Is/imCTSlymxlvZ
WiuFKzo0WN6nHYXoXMlNvZQwcqu1ujFXzIeoCU+VHoQ4pK1t33RCVR3xn6x5yOyA/3cFEbFDFZc9
2V9aao++jfo3qvP4AZCJuWmKWLXrf8hp8NrjC0GF9MRBjFgjGuoHsD/FqCaB+MzB5LLiMtgBKWkZ
3tnXXz6SWUHdaqygT0fYmaqDRXRL5MDn01fvW2r1iMuQMhRN66hZH4Hb2YhJlkwnF30KUCRQvDmZ
BFFLKv6kzkiPnYFKpbTDnVmEz7VmC/7LSr6JGCUuV1EWB/86qxkaecob1piT3oQb4xs7i6xN9N88
+iaimor6s3vUF5LdUc9aNDqiSP0lAHNRm8bxwEVHGazWgyY5hbKmedFz9rpJ1F16neG+P0Qwx7cb
OiqXZTSCSTiCU/Jrm2qEy55lAvUsy/sXimSPu9zJaR+f5JbXno/6y/dDQXB+DPnC7mfutSBiJgVi
HhyMvsYPNOIuXFqjTULOP+zr3ZybC+ANZT3j5rBVJVB3lHx/febVLu75QUpLsbtx66iaweizEO9S
URlWZJS8DZKVAt4ZAyLUs7JeK/am03S8qdgAFF95iDWbNH6Vlq2xzw6rMx2wxv6GbOZxKBqaifoI
sxEoVLbMZNYf8x9OOLPkWC0SHYBMxSV6fuGIZFspaYBMehyckdcB13m9GhglX0FQBTa4bJc5V7tm
hle62uUkgkIy68Jyh1CgY4od+GofX2BbFXI4R6fNAGoFoxo09vgPITUmSZghE6dT8Y2qUIPr6EBv
z3OOvsy5q8Je792J+wDht7wOwOSkYsWFRqRrGqDdhEvUPfCvTwOfnLWF8bKRqBy8Z0MbN8gaqHiT
HYKgW5DAZ4uInlGfbzotzoKFSqEVv47AhiXZsgO5qMQ6oT2n3bv7u56ypNtSIspRzGX/3pEpd4zW
TaOc5v3FEo8Rh7+3Z00RTVvr4P68j/JaGTN8vUTf+MhRsQWwEIPHo6nPwXK3EiSrq7ksliNPiGaR
2x2Ft+wRwuov0AARys12HnT6FA126M8vhfnI442+aD009ehoHf/oqKnndPfWPY8groG2Mx2cwLRb
j/8F/jHK8PIDeIdB/YUftUAFZl0h7OaE3fjLxS8F2s4PMT82VLxfclOt10p0rv63nkVeiXODHsuZ
waimrvTvAR3Dml2z2ollUK09ItyvIzvXra/doPNArglsYvvCS/p238h6gtkkARA6gG8b7csifJTv
DII8EZrhnhbmEQrRplFUFlN3nwfmb9dMD0PmPZ6LOjj0HwYXZ9IjLwO13nHD61g4t2rnwUvJGDuJ
/G9fn8C1u7GzEBzgHROOznvdwkKCnzSkH5OLjmqOMShVbqezlcVvycnuIGKBksesG3tYzlIe0a91
QEBzVVF8D6iE14CO94m3fmIUB52kxl8W11A+rzjzugin2Gu13D83CdZhypYNkGMydO9QorCtYXKJ
Wup/HVxlD7BROdjJX6gwrsqyhFbpsLoRV2Aq1Phcu8KbO989DrOUlt37+KpTK1up85Zs276HMrFA
fxrh/VrsPHfH/wgBwp4dmXkp7hnOROhofnYllgOm9JZjrGnJ9D72v0D5tW5nJS1t/gWacdXTDJ7H
L2m+qkvMBHiQ+c/A2ONGc301f7vJDE7nOYB/ftD76dsGfJdCtz1OVAAJv+ZCADkzakxwJDnYrbmc
g1HA90WKkqaSCLUT3VA1Ga2h1xWYRLzoT/IeMskS9bVB8kSYEffrhgxk3EnDhOgbwWksWbtZs2Ct
/IT1JyAmoTsSTvM9bj7QoJhQca5S96jp5/g6xuwwlp1JykHm0CBMLcCPod1l99F/JmOch8dIoDnS
duoJoSecptoLnKnOW39Zucl/ctL3FQhP/sMXxNW0iR3+ljoEvLwV0pRrJ3hVLjFk7HJYCUVSC986
wQuHO6ihXvlb/EjHtd4k6/UCVKlf7kJ5aN5kzd0C6mVO8aLmaM367+GAo1/GGbjovw+/5f2hR781
0mN3Ut6qZTlxViJGOK2wZsbsCMAqU62G41E/7u8G/oYM/YMte6g7+fkufPxHVvqPQI6oky2l15Q4
CTJKhccpaJgJsUUja3k1qakRyMSEpg6nhGwgcQSCPCFKNZ+5ksNLHZMkvywpLDDv8/XV7B4zu2JU
9fWp/ivb4BqcHZ1mL4ScLb044rPBcHPIw1jZhiPxOdJcN3IXXbu+2+IQ3PAaTVinLZxXULkpVMZN
3jLMxnrjyYysczZWwELBV8fKCnogTaRV93F76z5PcJb4I0i9O7RsrfMMuoMOvkyOxkGgeQ1STicW
XSWgD/1bVNcnxE3f7Vh0Erjji7ekKGeXpS9yLLbb4JapX8NVBa33ACGqLGgBejXL/H/AvUok7+TT
2YW3RKEw7pb9psS6ZlCBkozzDKGPVNxWgvKX/v9soLHgCdzUyChegx8XiMTboF9dLT3DtfbSI3vy
GJ4W6rWpv2cLfKBMBARPUdyFm7hSpeWz2peN8+Qw3+beXC88UyQPktagWcObzWcZszLMvzD3ehm0
4rEA9Y4KSqeVrtNCR9IM+2PHlV2LbJQqwTH8qtasNcCYQv7lihN+gh1xR1vQbl7ahVhsOZDdMv8R
iOTVY00slVBscGuUFjreZCoQE/Mgf++3FkJQgttv2Hks1sc3ZtPH82s+4j9B+vrEkp99sDA/au9W
QQMXsQdwtr+Tf1SpybfDQ6dsVTKyhImSaIPIzbFmmCt5elFwz4HSiMFb+pVuFncqf41Q5qyUECAq
bCAQ8l42HpRWGAFyS4aVpQAcqC7V+/v7GQlLPP1pUqwsoWixmTe1qOR0zqdK7xIS4a2mM8NoMcTL
gsc/3N0IzQvC43QC9rnh8OTWP8cOVa0Z9dAFjn3q1XY++CV9Y1Bn2EL2fff1FcnI89YjdsigvrZ4
cE/kMWtYO/UnhckSLG4XuYg5yhSTIsMk+p+sSieHrFdUssBKWcOpbTUjPY7ENNfojvY5e35GYVSt
+T658V+IbalZPYlGQRmYUGuK8rbRsnVapfZYPWrjaASgEyKc7LalDovJLxDc8x7pqzawMENN8cND
a2ays1bVl1ufxJ1/awO03UUssKgdFdVSbJ2URU3284kZxsBVQhghBV8RCyUx/0VLR8ixXARmc0Ng
1IS+crdnSdXeAkwuxy5d2ETb0cqBfN4oY4Vu4VB6ji7Y8/F66bcn6xOm7n/XmL5RoIdnr02UY2zq
/+X9GMw2p7j/YyV53QqOa6+p6LW3zgi7qULvHGk7+xGFnEWdrzvGP40Nm/IzCW09Di1BrYWdeXLe
GEY8sUSQejg2R1ArKkExYyjGgUVG/QXGxY+v9glcaTHpL2PoxDkvoG6hW2QPNCf9F9XakXKZYKsH
B9CuiE0xpmC6ntfvOf73dK2SSlQnwdlMG71fFmaJjPahfClNY0kDm1FpyISXNPR4XQCUFxSHZhVQ
ja0Pz/goqyYL81D6bYICRskZ5VojF5ks6LEqUGb8tbjUTaYPnZNgvko/104n0JbM/+DxRyHtjezN
m05bsq50r7v/AinoiiBIi3LRU2oxIeABJhvy/FaQIThM3BE22tOHOz9e2qWFh9O2U2MXZW2O2HPb
vmk5xm8d/3v+Ztp59AyIJtQXDYVMXMH6rsNmpyAhUDt10Kvx3n5gkfSsMAX1VI+dmrM7T1QNkApI
P7fyhudrDh7PO6qU6rLCGLrm9givAxg1h8e0W/5EGmufR+uWSIXQ4I2CrPp6u3gwEQcYC/nA17OD
fq7LxtBJktQ7JQW0p4f//7aX+4yfGAL+g3qtYpMlXnMQWulg6fPHd85VuxHusCxx9GU2p75ShZ8l
dDJgTtAU5YVmGAfJRsJ/kQ3bxJ+bp9lEWHZ4lolXBl5H5Jwhcy5CK1+W9s1VE9TLUUdbeF3KBbTu
6MDTnyc0tA/S38uoiuP9eAiMVcgia0ealjzOqUKEAw0n/c5JReusOTaX5GA/gnTyjRE1T9FEwEUt
9wZu8v/x75dLzEDIfxmrq9h7PTk7IcmtfC48V2dNZ08EsNbTu2VcndfeOSlQ9Fk7/bk6gLg3ERqY
GsJ6Cv1kvufBrmAXTIY0FJ2y0cXRaNXGGv/nzWXZi/B0pO2CIuu+rceQVXBkpfTk0ZGuD5BEiVXa
LJ28BK8tvnZo46MG4AcC2F8jmnnvMGguisRv47AQdeShWD+x1K7LvPMD/RAQJlC4lgjf7IpfHYSB
p4dmSaEl+FAmOTcomM438AhWgIlQ/X9pSwoy6RSV5iMA8zgMmCrpJFH3SmuO62FVLXOUSraovcFM
tTSG+CBoPkEfGSVmsPTFVtAkI+MJtmUCORH9/rs5Bm3EInJbBe+WQGq4GZjx4HGqwtmLLuektP3g
Cjw1CPEgszR5xaIpC0w2MfAg7XPivIhK9HlowAXfXA63XT0BdFVJtA33/HrUEU93UL6GCvRIbivu
XbacrXwFh+DibWFCGWl5gn0ImOeVp/Ablq+h08n8/Oir7EnCTGjR74KWKsJy9a/lha0a4lAQ8mrd
pyP3kZTrrMVWpvNk3B9mVMDm6U8j2dkOMwBb2Q3veg4eAu7/pjIkSiRMxX8yAoLZ9OBmeoCSug+C
Eb22FrTO5bMeCVlTxw+eTCvJslAR5e75bDH5y0KxBqZC2OaBntb1vS4M2Z3GNMOZzMXzHNysuDHD
S992UKTXwIAliuOFQLADD74UzgOxeqdJ8rsq0CEYgoiuLuaEL02boNKHNwFam7QSYrDAQqymuLmv
AG3ONzSO8mtbxt4bJ4z8NJYIR1hHeJHHWixynSmm2Fw1/7C40CguOWx9o78fHYrzL4EM1P7xgi80
Wf1d9qNrVeC209MWQruL4QvyeGDC2KrZUCNjx8X4fWPuZkkOhFP4Bp/c6pCEv9WMwqIzuY8iUSS3
lm880UGfQ9jkPlCVC9iRX+Iqj8S3gj5quDrRd4r5WjIn7GgEAxJhQyADtnlfewtWZ08lHqXijfCU
TCHIBFDHFCa45Ce2O8C4bqv/fNOOFbwYzeNcIeQyU4gZD7NZ4A7iiIQVfgmej3YD+t/+TxCbWXpW
Eti/r2HTRkxlasPxkVkcHwnNu7ZbIL2MkE6SILD/jb+/5YNo+qjgOIh22ZXtB4cW6wWuFKCPFfbp
mYJ6yaqHohUpmKnztwEyHnJyokSZCGV27L3Q6ilCE7t5K1Yk0UkpyjNcvsajp5/k+8XPYssnFgO/
AYFNR5TKTfM1/DDxo8MZsH6ILhj/TwpwZSvqZqLnm2kUUqw8FqdLUDGmLJrXTduwk/0IpIVtOFTH
XuNy4iRmFawrwX8/y2BM216uOyP5Kp+jTsKD1+E+ncLbU9fT4FpLEsZmf55LDjNc9YkyjbWYpl3I
TO0vD1Y6ZsczFzeXNewRhGrpUyu9caytKwbQHJm4LhcNSpaqLfjj1+qJIcC8KncNr3bgG7ETFzKS
IxuKdmWIn6dCINyyWFcLUna63vbYKsBmPcu6EMhRWoxYPNYaazM+VZz0x7k2A3wfDtKXF2xBUJhw
M2n0V+LMrIE7A00IcTAkuT3Qo4ujlubwrrOTeyZXqYj2Z1KznBIJ0a9Arc1j+Lib54QGXK3Z5oog
9JTHbMkXNwZYotW3VfwacLmjTED2MBxyspjBW9A/pa+domnmW+3YEptPlCPGjLOV9sbLfc/HX7s6
Ck4yTxT74eGz6IJIjfZZNlPdjVPnxjbGxpIoDh5DBomQ+4a+SaaKil0robghGW1jnZsAse+qes6Z
TzRtW+/i+vk7VdEzsExwBTKZXqhAixoOZyyImO0qg6wjaiGO1Naen6nxcKS2UcLFVWw/lsMAT79B
JPEYv+9txvchwNSbulq6wKn/OLJnOKkjs71O6aezdZ1WBqhfZnLLnGbJGtBIrPoWnHcGhlOdgN6Q
EMO5CyeAb41jGtoziNk0+X6mIg5/551P3tsKx53H3hvzBhpY1SiZuwvd5Pv3IlleLpAJE24nW0KF
rVn6VvilJsH4E/LBrTibUFkkOrVHg8L9i2H7enAWP0TjfGHnnIOEdGSdDrmGLedDHODFR6z3AYyN
tD82GH9UnRymWNrc5+AoNFTxdzG9pDVpGwJa2bS2Y4zA5GQ1k90exOVdKWmebBWOFp+zdEY3kJrn
SjYk9A9005nc3iXb022/MN5gflQyg+jHAlF7k9sEPndzMoL9AmOGM/n0QdDm3IQop5sD8OWkGAzL
TjbQm9qEJllodmVI7awem/1/3eoZhAUNLBAEusNrWJ8ewkVbj7uDmbaPjXbGTM9SfeYOoRtdo+fT
BtxBURzqvCS5y0u0wAE77nq0nLJpeRrMnhotm4Cwts2Qp3gYNjqqkSnWsJSTrYGhwFXB+dtOug7A
/31nNcaWTOGHAvBctcNdSPlJxOlPx6XQVhWeVHK4KeQRGXcrsG+Xw1QUCsHJdRDxYNlCWZIylQ2r
Gypw+Hq0UCII6/RSYEicLyVBy/6EqasfLE49xH3v9+Y1vZN1b4MDTEZ1+3As+rAjgp1dqFSzaKDh
k2uPe+JXYOL7iLwfZ6XWA9B1eeMyE59cGmn26gWKGgKhAzy1d0UAGlDdanduDwIjA7AdCjgacNzV
OoUAkSmt3y7Ol/tglEMJlm7kmLoGU2DQcK4S7ZqfSjVAWwKneBWeXvDV0/vu5IDG/w6fDuWd5tTV
E+hu+SVfshrliY2jLKDS+d3qBc9jY2PZne0r0RSPexFPYNvEffVfBAhtMMrBhAAken6QNCjnRsIM
AkYR3rKozBZUKHZ+kl/E0vCUq7h/xK+DZny+EpWGnpAIb6Jjh3GDUKFlpYz6+XBbkUmjqREkOh8E
tJ+He7tD+CWP0BFFQ8NazoVvTpyBVzXQiWg7tY7aDEqm11AaowWdbWMyFwGhvndX/lZDduz0+gXB
5DNx3UYUO4KL1N0QOde+wks1TqR2D5dErkzB3znPkfF5/EzIowCI2KFJWsblfrmftZ3s4eBqxAlo
ymdR3rQV7b7QzK24pcvNKr+p8aYP2al8WpfVn4wCk1v6m2GUrinPYpG6mTCuLGfn49FrvGtaL60v
3wKH2PxFDmltIEfRzfKJdGxBFhUtjI9xxPjxxraI3O3oYFQfiA9eE3AjbEeaxCxp4ChdwtYtsI1q
MMiRJiS+Tz2/HcisNKnmoW6tKhckULGtzx0hCJ8D5y6jxAEmFhCjKl7GOBCG+W2mAOHoyxfaeomW
meAjHU7RJ1u25qYJcFnBaXA0uiwCqPFBUhs/rGN0MQ4fMzl4NFJZNuAB8oKdPexjSYnQEgDOIcNf
rclIS3c8dG5GnImGlzoBhaNjhYsmIejqttw19aWrBBnQv/Sf7WtCf1NOOic/Oz1Ws4CbbR624G1K
M3yGZrOOX0yoMWYz4cIhwYRUnuAemhxR9FHKakinCim+j5kghYCIIMu9CsXonqTTBGSzxJ1/+5RN
ZEzbJSJUKNrQ+Wd8Xlg1PkxEKitimexBYLJ8ZvU0c27e068QmNre/4jLpwcycj4Ll9iv/DH4UU51
QejrPAYq277RJ9WI6BmzO4OJhURdSzweiU+1Y/fbXZEhxLUz6knT4nM+GHyBStC4KnUHMMRKfprZ
6LxIZk5iKG1EfqTWooyQVVGfskKjpyIyBL6oGvoweB3v4tmW8Ro9wpmRjICtHvwBtMmGlxEu0RIo
dAyk6CqCUdc+sdXUMnx5Yp/QpSMuJ4GE+ENKrlasCa5WOjqFC4S9WSjB4IvfP2/5s5F3GjeScKaK
lvhhqb/tPmhUIxaLiOrblXlHqE8/MpWr0JDF1qJWhfZJPqVcvBeAuUM4EaCc3UNFzaIC5iaDpMXQ
qpfxwlEYgQXdNSnzorcsDWqnzTrXISSOEKD3C6MKavI82PqNOCYbHSemiEOG+iujCrP7PahSDb8N
UEQhZ6Lkc20dwpwIIfSqCPDuKvIep6rU+MKAkxlOyQGtgOgxHN6klA/6063r3paOuLieICOyspLJ
JpaJHP9kVvF6kyulAX3MFIBXrlSoneDi61KF+VFiyd2vK8L1UEPp4RMd+G4T5FKxLoEQUx1nHnV2
2UngwPzhchPAJmQDxWE9o52mDFYGfosHgSZ8cM6ZzR6/CgzP+xvMuPMWLCpAcFiaJ8G736PZj0qd
Xo09eRUA1TBiplaCuQklGh4fnxyONNhNEdROB57lsqNulloZcHX0Yi8G8OZ1sbQUvjzKm622AD2V
w0vTy8o5HffxTENDvqU8kBBSilshKXMzceuR9NJb4HmHOHW8hlZNtpssL9aAo8ntR9BBQZWKiORn
+XJrb5Pu31nBeWUK/Ok/b0Akjm59aI1r+m3AI1rBJxJ5pt/gqv21VUB7OnH2vKaQR1VHSt/4vXmW
E1Q1zdrhnMWPe9+lzEBYJqW0q3cO+MsUF8lNsnLI8sx8N03VM6K4zu/W+kTw8kWXRHFWgnbU2nD4
pCQaiLsVkCSsoSPel3XDcn5AwbDolxw9ksM00OM7lz4l+YlVTkoWPkMA6glPPctnvwxSeI919EAC
1i63pSGI9WTO4pGgdlEP8uGR3j3RXJj9BC17NTn8cqBHWKzKO7tYEb9hVOS3Ch6aCZadIrV//OYC
uRkcLpoj3A8MFR1AQPUvSzrG1/GKLBs2hm8H06ZYF2IR9z0CogoXfHcwVRB+t8Scmdmo4sgsqZ5N
IYHkB/vEFLKsq7JnJd8SlpWcAgOwcdy9L5kMTeIbWzNgfz4MgXWxSeaEKVl6vtRR8Hx7UmQ1kzwI
GNgQMmdZOlhH5E7aCeToQuBdf0rmcJTdbqfbxkGdo81cDS77sshlYAQ081YenTCLwwDjGCXJwfgI
s96mMEFHJ48zo/O/Z3jo1xeYbtgRMuZTQSgXg3lL1wNIC2nbsUP40NJrpFxGrbzBoWlByoOitCnu
3H9v8s6lYp7xF7xlJbzexGjOvGFlO+nKM3ocMUhCsUmwIViLruYRYu6WoND2iceACCkBZjjHL7Rm
vHQ/5ccitCeMROe6zN54sBgJKfXO9GXflR26xl88wNWRckMIlR8v0ATgXlBe2MyRQrVEU7PdP5L3
w85wmmlRK9fVneyXsg2BE7VlvkQDRXSw2DnPXxHLHcaLNBa2YSIUCmNRblTCqjoI7uSM5Z/xbq9X
12VBBMWcDmKJp4ddSPD1/yGPWrVR6Rckdr8L0eLPTN5pk67rxZkL/QN4brjG7foombokgCFYDvRX
YAr4NNS3hZtJc1x+j/9W0fBBUVy6XYiwYz7+YWr4/QKCw5O3Z+mW8e9KfIbhyUL7lDiymxFMYAlN
pb+X3F9DOGiNmIQ5G4GrYuAvkHpdNZNeZoKeB6mpQN+v38ryTm4VXudhb1zCTlI7AQVR9sQr6PGY
Sm15qvZhXf3+6MS2rmPcxJNFuDUecdh3f+IsW6tlpbwl7gY5L+TNPQYeDWq0HGywZS406kqqE72l
uBv1djQmLhQEEUxL87OBCpLl5pk1Jc5d9GRvLbBsjx9ma9sSQwx1Rud19SBuaEiGQ5m7EL2xqpi5
IeB2bdjQIbSTcZdi7wGg/yf/lCpSjh57EJukZCWDG1UkVP9D2/J3D9lmOC5RYup5GYV3CYjMii4+
hYD+welrWnVAvbYM9yV5harPcv1gIZnww1v8K0RSSngX/zt6+L4FykDd8U2a1MPzZ1V305oJyesC
9KXTYqFlRHSkLV+f9vH5ywmVj5fNksNXKVShdtytrX4+mUPtpE27zgEOVr72FCIdO1hf737DnvYE
bGHVtJ1Yn1Nfpm1cgUJtIE9pBkS9FPSEeyTHXXL0b4jTvMGO1yRmFG2d9USUcwOQw3M7jNum4pmg
O+m5NVgIAiC4IeQyhyUzfu42E9eVUv9rrWOyyndp1Ye9eBadpsLUMY5RFprjalXPUyP6Yn4vycuz
e932Cee3JxEFJg5gcZHJ5PUQLxyP8q2rMORu+qM5ViU7zb4ipMQpQZDx9gsh3bOXKJIluqUxniPA
5JKfuJTCVw/pXfTywdM3ACu5KKYXTzeEGblUmwhmNtSXRTnSuXwufdqo4IGghvvQXPUzytbqXBRT
EWpnZ6FrUmd17uDcy/G7biXl4uGUo8NgC1fBi2xf6WqrElO2UROaDV3gw9YDnPu5eznO5LxSBc1o
jPWxW+xYEzzNRf7hKq75VXuLzQiRn48ghTjZDHZWVggrz87UTPG3PvhmU0CiKDyVA/0FXLkb3WBS
T14v0REDoKo64Y0AcBfkKGDGZi+C1n+025fBt6h2ku1BNiGYh9VVN+1yrLX1aPl2BdaGVvRSWpcR
6Fyq/AOl9MiBt5g3/qfh0rng+g4Kmg6FBuqvQhUABWjOJM2FhR+3R5UHH3TA9++2B8D9sUwFthXY
9thIyXXwt3WwguCeXA1Ld5PlOvqPDNyW06Um7Lux4zMRQKhc7iB+FW8vmo5YHPuYbG2dTPayeTkU
aQOH2KUgTYMQDQQoxAdZz9EbJLtL+H7VayWJ2/A2VYdaxVEQ8W9BiT77pOJRtWAPaBGkXBPYCPRG
yMhH6c5q0Y8ePYycxmxUu3jeUylLmjdJBswnydijT0e3x21LhdOa4fiQlBwoJhUhQCJ4s/72rmaL
BbGoJBJJ03t9eCZDS4+YAsknWH20tetEWMwhwoj8b4UXYrEHqtP+vqSVpQO5g1QDHxQsIkP0D93q
7H7ld2ayltBztbHxRNsGOxTXwNaqNrJ48qm8VnzZjyek2qKqutpSqNsrSrusw3oudXpb8CiFo9bo
g8bHosTzIekujcZQP3O/025EvtNnBUUpZFnVG2pUpepz840UNfz9F+zoQ2y3fMTdrntyCUbXG1u7
kY+GBxZ2BIR8P6wLMaGzDs4xYEsM+sAisx4JIqGrwYbF6Eq63SrWP1UptRogD730AUm3N4nB5FSk
4HtXIIYLyZi6pz3S2cE4dknO5Vjz+zFH0jrsmkig68MnpHydyzEycaxc13aS+ELxeOyWk8JCcYN3
KnOxM4z/R0cTO3Xl/QV2JDyRvjsnQPSP2H95PWxTDslp9bCRbKceWBHpgJwWqbCB5FEJUlDX2m7V
pxWObtjfTJACwqhiPbimBEMTexRxoi8HhE8SMXVKWoLJqx03xHvEYF9D9JW8FKuo/TZV7T6PAkw9
+9jZWys9WFXjtMngVbt4evckfHPcK9Kwt+uXnRjT3z8DCbmWKxjK6d55qAtlXr28+bhWWrjeUUO5
IH8lfxLxCl1nNqj/5gKS+GXRPa5EUzw/P6gIVeAoPc+ilfKTsG+QWKAhW4zgPw4jsQGLNlGvBE2l
WDbR1GtrWUOhHvBGaWwtVKdWKlY2Ns11Ig9UGqv88qk3fJB/ERHDjEbCRM+uz5mg03LpZ7NYFSnK
NFhH/lHGsTWlbvhlj0Ypa1+7ch3ich9CqHMxKpufqXhAPfbabg710X8Xz2xXg4astRIK86ydHygG
zTxOlEex3ydygDoCFrCCwS+AJ/pjKFl7NsRwqpGbKEJxuZKlOh4GIV/J5MtqKvpqKTXXgV+BggNR
YJFiLcohZMAfhKxEzgxzSf75YYLbGGTlgtP8F8LMALYMKJJEQ/CkaNZC24P1HtZWyClPZmyYQwVh
M6Wt5eaV/GJTXxpdekwE8p81WBQNIq9cAo9EWaOlcHpc3iHVi1HVyiJw55PThtwhlQYO9nfH8LHq
nyXWzzDH75/vF98z1YH/uSehpt6hS2bLNZ+1XWMXIwzQhoFqf4bM6OxrOJ21xYanvSs/okAFdNGe
FMcIKLteEQ87vG5WKDyn9L3R4yvUXoE3N9uQG8sI0iFr1jw4BjfFVZHMcv8lKEKC4H2/EtVEVmb+
iUJWR1Oft1nS/wY0KnhqNU+TcQUdq5W/0bMEi13bMKDhUVCBHn95PBwYOY0rht9sjrDv6iR+AZnX
iQZh3jr/zzKD5vh7Bk8M6q9jAXIx9os5t+sg03fG+ZTt1AH1sAi4e2RKmZC7FGqXvBLM16I/RHYv
r4wqp2MNHrjDChq36K9+GmKRVr89Qzf+QUnPTQ5uepxnjfujPyPTf1zNhvdXCMxQLLpDnCYVw28U
plMG2JEjj+WjXvie4EXcJKcGTLfXMx6vSABf453vLkLKJNp9dp9eDdep7q6VbiowNCqqeOtvpYYf
ZZsRltTmwJ0Cn003Lsj8wJe55cSIYi6d+Qm5jvHq3Pw4SrwjtVkU+tKR1KC2YLKM1K98jtXnBcdM
6Mv36V9nCjkvUh2Phtxkm6G5Fd9hONOXRr3XaoTtUKD/s2IhklvsANgkswt4SWQ8vOsIumjTfUGS
hClVrFtBGXuBoLcfbK1z+4j6AsHdl4C0dx0WR6ppN06Il/t/1TXEgQQVwPdvf03+Gz5PhnbkKjA+
V/McB9Mfpxl2lDg2yh5D0bk2SiEvl1B55UyzuxUf9XYFzmKuldTWc/chJp1b0tdNnHgufzcu284D
UhDmhQItWOXH/bAcWkJhHBzHaX+BTMuaLJK71+gRUiqPeZqSRb8kFXCOQZLnurtfF1lB0KrN6Ul6
MKLQ3UjGzWswW17NmzDEawNGt8QM/1F75yQ/6KoA4IPWmehDOrRpUrKDoZDu5vOJSkgmoJkYXnrB
Z5Qn5R9wiFShQU+sXfjpF9x5mZXhUtQkybUcHjPLfWL6Cv6xAe1GNoi2JZfyn4yLe3qX26rEhZMW
1dTihygWtU/Cee6IrH9fDsbkO0AxeOc/lc8dYS7LX2dQc5Gz0Ru+imUVcxuP3f7tlsIDcJ9x0j6o
ATm6SbALZi5Funkemr0TLSWne6JOvfyKUEXqPq54C5hS3K96XF9yZg+eqqDm3mO7TDqiNa3sWHVo
avb5u9XlnSMHzPxI+O20ejkH4JbVZbwkw5WI3oc9OVdJHNweH7kK+rQZIxLB3hsD2fdq+oYR2OGu
UYHNKy6tSrMrAiG8cYdxM1YH/9RD/QkEkKq4eP59ERctIaUfuv3zJie5OOd7wSvkpJUEignOl/fB
Re7BVjRxZWmv49IckSHkLWrSJN4IGQ1b8eJXrL0rjw67KNsu8yRCFg2ciNgTqMKllun2DLMOPpSP
NguN1MKgwYEoWTDMq4Ldvx/rnC+rw7hfRjxGX71vQ9WOhi0L9PNyhAC18fIHTSam+qrmjfnkRzj+
rIou4/ImJFrlfcJ9Kx3pIDEo7HayHI2RLbYF0k3Fk5yaMFN34l5g+h1z83fm6MtWhf11/xAg0QlS
/J0UwjguMas6HZ8VKrT3IEnIqfVi7Sko+gNlCdevrTx1AwhCKxMlnCYct0i0HtSwLlT3dFeRPTtH
DjdzhSZWvNiO6FJIH5hmdiNfm1Lwtt4sPkT3U6Ey0TMjzU/FZpCkQtDJvcZzVyjfeiaVxE7DBbV8
WMvLyV/HvtLIa8RDhMjRVtiVoqAzgjrigjJVDU7g/FOqa0t3phrMA4532b/ukYBp2JJMwvL5geWU
OFFh4oCKSNxx/qpVEXe+f2KnJ3LYIeT4dDPphQcYO+FbgvenPJMZnzV3y0neetJZfYnByzHJK0tU
88/cuUvlyv6E+lkNEUw/81m5yL+3ddcslskV8N4M9U09nojGwvyuXwWZ8mmfywa+XnuK+8IwhZZq
baz+9iZ3f3gS4fdvaa41xDom89nbLPYxf4gWlfpTBI6388b6SMSJ79T77UvmiBFucKg53K0ElGw3
TSHP1oK+K0ldK61qfKOa+0ooQfjMaijq/1LuB3SWDhC0CwUznkCEKgaZbxfYgIJyWQ6HB7I8Iy2e
7Yef8Tql4ouGMPiEWnup4jv4F4156s9QNCOKR08AJMFUq8ZSh2vaAdEZ551M6K4Z0B+PrGNBrwCB
2NQcl+CNKcfFTi6wYtfBHIMD+RWsYZZqzUNBXGJmjh1fNNH/5I7FeNIQwfOuNB48tvYNc+sRhsX0
VEzK6Kx12/EaWNK2L0upQn29jw8OeeGPBxD2hBHzqNgqs4Wk2PzuJBsRQV0Z0z4CbkZyjM/X837T
LjDxOi13zI/b5v33lanf/1bbQcvIoAwMgZxnBrvuX2PRWAtPJQ5YdnAb3P9uoXFfCmOWMXonACSD
FqkZWLZfuR1KtrAnZ30uDz7IPpFb5vR6yEmncwi4zfO46cvtXWcNm68SLW1Jef2ij8n5uddTkbO8
YLyQ383x7KM8IAU7ew1ce4KO/ggCgpGLah6y196A7waVzeTYyEtFtxtgBv1YxkCbenqhBmaxu2oO
Rml51IOhXfOsJGk8+2Ep3n45Gj6hV3Z3NmZSRypJsgkKkmpMkSDUITM5cYwwkaqDVaqUs7qErPNi
huYM73zft7XyAg12/pHrlcRxe5RatvHFkPN4jpKkvDhbGBOjdaTQRZasLcXp0Z28Pi8dGF5qn4Ci
wF51FFnrUp6vTVYYCq/tqsDneahlmNkcV1WV6pd9B39uW7n+4VEbqJqxngeoYO+x/PmjsQsFZgz9
pTXoi/9krG5wlhFcbDY0vi9YhkjBfwvm7FQne7iwL3W+L+XZVtcUJUO48AQUj3p85fv9oeEY3Bf3
qca9dFNaeqI0xewGE9mbruMjTT50yrMtiKHf1xR1ABhqVMnwm41kVTwKet0t0GagwxrHHB1/ZEPR
f3XLtmQguwofr/YVh68BimZTWSHtXf5HBSUOU1fmUsCwZb/I3gmaSK9D81RbdytHFxZMGr+9upLN
JDckSOUieFnBnRLt0YqnYd5LyuGNTQWRLk8xY2+f6MMtpI0t7dLU5zMZcSnyVHnoEm/5sYGzfelg
GWayEy2rH1rPnV/G9WFRoXzwwP5jLG9cQ++v9Ge3FqRjKpDr7Ml3ldxsjvziYFJ2FKjQUEJKUPa7
a2GVhBVIA4KBkStd4TBOBcvCFhlhIjkfP9q4D9p1dfKAI3KtgmAnqk1qySDJvaqaf5emuQXEL3xS
JXN+/hEYLWUkropgzk/tfl3KJq63Uiz8hFwt6rnNlr1a6Gjccw7icIUb2zo66IewApT1flwBXx3q
/mGwv8UpWdR3ERyOIWwVN8tlXusJVOd51nffLmXXHH1sz9zj5yGh08D5+ToB53gHmQHIUEgwXhBt
6v+EZJ+QmcFmEOkROSR+VXzDgS9gj1wZcpMCm1x/ydskphB4ap2MavkJzNIKRlTZcGCRjfxmY+Ai
JB5taNwB4dugalwnZ5ILJKxAqigmfEa7Fn2ZXpc0mH8X+528fAsF4CZACU09DYe7NWWO+kDKUgOg
5WqKcU3l4KfQA9P36iK15pVKVyp89MIw74BqdnEW+gH8gleeucMTYd+0918zsk1jS3KECiedgaed
F9jWulYhjk28zjPaKyMYO40VJ+IYKp5ZouKbBarTJ76rYQ1z6bDboyIKZCnQco4yV3OaadlCTSIf
zFHxo1fZqvNfdLMuJU8SkpWios1lOQPUZfCrgT/ZcOkU0Wemerv0SCFOgOpQSXCmnGjZs81xvRA0
DSyomyV1fh/f/h9joOuX4Z3lzCXU+dAMyq4sEgpnMpNYqZWb3qilzppArYnUYWypBBgGAmOpLjdb
klJ16gjNRf48rix3uCXN+5Go0e+MD64egv95L8YPFgdgz37cfOQXMsfa7bmOWey9p+iC5FAx/hqz
ib0czEChfzKOhiP7vCxurx3+T34Cdf+AW8zrz/6q0TyykNrS+25SvXMevsJQHST9lQ+3beNskG4X
1i9frzp5Lubm9uT50o025vb7tm4JN/a3E0iIicnVJn6eElBIyFvMOEZKLMI7bRkCW2Bna98aCn3c
MrS5qn4nYZBZfehGBUWk8PQgbfHVRL1zbrZXy1HreDqFgNrgeVC/svverWaO54/948/sB/1xq7Y+
DtwGc1dG6qGnrYVurg65+Ip7TS8LvqhGPb/ZS0UUACNwtX+jmDfezHfa/k/3jAZqL83yi50l/2YR
L/IxPVeVII2ryCgsMOLB/RDMqkZUIc7uJNYNV90GRXoqKDecZiNTu+TsJU36JeG/XISwNnNhDAV7
q1CA/G9u88frk3foHRSTxnFQHMSlIfdkKbZCQGxxcj41blCFh0lGDHIiZTiuh7lKgKjguDfo5PBL
aJEzLQMRtwdgyXDe7gijsyCD6wAzsvs13YvVFwRRu5pBzUL35ex35CRQf5BIT7vgrsFH/JnTDfWf
UkCclEJh7SAAJZiub18gjAulK7U1SqfpffCOZgot03Ov2BvpD8GTvZz3SL2BYlsdnIkAgo4s4XXq
cjGFx1orVVMDCBEgmshCEhwwQhwd17ylds3lGAvP9NpaatkDA9Uxc3Sd0IHKXRe38NSlCzD+fa4H
3vK6knx/mhD5iQNyN68NF3++Kl6wH9u/NV2mMVA0X02VTnTyB/ZmYaPd4/29Fy2CWRosH12RbT0I
OCf+GnXlJItcX6mYCCB8Q2MiQB4gMYlO01MRBwKqwXdUGErPAZHmBvp/cri+23BleWveOib3XLNP
v34JN1hrHPjP4U3PnnZjXziWzVaQYCfxW26NSVbmvQCMqFCHxwgHO9ZIenomzzNdEqq3WeJL1tDh
Q/w7PBMkYsG/tkEXULrYB+pG1b9eIYr+2tuqTvN0EFxAitRALNem6bha8WW7INaon2ztjODQ5UqV
JIiQcro86LRk6E+hO6BTLNUpgfspmfuYiV/KA8n8e6kPnLIeSMzpph6ZtVF4YxPkpbLOKBx71n9d
23xjE7K5lJn4L0+zC7geeGnPztyIPfIRus1uwXwPH1cSnT/726SSVTWjqIb3TStmyzVjhknQpzQC
qqsreuMShF4PjlF/Ovz64+wHUi9M1R91TBQtqFjuIfaZ17OMFZFI7UnxBg7GjIIioKtD33Hbk/iF
oJW6scsVEj4ut9T6k1yrcJTPqximzDYA5FlUNxaBh3AxuaddozKGyHcU/dtjQgZA2r8fAoJtX0rP
hEZc7DVCUBjYBwTiG7Zty/K5kb5QEc2Ik9004HUal1KiZQYuDbGSZHQL+IP+T/OuS5HJPk30+ZCt
z28d5nC9ymmV8m+hrEwTp55t03rLF+thX+ZXi00BgqW/jaD1oQix0CpbAmgnETSR9WYYRxznU1Ke
h9eA5Oe9/G+izuDl4UXSdDA/sEpqf+bd7azXOKnRn5QUDveBtXCDV8tbxlVOQOrPN47gj6onX+0a
En32JHqn0g3NolJPmIRtu+gt6pGG1lJ+lt2IzLD1XdofJWbh6mkF/S1PF6cTPmrJ1oX3Tb4Sx7jK
LyBaEwQuRYlVHSzY/7YZTP/8bx+3SG2CnhK0jk+hrE5Q6tK9pXMoKD7ELx4fHQFTxZB+TNTdmfBi
3j/ZJHcq/h7v/Iuq6Y9J8wJOZhtSWj2mwUzigYPXXtqm5jVh82J4eKKcavas5X7ku7pbhI1nCSKN
G95UoZwPle3q24ZvJuhq4fd0eVQEWA00YL9ImZ9SObvGoJCz187rR0jXolf+6qlsCqz2Md0vTUQo
xWPBs/O2kNKijxZRSxI90bfccnanB/bf5uRXXVqejxKb2Njjewh5UeH7PO5O0ltVjVlOPkGGTJpV
j38CimTesOM/9NogGrDQoPcP2nGEz9+3Fpnxo5a68zYiWQ6+4MbDMzFb/PSXmixibz2enAoHthCt
+oNXw9szpwf4C4b3LsdQoXaMnDt+aG4zZBrhGzJAXgD7Iuysx57eoBbDIrWrlicWYhw0PAjCR6Ms
PbDcjyEJJHTPADngs8jliQcyn6Z+FbxcLPtL+HlJbXEVvn+A5xCKskTIiyu5TpjMm1iUOn/AYkvH
rEbLIB7t9Gq6dnjPYAz+aw1mKITS9zm8LViOZEi3dPLakcqdlEKNaErfsAqH9LH5Z5S3gXxbNA1r
6mc6vtkb0b6vL2wDAZv2hI6yhAleYMaheBVDHbeyAUWGxpKp82AaFNxdUEpt/6Jd28Xi4DKCclt2
1fiUHnNE9261CGOBVV1Zk4Cz6ngQZ/9oC049XrsBn9gg9zkWcJa1xoaodfYvRYBa2wqUVMGSGFvl
moroA2/IzE60uIZikADyBfxCFQ2noqpP9hoEVTQ/Zs3CLmcj0cqsnzLCby1ctndhZwhjKW7rus0j
acxhb8Krq6c2nI2ptQwurYSbCN3dH6ss8v+m5tne6Oxya1iZ5FjNVHGedxtbkBXZzeeYfArTr4QH
0JUhhd6dSbtJkrimNjAOfqUpKgQkr3OBYKl1PFnN5mXpsj6BNWy6jTn3N8unXfJ0fpcbeNLp7SgX
23aeYdQFxTFCzmTRjaEjeavxe8QFTlFNk9D3Myvp1y/t9wGXtcRw34L4Tj2dUeJGOfyIJo2I5ck0
UJEqkUhmBYFXzuzdaiqDak33DlB8B6UNH4QC1+n/RFJwWtZ79M30tbvUvKBuIhVHqnNrGlrds+CT
NDSEeniXSVVFvIgmIPOEVXjTGprrHfN5c3wvy6+ROh8u1sQqla/JccmLeSM2E1i3k/XeXCG4k0n2
8rnjzb97UDGHmELZLTrb2bIJzJ4PB3iFCe16FMxpsNomtF+Pk+yzDFpdsI8/7lXP6odKdHQ1yHzU
O92kHFsKULTJ+LOtBP6w3W5EC6OWNXQf1z9sSUiUkqOxmVeD3q9uW2F8lQ89fg7cN7NT21QuQQb8
RH5r6q5xmYFg0ZnXk85cYoKcCogEjI8YHLegCtm2C+RKvWuCFD1InzkZulzfl8dRp07bs2LLBhdg
KiE89sp7I5bSXNkeD4BXj0q9VBy/FaXhwC7me3Y7TDGCDdDhX9JZjX34HYHr0ek1Nj64VNpVIu/J
dzNULepXlfhzoIJTGmvL9uxhYnbOOGVy0xwoBvVtotMe3FYHFLdxkXuPVUAR6qzZnoPt1uybrfaL
71z1UCfKSL86U29Pueu8FM7+QZDxPZho6slHLTcE1i0TUYSWhzXBM7SexPI6D2krNmw+1sZTt1A1
tMmOSAbsYImO3rZyDFNRoX0aFHFJpAOcP1oYzl21gWHR5eAZnS4PQSNKK/yuc38GJGtZDHTbGHy2
LnJGX7aKJ78tTgkXXq/pzaPHX+inyVXNBH5njxyw/fFGPL/G6Lk7BF/zTil0fLypW3p6Pebapj9l
Io4eFEklBUs6Ly2sjZWZpwGMH5XMtNf7IySNp3pO5S6ce9aJmif42wuS25YvQ0uKSf+5O7yb30O3
ru52JgfWniLC4YqK3d+yfy4Aa+9m7jl5UjqjLLedzQnQMljrUMx7K7wcEVuywCn7CKRsZ4GcpApy
UqxFWxY2+yd4hMgBn7eeP2JPHUnD9QiwgqwP31fZOWMxF/64CwgXSN8VGbyKNolOt+iSg+qZ6i4+
xZwHx6itVpn/xsfs8KpMNZ24sp040B9J01SEZyQUOtfDWr930Ts+oNxFJiHL68cH1NNqrhLm1YX8
pJQfT+dlX+xwfksgoCkDm0VaWUg5uWR2iflVaiJno/jsOvPV/+Fq0JGlicEBslQlLpW86T/xp7aB
Y0rL1KaZVx2nhCNNhkSAQUDwCbcp+xrQW4rLF44KVcnF2/a1fn/n6K21dP0hgJFe3qcvZGln9v/9
MlXdCRKxl7lY3cjzF+0/TbybqFho+GU1oHKoe1QDfB0TLKk0qtIAtWsw663+PB3XCwhcuZaLVtsl
p22axPjLSXzdWD8padASVXFxqlLWZ4L3ib/uhzX9hZdX4j0JSaKP58FfqNu0s4/O6IMc6ocFFThf
WpTMWL/tpRsbcjqL4IgC4OeNUz148F4vOJa8/ctv/Bz17N4YzMeOOb6k5C6qOe5843OHFxVAogWg
yhU9rFa3BnQyXT9w3cKQ+p/T4nR085Ab4HBOJNw3R40vTBJ/XsaSogL1z2rEs5y3+Ww0tIHtZ8m4
5cQZlwsBA2SOq9WausIJceTVs+UVKCcKK6d2FkungyUxF/d9e0sFrceg7rIJzykCPyvdcxjW+JC6
5LeKRp2CMNPX8vVCGluRu/0glqqlJ8xv7OTunM9kZUWNEq1zHnjsatHMSE/D7WKQXZZVYLHnzs1u
uArBYU9qnNa65XZbz8XP1PTYarfbJI+JzoSb0OvNVeMq/Ckj2nEnj9/LBrqrhQugLBD+Df04c87k
X1LfoI7F6J8dZjZzZh3dvF5TJcLAptM4liHqf8onpzA3LnQiD9gvwn1ddgw/ALogsNGqKOBfpkez
noT6uTTmEat+ABszvTqmU/MBQ8DTpdxwcP9fMyk7zDU8Y3B9N6OrIDtk+CPajd9swAHzlbPrQDv6
9A34b0cBdnapv/uCmyerGVqHMH5VSSnU1YroYUxGgwwmpvz/ilKRRlz4F2uwPEdfl1Txm/ggN1/C
wLhG1MZBMdlA2QiGNihlMCJaewbhAFe0kbRZik3JH+jTUzBj8raQptVgGU8HTWEKmAEt19PFYI9o
53ZXY8igS8EjEG/sEmi4bNOPcPE3LSWTD/pk13KN71ArEvCK1mGw/Zq5o6sz4toZBZEa9V+7ly2z
CPmMXFx7QK6/qhDWJ1Tw7QhAT+wgI28/FQ9EJ0rrlxSQCw5k5Tpt0WxtVvoPeXWz7DSGbbXvXLzW
Ix09Wzn+BMnZ0zrKcjB+9Fn7euq0KTERJo10tWB6b3BwrtwyfUUY7mDLyw1CoVJP74UV2rud7OoX
uGk0o2m1nVYDDOHN5uGzLid+iM/AM9V1UbCFBxU+25qNWsyGyqWuDsJJCB4PF3SA1O29g9qnA+Ce
LC0j0sWtx/YlWTV2OaDSL1BE5mtHDrTfW4O6otZkQcVzUnujIhFkAbmxFgvPkEs4wysIwKle1jmG
q64Vc3JNCNd+WO6DBWX7/7CTGtb6qf7SdEnQwYX5IpFkHXv18Ezave9yCg6Y3m/cH8OnupRHgOou
dM/PCntupXXcsk4th/M2rXMyuGMn6+fqOML+wLknJ59Jn6MVJYNoRi8apaF7sx7zdZwrRK2eJNnG
IwvNgVGk88pLlPbhfnA4jWyEC00YxiT/iADn5M0s0/Qnox08v+44ywK4L9pnZSwHQ3Q3xvhhvr8C
cSebPcn4x9jrWak7neVN3pj9gMDQl7gqWj7Xsa2YokhfJ+aB0ABZoOO6CoWkQveHNeIoT3QMOvQ9
7t96UaYzgdYN8t1Sv9wmkIlvzxrXb1sfFy5TCGKI14mTDXk7wdX6Ly6RBTiqmJ3C828D9UOm9Y//
NH5OIwYjJMljLJ7sNaQX+pcUWXEnIuFQ+RgZjh/S/L7r2znC8UNRUe1u3H7uM+IevPWzlzPQR+Wg
XVfzDe/MKYO0VVz6IRiV8ltPY8SXlbWYqrWnwiB/B9ziiAwe/Lwjjei2iua1LWGHk6UTtxuJEslT
P7zsVgN7rJaS27osDjyXWLyNv23K3KwEXOqMIPRmCKOdjURgaOfcZ/w7VlG8/kNGhnKwS7cCtZ8Y
6CSKB6xrEo/iYnxWLxj//jNf0ppfgpA2uKkfQkvlwZjBmFb9SdVCbVMPPN1asel9Zs70X7tyxoXR
fgDWenEQmf3xxVaXcYH7Ax/j3vfTBlvo/vWNzpbjhn2Lgbg135OsXWVDvJAWo9N9cupZjAwp1xBR
XM6xJ6bP8omV9lSbDzrE14Z0P20z4yU99rZtjxmQPIXLLgptMxClwafye2ZChGoNnEWbhHBweBEW
wLluAProAoG0ux8x2PXGLXS0UuNbNpLJNqWKTQvT+1Fp8mWvEG0hqXick7REoq8IDkmrvGJQ6GdU
QFBt18S3yVWmFbXB8SEGGZm/H4K+eu4viEgtVDC4paFmUkZK1q1C1Hi+zBC1SK4C27W2btvaFt4Q
iw5RNly/rK1h3Ul/hgWQSmlHqrS/TRvrItriWUXrsnVm/WfmUQYlJd6pogQGy12HJL/8eglCDS7+
jh3ANWszJGNB6PgMa2aaLz9e6Z7nY7qkODXVWT4iKv8Q5no/kHATPIb+N0gFHC0rHDh6FLiWP3kn
Bcn92Kf7mScmqwRyAxYCpQf4CsjZ4O2z8GVNtJGj/Fv4OyHg61t9cgHMHtkx2bDioiiGq1obMDMc
VnNPBW7Ro/i2Ul4QWZR/dTP4BB8zGj3tGRQOxC3phiv7wCkZSAl84AiVJRZrs1Vka1ovSsaXUKcN
u6dgW2xwZCt04/ycJd20fXr1X5c3SY5QLpyC9A+XRoDLSnXruwnXJmcjbSedCL0OST1b3o63GAlp
iM4pxGhRbJ9hvwLIdeKaBqRO+zpmi35/OtxJxzzXx6d/vXKYA6Ggjs4ZglE/Zt4jg99Zwa2MI670
L8njoPMgEexaxK+dwp+lB157ssKuj+Ct59Z8FVHynlVTPYS/SMh0k+jbIp8kopjnBhB9yAyQsj7C
bo9xixTaZ25+E5HQJI62XjVrAZBElatqesXd7PRysNiE1od2PLNXxfOA0pZJg5i7JD3Aa1TB9T6h
K/lHRCGRwIfL0+7qbPUhIMVRhcn7DMlJC0tQXoP2LcYmI5btoTddzLQE+dkCGcu/fb4J5D9ehp9O
CmDswi3CN5tFp/EnD6UX9FCZ/1y+MjY01AS2HHOft0BnXo6nOAfcUWplh7cJxOWFvm2sz2RPmrB2
0kUR1Hm7MrUQ3Pf6n3JqVpsKxS6LDgGAGKBlkCGkNPsl1381X4D7t/ApCsDp6WuwQFsC0Bh+18US
YrV7zwUGe9ytkOmnhuuOGr1H24wrDU89Q8lN3CQQEJPMSDUYOLnIZeUe3cxt8Mx0QUlrFAkTkUY/
T61+doD2P8VaLdZ1LZNwRnXhmwaMdIkHa454n5T6888Q3vKBL28rBcGaYfBSC2ybsFGqUpp+b/uq
C/74dD7qY6/cjEH7rIuZJU7IKRwJtxNpxJJD/XhWG5weQcJbPTzUzc7zaDGR6SR1WB8u5H1rvJV9
4YQpjJz3bJiRPwGm26xyb5x1m0peh9KAvJignu2yGtzrZ2HffCkJV1bBHPPiUkN7GyRIW/s21Bn8
YZPLmr76U1DPRiceNHxAVs8pobelsnU/gOsmdE4gFKKa2CLZFEgwQkujVNJXZP4q/sVbTi2AwV8B
HZ0Lv0VugP2KIJhmmFQ3Sd3QXJb/F5qZwAdl+MFHc7xqK7dbcz6i4Wh5109YsDhFkPUZfUSNR8q2
FbdXW/n2vtxV5m2QVw7pSUwDOQhBSOUuKIjmp/D0+hyjk9/fkkOPfp3FYhcPI9kGdXDeUYNc8je4
0eiDgxLxT/hKHgWdAWNdDZ+Ri7xU2tO2kutG1jPw7jpaLabc+Lvyi6bwh208EWUD4MosfRPdoxi/
14twOYsPMdVCdtrMTOyfzc5SRPADSvC0/HIH/FIEHPw6hqQWnOaeuCZEb4I4R3+veuvJoz/U3HHR
wxZtkw95zpIXySvnt4t/PKfCWI6xj7lQjLbxo500ne4R67mfoj5gcYwkYo4X80Sf9FFCRxZ00q2k
9sa1ExQXPtGqrrgNlxb63bndQzMRN0RWQHqsoe9Y3QsVQVR9wiExskfNQ2NAZnIZgSMV0ytFfmF7
9aRwD5J71lRpwO1HUhd0yIv3P2rYThtfIreT1+usYRPO0DwrW2CMcT26RMCiDT98NK/WXnZBuybD
RZiG1P7Hymg3+cgHoIw+6aEcVcCae4vxgxB/lQZbMzONQnlkBYzANIJmunJEbSkq9F1p+3rBrKPQ
3Ev1eVmeubRBlh2fiTWa5mtAPXPi/KwdBUP9ZpwlT2+u7iLhtmOI9HdzJrwY8ArZ6IGRHTYIQpyk
jhireDzMTvuTqS1zTHIHpSf6iN0XxuIRkxjrv+0RIzWHBJjdtZ2phT25wYBHnqQ69kYMaAjt2gXH
mpjbk0HIGLe5VVHtdKCy6xujSjBNEw7cVD6wrJaAVcpRxkcO7VmNnwmjjvAT2DI1f9JqszYK1H/R
jGlsOiwsYFDwQPK01+0BzrAaxWZlMJEpCrMYd++S4OsRJ6cp4U3cX4Pg6i79bxdRChh/Hzpn1LRz
Pz3OrQApBijAQaQtuHOY4OMqhlPbGeaDjP1b8j4dSaBNpsSxprdWEOoUMR3SRk1CZonPQf0Ipch9
GnnEvcEKuTvIACjptJB5T7J7SSECZm8d8xRLuhuueNjb78dgNHnRj51fs/ENNAZszvOPQioqBDau
wrx3sURCuzZpukPsO+auAskHVDRUAnpUKblAzyIQMk4Seblp5L+zCPD45q/qG5oOt7zbWK1t3AnM
IaAiIgWbEC1zdywTlCGb22KYHKVo0TgRfyIPxOAzuONGNV21gkJQiHyXl51j7IuBlggB0wKW7/+d
6gCUbZMVRtUBkygvd8PqFHg1zGJjE42Mhn/LGXaif4A+9pAq5TPGoO/iTXvoSQQLt+EQ5vRLaWik
bg9de38TZxgWkgBzfFnory8x3oebNbmJAs+GPgEH2btuRWjxJAQJZSZVrBXzqTfs8l9oU1jk4dMF
kZrJP780/5xt3Dxdooe1t3ICjT4P6ltkQ2ijr1mg5hFdYzPbZIwKtkuRzvU498aEy2cS+1VLSY6I
8OPPSB6pAdPOucFqhrlto2jg2D0leshQ0wSWezrPwEs8+avP4+OVz071naJVILXgeWuVGU9DExFQ
vcnOKH/FcK35w6GD1oPdCHyGSOukkIckvtTMwK8ZX7M9ahvCXSsltjDV9/E8qSYZmPA6scxSCwAY
/g5zVYvdY+i5yhAQUbSw/ktG0olsDCrKQCVuhim0iN6j7mZaWtT4OFP3dn3UFpsn/MdEFPhieIb0
qgOeWugdY8DZL0B5K60rDsfu+CJPyF/8huNEyzpRYOQqGDlI2xZeEd1YX8q3vkmUseHLwpyXymY3
s0tZgwNwtV63fNykQGirg5eGQnVhW6dd9hDfelZfLDksakibq9mU84/z5/0b/HHEj9Jv7UWcYKLc
WyFSPJp9QQKI7lmzaroqJlJTboXVLijI06qriFnEiQNhr3lgE/VazkiNSi1y5kB/vr0Qv7Nt1qOR
exFK/e8xT8XhnbfRC79IB7zKhvnEMHW3ZQKAjB+YFszmIj6wFB8p3Gqk3fkqQj/KoJQNKtQNCxhO
i84v5Z4M0wkanvI0XtvT6fIo/WJeHymSZfvcAzts1XGL35WA+pNAklC7jTCFFYKIwt9rhRqDxk3x
rx3SukKIlcHzZePghOKRPnNi3OOU8PTambtGDX996SQK/cQoFGlnOwd6lowMMQ1gJWt9RXGIc67A
PRpuSbk7UWHbe0VWc7s7hwt6Iq6KFBHoXBUpNTNQKXfPJm2AWMgV0+so4VwSRzn75qG0w5KrQRkO
ZTmZzjYrOEjGgOm47yUs7KP07rwaBe/MHJyfz0LdEDNppIU87AEBhcUP/OgrTfp4Om/sMHfhJ0AV
8VaIhWk2PYauQ7tCEtmiJWz4Q7wxwxpjMC4JYEq4voNfu1KrDHt1p3cP9O3aUQBYV5a9ThS95qD2
XVi5SoQI4HtNpXW76dYupe+MygflwogqFR3Ion9szmuIsooLx5EYlB2YDKoVQZWFt3QmC0GhNUeI
lPlKXZ38XNAif34jN7j2a6GBxZeLiT2Dt1nDvOdo3Ro5GqTm7X/jLLSeTO/o6Kd+BASNV/42tiq1
2jZJNW1i5eelHhPR568enB97D+yS4+JAW7cZramd95cWjeLTlrFfKbvsfrzcz7SWEQuMhcFWEPIX
6loXqcj5MabZSlCVulpjQGJDjU4QVuKPkYLdE7UlMuA94c3QeAlA1cSUURGTE4eKXRI1WnZKspL/
kksQNo5nL+DKJgfzQ2JvC5//YGWs+59L/bMsm8MxPIkz7Wid8MhXnc198q75HTVwFEPYeofWdaoS
4DW8KsaMKoXNijxAMmHUPxY4fbefah97DNaxyu/bnsHYoHQ1UtL19LeqDTcT55vO+sAxwr3a/Oy2
dtTtYfjav9hMp/mhHir5tWY2pd3WOiMG73XcYSClRV/LaZGvB/6xhK3bcEw85XdKfV7il3yPv3Q3
rJ57vV8ObhLPFPpmGTNetfFRCQfsFhDGXvTOeWb5wJMs5eMYfsH9V+JPCgD/a3MUYyL5CRIjUR61
e1YRGYizxnwjjiUSHhLNNY9U7YzRELYTL56rZhTjt+rrfg9a5Bq1ar3mY65jYqN3ZcflikMXJJA2
ggc2bBCh/a8sWgNrG9Rm5SsJol43jyXYAQFhqv+8zm9bhYuiJ36L2aNiPv/rf0oXYiEl7W603egr
4dsayR4fboItJiiGFIYRy7pacgEmV7GEejouF5nr53rGElLug3kyu+ruUijtBp+yal6TLeMQVs26
1Gj6GEpo36Csnijx8DqvNeB+slTvguz6AgmGsuICtUQPi7ov6l7sknwaq37K7fFA1GY57BJg/EB0
Ed+4Kj8ycPaCPCtyo2LoM6MNg1oE2ygy/XfKib4zarb7yeCr+Ml5w8Ibj6KZ1DbICF8/MPoLXMiU
xmKpgZumj1F3JgBhuxBwkngM0bCXzpoKurs3m5DWvOz8duWD8yojekcY3cIh4c1FCcBc1t+Mvlhh
/ViYjtgyHaDE9+jGM8UX7hohPl2JiheyR2jKqEt9Qd60JqG33DCeJtDhpCMyCqW0TH3IhX6Jl26C
REPfPpl6CLkeVdPjgxGiarlwT3Ev1IIOnjPEedSGRV1C+oM3q3/qcPSw+L3SN5q8KT7Yjy+r5yni
n35oQtEue2WJhp/c81ELMsDIhULmrHaHDTL+OGbsBRT9PaPCQEMkynJx2cSxVa7PicR4C17PLvqm
T8oEMk5A+VgYN4lzM6dYF/qrwFHNksMJWF9W+18vj6RT0SjoywbtVCoGoGIf9Vvuopy+20ji6koN
9A9JgLkptjLcG7jklWzMFFS5SP5bQhFeenirCsQTUA7oPjHd83TLSS+spMVe4tTnHVHrI/iHOwg9
JTNu+CVM3wvTGO23ik+ovkCDkteCEQZw/o4pwPIGuc/FwgQ0rMhkIs3Mp29kdUwF31wfSR9Ll8Yj
S/Xq43g8s5fcPK8EeZ1xU6vbKElvryIQcHlukyXkGU3vTl1+LrazgmipHTPXyY05AvrUWm40YUWe
ntxWJRcUlC8kOosukvJu2y7NXvMySWf4oi8JnKNjsp52kwvqFgnCDhz2+Hu/PO1hzi0mbUW8S2pr
x5HneCphjYl4/aHo3d22aY/lmqcacDp60YtsyZK8r+WfL5Aj5I7B+lq0P/dlbVGCVZuN0n8tRjx/
UBq6KBgNADIa7ERk/vpAVqzunN/h1CIdCzbox/XGY+pzvoHqmu7Os9RgvXrm/03sw+zbiTZZeRf/
HczKwXwSVXr/IA0wz2ikYGBwRkr+ZFH3wcZYpzQIAW3fmMd8ZHr7WLE3HVo0cSRTNjuOOjyZ8V6h
HAKa4dWdZsQ9vujXYY7MmkwRfHfMVOUzuG/f3U3qZMQt5QnZR0j2GTf29g3ZcARsH9LOqmfiyBg/
99Z0I26sBUaCawFEU301C35nm7HDqVPm3EHavh2nnd4DkZRlGrDXA8Zq4P4tfLv0Qtxc9tSkG2zV
3XkoWTvg+OVkoECGorICvOjDN2I8tX9N2tRyQBzb0yuFQx0MHW5Qm+eu6miA7DQY8kjEpn+iVLDD
5X/xh06h6I7yJIHxZj9xiP7Vcxb5Drq9mGVHwkng+xxHJXEiTaf0U5TYwPCXaPWCIhyp6Q8tBkys
kaWEDse8eW/7CGU4bAVNE12vVqLmJREPCB1OndqIs9TrHYP5K2wA5LKyh1WD2G1q4rV0EFt3kpw6
ho1V9Sag58ciySdhRu8+MGccAeMWOG0J47d0ZRD9moqWxyBrjKJ0ltthQ838ATAnzAVUEp2z0CgT
1IrmJA0fNYjkpBFL0OMKnIJQzZ2YLwYotZ5WDODV6T7YCUlh2g3FMBYpK70LYiRQDLpRDqc6J7w4
t+z8VcGm3FonVz0k0TfjOGFZYcWlvWjTiBIo8+07A2lhYkLeJ4jAuOnwhDAg5MxNLKQzpCqba7rJ
IhkpghY+ylduqY88pMsiZ0HxCZis9Y5TFz7/WNaFcS1IAae1sebaYWa9bC0h8pn0nlFooP9+Nq0b
HhdVH7C2Gi408oqBVa5i82vkTHmoEeftavCFOrjWi2iHojl9zeN/8OOHskc/p+5/6jAi657x5Qix
0OKeqWGw8MoCWpe4rFRIOv9e2d7c7wQ2c9z9MAZcby0Ygd0kr6c8KJJ5wPgFp1GinFQgYPhDmhzm
RYzL1V5uoUt4aZYuFcrXLzVom7gLbvUC9Be/GnMwPR9UJ+IXr1G540rFnbjLrshdmC1vAJmzhF38
BAoI05TMwDCK3TSRCH2uPK1m2W8OL/Vu1W/hCN1dnZVVLrBCLu49GPsex9T08VvsdPLuBcg+6ehQ
pScXqcBsCSa49Iy1LPYwQczw+JOGv7tH5tUs2pGvJtim8h39ZLN87pw8gN/wvaEL7Ztbbu1fqXHQ
awomhT761gAbZqPAu0s0BFTUtoqnIt4u4KRO/9tqb2R4K/lLKK8coeS/6UQeI8fkYk4nC/WF3LiU
/iKYaHdzpWDUPm2xmc6v+lg0vP2zPjebdjBiPIIOOLiJ5kNMHi6B7OPOJ/pfhg6nIdkRsdEtthrd
xwermNnntkCF+LsDgn8vE3hqqIEs1yZPAWFyVdsLjBTW/gYA++8SJxg/OpM1X4cPTy8EkacyYP9y
cW+GLphCmcJMvbluka/5wZYqO8Irjus6t/5JLyThNwdC6XatunIDL1cq56ss6bj6vUs4OThMMYim
KgWipd3qXzqqRsRRHggPhiPWc6V0uDO2Y2dY2+H8/3t2g5hM7XdZIOuD0WHH0AB43rKxE870L4Pk
9HOW+9ptF+eTjWUR9KzA12E8R4Zi9SfB72OXRGatdnaiDlHnLsbHrSjbXmE3BL4YLpuU5Hkbr0Lz
iwV1IiUan6QwRiYe5LIlTmA3wiepHn+IICUhEKKGH79MMfWUPrxYdUuV7lXCKQU/YhRPofHbxIZd
NMy8iHSnZu/m/kmxeb0F7Wh8zrikm3QtNxIYUexEx3TOz+hUAfhlEm1JZpScv/pK77T7ojC0z3dw
THJDZ4vpJU95SA+VlLQqeXWDcLRggak9osypqPlr0KpfX8uWDgCHewltnzRqRR8z11t1o+iZKd8U
GGDx1OmFs/KCYW7FjTM0DSIClNTLB9qTzw4FrHhLLdRifCIvYPjTiptUOsEnS85/kLCd0pXE1jjj
OIXWsH6AsnLJD6YTwhmV/lA7FSkRW35MKnGInOzdi0I2hpUHR7FVLFu40lJxbYcs1lsa14+IRNZy
8mJj0bjK2GNLgM5SeBfrOC0/Q1JhQL6h/JWfy1XoZRDLLh773dI6puhanXxTtprQHmDWseMbxVa3
AcJqojhTrb2Q+CQsPAhgoTwL6j7F8MnxaNfmYsEXlCKUiUF/Zdvbw8yNaUJSm6hhb2hHZ645qvnd
UCDgAlFoWAbssXRC0zDpzSKiwjJ4TKbL4uHIBIi1FGFfQYuRVWW78SDWhRKhZqCyXfdFkrefStkV
E6Su2jfUfC9jd+YJlz4BG1AUNSnC1OY8zZZ7CFPM6RLv0imFoL6IrzyZy2pjp60M+O/wR4scmKgy
vv7WMnRQLROnHmyhZtY1v1KHk4CfqreeeOs5/eoe7eJpZxf5WUKxhlLWWGFY99F8nFy9sxZ8cc+d
EsGPbJLXqapuCB+DDbShrO1vCbgDK8xvjUbc6f9rMDc2avaBngff+xSYXn9ndAnF8u5S5Ook55Wt
aGNaDehqE0s9oZfwjscoej1a8xH9GQPVwXhqzMXlL5cUUF5PXA6RhYrpshiBkfjgso6T/de2Ilhh
uwuwguXwTrvdjkog8ku8gua+K+z8GERehqPpUXzGScqQ0rjCs/96EcyB31v84226ORTc17QQwSBE
yJDx4N9e+pCyT7Fj/oEcn+lIXNhTcwnCZ6zqdGFsIx0fJzh7SVeFBVnJ0hr0kmn6EeFvTjxLdE9f
nQ5Wz2WNhLyuPAszXzkBj7koN9HHnebFgjhN5xyA/mJxHD/F4DYSvFf3d7zBWA2wcoCb7+tlNv0e
vvP6Vq3bC6ji2G1SAGANZYN8RwwgUajP+TOCobJJi83w0toimdaq+9mVwXUVM7t5BX6iLIxo6gSv
RVIlMIHU48bBki9EUtiEFquErPBDUZJHFm96jbBzgr4mA9aJVuTXANrqsDo7l0vfetUyXvx/ckHG
Ej66KYbiSW03d+HVhr50Mem8rqfLJefw+KHtqhkRwXPA+nztT0nFx1yL7V/pKGDcSKIRc8ujyJX9
MK+DL0Xn/BWGZNYlQJH53z1atDaBks1lFt6RrxjrJgGZxbUO3ds9rABW14lRN2XH5EC+WbxJGUEf
T4WgxT159h5zS7V5fWPwaE8XMERvuJTsAamyskl/EFrx9KUoaTfoHYWQMsNHSe/rMeTiHWHXYh0l
i0KtOmbGCYT8O/j1/c+EkiNJ84X+yy4z0aCe52bACxxVqqIqQGdfHJ2pt+eEcq3Co523QSouoFJk
5N5TLRIO0BKSL1VY50XblyFrpCnHaOGdJyrqqefQLRbHnu2W/XloF5izrtwDSZnD0cCHtKWt2LmW
IqZqyccIdpeHvD+QXOoQ7TeMY9VAVzZ4GJ6qsPG+9cxP/sROF2BTauUAYdl8ML1sT2YVu0/UF4zS
vQVcM04oGF72ntr3twthq8mS3v/48Eugq7RbEAK6amoWPb/CAB+5OXyzHK1hsR/UCWg1X23Xp85D
S+NFndx0mewULgvIXsR5b0DrYkgFHUzgl0o4YSsDAl7LVLIBQmon1TS1Uur25Y9bI+SdUWwcS3or
nm6o/SPCuF1TJ2HpStfaLzqTZyT1O2eHPtw3AmCvZyG9aKhC+KJMSuqyA+Ovcy0P+RmR8xXdChPs
eeqOQ9QgDXnlcrutZE03y+aGOtK7CLA8ARhSWTLWcaJ3O/orhMNZ806SpCvYZZcO+/W86dAAWbfk
HHMqy3sBnNyDT0rqckKfq0LVF7KyLXF2gW37/GfT+byVtk61yna830jjICHBzlBgPrxOy2NbPva1
iTrXBCKnHIpfT3rPpeOyB3RlwIb/Lyz/EwVThLdl2nnr0PkKW9deUaIQ+1tHef+pOlCCWvBg91bZ
xPLzk3VIzeSrUosYdfDGxCsCuqoXqubVhCK/UxWvtITq23G9TlEdfSjWp1OWAZsuN+Y/pScrBd45
iXvSILd37E1XbuwOMQmP4HijrWPCOiLtwWtiTx7hvTzwQ0Fh0rBjpkzYtogeSlo9TPkgVGTU5fy1
aKVBhevb+ihpg6iNlAoGP3pomAyAdHtyLBwMkTnozrSzDYsVob6qR7Ijehrqg+yFhT0wWXplxfMB
smUpDjQLAsE+Dc/68o1Xg0woJBeKTUycXAveC84dJHxTdfvZtWGzT/8g9yBOm2C3D30xGztc4t0y
19FBfWE3gVnScOXz1xlAhPMfQJDH9ew4s3qEuKrz1RJ2/eTLXP5uwAD/QcyQquEp4ILsERZrNdsr
5bL2tkPLSaYbqvyJGFuo8mhlGOrR3XzZ8miXqIIHKyYoJ5YpeDhV4DwahEGhgvvgx4/arYwNeMiP
1kJmF14RKYpn5Fxiw4Mbv6RON8duhygekmIs1E1vm8fWHmDVJY0ea1Jm0LRon2dfljK8XTXVpBYG
90EG5rdXuSY7/iomYMg4YZ9jdxg71uMZl0M6Jk2Vrcd4GGfCbS7WmoW5BBuUj6XOuiqsEzDfuMv/
WLQpGJ3FOUKetT2mdiLYzkciPSvdcskjbrsHWkCsbE0ueCQ3yqgMbz6BkmHCcXxD9drMvry5iNbA
Yx+gK2MmG9SWSF2LduwnVRhwcoZAI5MXgPjP5z8aEM9auScvn2S5CIxmiR5xyRjjIKzDYfOHx7Pc
dxsrc8cgoo0kvNbTcygebaBkV1ah/Umabzbt40CmQSAF4Muvoc5IbjSpeTqYKi3BCaJ0nPuj4h+q
YTElMBlZ9t3UwoPsRVfGAYNEuSmdDnrZRqIuzHBGmLyAmkrTfQmXUXTuBN5YEQzwzlEBjb0fvylO
GT1/idSl8lxyDlnziEIQaEevNEVEBglCQMWn905eB5HbHc00TXNqupbnalqmDkWX5Shi7BnAL0GY
Ukq1+Vr+qDRkpv5dY+bfUCsdeAU1nx9o1PC3BaUIj+MU+ZSo0i7Efy3c1hjni6mpCC8HA3i0HXOq
pLSAVh8KvWpR0kE2Gqrx2iOXrVBYyasluAD2x9nSsPXJQ1u5Sz7is/3C943JVQdAFjBkKuQpbhbF
d6s8RdYYK7crQOisOiiqBXMHNGool9U3EkgXdDuNyqHo7PugdWsQxCtOLvr4amQxWqyoi6LWe5+X
uVJjK5PxIxvQnHfi2SbTBcELHo6nHu92QQpLVlRRJwCBebyhFsdIu9wox6Nt0VR84bka7lWM4/sJ
xwP1dmzjuegHFUTtATk45nuPM+omOnyg1L7hr8FTnLwdfM5DETTntaAw1wr3Iagc4uwwVJnhUEI2
EMkuBWINXfVjX0HGAbdhaZ3B1YpgxKeHsMkjCmAMr8+dvHy3Mk8Gsy9LCedNVl1Q6i+/1wJ/icFW
ca1bhKpCZz47kBfWFl3WUrOoBI9BI4BKt1QvQyo/OnlKsn31nxQEOAVUeaMXuE2/ZVDjKg37PwR8
5mwrVqYIh1JuCKzKBVOqRFODFrbgFcWZfdE00Z2qKI0DJkBXjS94DebdjSBAEbgsahrY6xCqXqXF
8LPZ1t3MVZDYSMt1qwil1LHRDn/FE/j7TtBMIwipzmw8B/jPDyIt1OT3mKwwWtUfqudwNc3FVmNX
ZOiKHRdwO/OM2kFoZlPn3Jj8XZ74T5lnobvfr3OZua0uG9nFsECk9wNTXzPeMwnuIE/7HQeocLGS
XW1w5pE1avdgIgrIEWlJYtfGpwOkXPdh10zAaZXCr5qEyjHdCgIxzAiAcu+OL8xDKUxcda/Y1/F4
iDRBHMKKowd1fOkoLb+Q3a1KGxjO0Nqm3GsU4vrMKJbSc35iSmuXRCxtXbq3aONM7Ju7e5g5R8i6
ZiafzMBD8WgA9sKuxr5FEvU30IFZg0wB9KvTpmPpEsv99UWOP+fgMjSuDqGzyiuU5RKLhtffMQ6W
Ct99GYiQQ1s3pAV7mlnGgYQgpzSx+QisTh19IX1GUaDGXg1A1c3EP8GBX7FPNSO5CCuOSf6a6dOj
JpG7tBGf7Dtr9wQ9HmBJQ8P2GZm0Z1kRBTe6Ax173cXFr/ccO1CEZHHvLub9y81eoesE7OM7IQyc
wjzEl6ssyz3zABvC3/qe8VjhAUBg3YNMy2Mve0RJ/XrEq+SUronpiWg4v30Z5tyTmjIQHHSF3Tij
wNidoIH+8BoBbFh/6Jsl5l4IvsXKHchMbA8ibQ5OJdLZxAWYnkJxZ0e9s5xaTrgCQgJziVeZ3KID
bIOO1stmLOOvj6qt8/5jD5k/iPkiaqPNZSXVwdbvtw01cWGNHftyhGybpo76dp/iGQEqLanjxyKF
wQ85+AEBleEYEEDuwez0ij6F4930ztWoGx+48JgWcj92GEs9Shpu1lIHSN0WugjSx7897zBx1UaY
jnzoGu9s2q64B5jW2658AcaPxwXk+wUPb6P9Tu3vO32GVVWbAQfCjGsX7PbpqaFg+niY7ENH+EK9
UEwA97wlmfUDpJjwqTC/+/eV4t9Mg4CtT0Is2KFJkQf6T3hLNh5jxw2y/IvaBtlBsptT+qYqzG0y
CSLvGNKyrccuNtCnpt8O/IC9G3jRGrR20RjDg2gadxNBN1ypF97+rkdb3VKpJGbNd9oGUqhRwJrx
q+wR8k7ruHC13dyuiIrnzL9dITFi2z4AWNimaz0sWOhQYT3O4lsKBznoUTUo2wLqNhoTnAnMxchj
o4iXK9ZY8MEx23Dvf53O2gwj8nnTfGnWyP4bmE25ERtJf3fsSPcxyjjA+r7GRe13uBoXQYlFcmVt
KTFL6xw4SbT1Kh9Z2kkg1TqhnBxK7ZBLyBV2RCDs/STWWK/anpwULwWvDw2M0irJJhl5eCxzRHqP
lG8iMWAt4mOA+zeHaGMzpFgynBuQKjuU0qYn315pb/B/+o316wf/i+hEqbMMmLUa09O8JmURpgWP
jLg3+U/3eFEpD1fOIL/p+frPo08ubYmzGQtQDfKZQwEztYjgmd92ZJX0q+sZ/UCJ6KWP4FjtiblH
IGawjHCodTjiMByULTLr2l1W08zjonQKegaQ3SoyNyY/Jh+ddt6MirZC5924jvnuVr9PFrk1RqiY
DiJ6PkulZjaQm6+ecBUyfOq5SYlfqQm9wPz/9LWOV7WHfBWl1kF+r0taIZAB96QotSNmDlw448EP
Qjy+72TmdSOXk57gQvrNmdQUIUhWxOs0123uCWCu9wFFxbw1e9qy2M27WMrJ0fZRJZ2REOANwLD4
SJVEt2nIkSen36beywzPTYsMSvTj1acRyUGBaEGXw28A5BK1cUfwDu8o/1lR8U5bCTdXfeZ2mrCx
h3P5g3jAutG0D82x+mBzcXmHhR4WDHIWV0RINDNLdlVUs29EXvJzdNDIr2PamE7mcJr3V7T6YKKG
GyV5VLaGkbbsZpreUSj93eb0a5bK8HxA7NadSHWj5mQXzkeYUiYp4ofyO8Q7vxD9gXH3xTitg+rR
qvjh3k7h3PAg/aOmh/qXCBePftV+1uaZkXt8MHMwKxBP6i7i2TnZpJTRCA3yr/GUshbNZ/G/fcDn
CFJ23lG4S/7d9pGUjEGkpZud6Cjh0VIXogIWh5TfZxrMcxKQl2lni4VHIyz0nd5MQkq7dCrBXjHy
3rt1oxG0Xn9QCunI6+KytYHHnVkWvFZGAaXJOagX6fLAYiwMJmrCX5DHMv1Gidtud/DMhdR2CIci
EUgxcD7wshzC5GQHjCiSiP0lNzPa/zvfUo/yHQO+cNzTcvahP0fhLl9sKjkaVxf+vKoXsCChzMwG
6Kl0necI9gX1/d+7H2GMYxn+9YYiqSrJXFN3HORVSx6RzkwvnDj17uBka1OvJ9NO32+1OOuevjyy
REBVbudpglwTOugHE/eC8pSjbJyZpo4OX5NTL8XpCvCUVDXxs6DufFIDMhoWcs+JyUEi9t55f/B3
oG60j7GuYimHIUFWmRe/C6KT7Zp+qaCKU2n1X9MHQ7LUrfgEJn/yqxgV8c+Qu8GHR5Us3Ttynhpg
2+EfWDPJ+TFeWzsiHWpGJyFnAWSW/1oJiYZz3EunF9jSai081iwc+rmBbx82YRhgTs390VwnV7R9
jULbPTKAD43VKyv61dNKkoeamoc3x1h3r3mVYCA9j6eqsVUMxQzljuPSQ6OBGf1C0pLtTTGAXa/5
RxUNDlClBTH+FhLRSZ+w20hE864HUnLd1Asc5pDRLgzwOedgz1a4VYPpmOXPnEadSF+f0SPLadfo
pPVv3vY+QeArAhgGEZQDksRIIal7iid9CMPQgoAGEMroyAJk/LmcPlZqNFj5iTgM6vJb/jEYoCbs
D5CKZu570lWb+XylxCRKzkAYj1dj/EocX5OtHJTNXZVvdmNpyibTbHZZaN9/t3Ny758VfZcvs0jU
vyAWqL3pOsWBQqGXnrmiIyU94n7VOhSw7WCEwHQUcfRcn0JdZfcTEKI3ve2srhraAqmGOlpRtOrk
W0da7dcwPGDykJbWKdayk45JHKvy7zfTi7g4Exgx2H2mnyQyPEhaOoGh9RIJhTmVgbCc2r6YVmLU
BqcAz6X77Vogx0+u2YYq4FNWw5V6rl3p/jR0O8kdXE7T7HAatggRHqJDS/18r3GE3ELOXypNAFNi
wKzsRlnyIJFunRsuYXCcw0jk0Yzsane7PBsVL9RtbCMmBgugvHOsmK3XBG2j7xwEZf95u2Ydgn7M
QNtdkwMIXx6bJjdWznaPMf+qE1GSZVo/32TEQ9gmltAoscZoZqsDmLhN7ey/boOMQbwVCPAcGS4J
Jx59eCdH5/GZxsieO8xrj0plbpD3Hp+afjQeNbqTVKhjl8R+au3tzNylsUHe4FY4rGVWLGFHm9JI
XrxMJk8IckRXUIyGKJU2b4Q3dJhj3AbmkMfUt3sYjChtI5OEJpm8NakHgebQHtWqL7ZhmX5oyW7J
7V7N7lRQbdG7r9AMqhiNIHdfsAGVE9dGv4P+ZIg9t4PSTS6VYBUgJZOx7AGixSqc2oY7ddMu541C
sMv8EKLcAjQDD1okkudWbtpkVlMu6rHQ2IwVKLRjXe+nFbilc6IZ/m63c/KnMWWpO+/D6kHEkE28
jSM4l9HcIZ7dQVfr6CMSRcuKTtiU/MpGvPYqpcpCKvBEGTjCHS3DepsbBLlH9N4TBRGLrImkvHxY
AOJEq1RKzs4/CyMvuLh3HzArqrdlbokb2NqltCfYKVTgpm8VG3BIcEn9KPA/yaC7vx32u3Xqmm0y
OR7auyi7NXbPHtjuH01GN6phkYjjaNwsDuOPTEoRMIg3Dp5Eb0jkPm1eo+MQmHsJmnmjoOEeKjLS
EipMlRGr3et/maSzj5yhz+w0zCX8ow4GnuiPlPiUVryDGuYzpoEgSO/5RL69DvaWqvJQicdYp20i
rETU+NqvEdYGgbL2edSC2KFeHdh63A4OKaVTJ1WzwtfX3BlomKjublXm9+ng1GxtkQpx/rbqn2xw
y+AhqM6YDHH/lLtSLE0OH8hokpazY12nQdaz87p38hRHXx1VlqOYpB6Ip9nkSH6ooBGwOOfAegML
TNxya1akekGo7Nb/+z8X4QntHmCnKIyPadThAag2g0+aISAx8FDh44bkuYZTMen2YsPKFTk882BC
qHzJ+GjspHSwZn7Lx0z35HSvWUHbde3r5KwptY2lS119Z2ZT7PcWQOqEDZMhguDEA3Z1mvj91USQ
rL2r8KSth+XLks8qZyBcEyBl2+I1hHD388cCIw0D5tCvGveyimMmAWx0fYv8jk8GKnXrp8yBSvmp
7p3MR8KSVJK7aCje2xFltbEN94QdgnJpHnpCi76dkxIiERCz+dbfXcxHAJEcQTjaa3e3d8eAd3J9
6IFxu/YKs237BxCMFBPcNSv41Pi4hneDwEtwVL8GSMJjmsvlZOxtIXiDISWWy1KVgxC9Eaxblgu4
GdY+pUCaGW1iSbdPOF5yJadOP4gDRt3dnuP0Yd/NW/ZrKhwmRk6YHuBjvvSdbBQbR13nPq8AUC6O
zoMYfH9Q4a6R/kVQAR2HDtNzb/Uhlso7vFKDND0Y5loBLdtAgSmIfMAgo4RPimeqb9LmNXsibG47
m7/G9T9ziSqNx2mM/BUNGk5zNq3n0lXv9MIZs3jmSBCCizkt5FmVTxUmXd4MHzlmplddQk15yi3P
KGtosIzEEOtK818F8V97sCP4bYnJLHTIAhCXEAwuaMVPNXEm5KJvnwmRoBCl7c7FctBUlDiiP8FO
R1Sd+7pHM7dL1FPdW4HLr1qj6s17emLX9jQucsWG9rmp7yhFRrB+kJ7n7oSuksNxK6c1V639rudd
Z/eNVxqFwuNUtCr436pndnqoNFB2w+nDnrzK3t5vW8UbIVHpx9AUMbaV0KoulelH7tpnYoY4KzyK
BMydBvmVzqN3Dz9TPhXxMb/b5jpPA6uAWU4FrTHHpmXy62mLtrq/UAuaVie6bqIbaM1ieFCkHNqQ
FL5e7JlMTvvfR3EhPfOyL+7j9qH7PXeIPxErkqbAPBZeBKvPuAulA5JmC09tcs1tdGHoVS+w7MgA
RqdrYKO5YiBd4o1AmKroG2ImseMQiBkU7B3iwYeabfRS4CSwaN8HOcWSFXYXup++irlOdm0IHTAE
DE+quohxY0pn2ng4ZYENSQShzcWMWNI47JL9PKIOo+oYLv+/Tj1FSaGlBRTXVuig0xrI0owNbVS2
w8gxlMaeVw/hQQHCkgz3+mIRoZQZI7ygg/Qp3KZT9EnDyruals14sWh2JaxuBySZ9ZZyMTkWvqIB
MLZuaV5VDr6slc5HBrpyjkj/1fVkBlGZ9maeKfF/sJL4EtnvvqoiG+gk3BzXWBPJvtx5raTLGKb8
8LhsbVfisfwotyCZ8a0Hw2Bj3V08zEW+HpmTfvXUOstM5+fzy/qL7iXv5BA2LdMn3LXI9kIC5Jhn
VBgHWw9LDGp/KdOmYXZzwA+j4xh1zlKUT5I6jznmlikD2PKzIcA7ouRNfdyv74r0y5TTUl3cTliV
Vf8qXFH5zqZebntWg0JLnl5se7OfzBazOpk8YuTYSoVGHVozZT7uMx0NwNl9Ato1buJyhBVZOYAb
2FEz/ejldww9gaSMEptK6qPfBeRVO6ZTbUBoTMmweOwt/Cikf8DVBPRnwBBP/zIEVZpY1Qv2JNp5
pmHxjPBbRc2QL71ooWgv/aKvDs1c6/JpB2hokixYRl5jcaagq5gN4S7KOuFds8Jj4vtpNzqsbs2P
ypLrKf8BqadPTFQVr+whcP8aYz4/S1gBTRqOOpOte9pKBUqLUbXb7M9A8SSKDp82G96sdg0tya1I
oBKd1GPRmSOKpkkxTCnGBs61Po6t1RPmfASaekHy2LGsijEpyteIQQGiP5aW99btFmLO/h08JovV
IPiDIHfG8t8+yoMC9hRTZn0efHdC4lg+1Cg4IcOopIaf9gpqdy+Kw6wSKIX65N9Kln5H2y6tToat
uiIc6O8Oe4KK9iTBKSTYJHTmgJKi10jgbFyAY9H560SX93a63kf31mewKXadO9EliI7O2ynh6aKZ
15yuaUYhEPNLDC5mpmq8kW43JLLYZhmxHPm8ksoKwSu39czZ0jin5tQlHHrNds13L4PlwuAgYoE6
6OjRbJFEMF4aMcsztgdN682frgLFK9CAcIgxFz+YbH9XS3yiHwG83tRAbYu2FsMSYrAyEUkteVLp
MA8NqPWR/NgUjEShMaQpw3Wr5lSZtgZorWYpBZ+GFXyCv66KpaHU7lEIYgbrC3lTzHN31TWxin+k
dKMb2Csp+i7FURPaV5D6dUxBA/GaFTfuxwq2EpzauHK6Uhtj8F5qyQ53bh5K+V9k7Qdsy2aHUEDb
NqqgvSM0K5W2RAFDWKoukGLaNVWLsjCNBA8TKULEiUfiZbmaOyE3gqksBj+6ZNDUy66pzc5alNb+
K1mef1kRsFIxvK8P4PFmmaOIaeOBt5R4ZpOamGFtqiobjp2SS99G/nPVrwwPiUGh1ojvwjtwy6Xh
3SzTLBtgJ6vMtGIvpXvjRTVBzIXKLSt8QKyjfqQ06FjSdoK72itW7ybv765l5H5WtOrIlFvhozXZ
juPPLnVSqX6wJGdStkfKsWReDzQWlpmwGQiLRtryHJTwIRPJpDXK0H88F2DRpmT0qoXfxUNOXFsT
/0I84Vv8g82+qCtlpjIcdZITCNeDc7ytM7P4H4+3KHMRS7w61UqEEPssfuJABJ6xvkePaESTQgAf
GrZ1oYBDn7L+VY1Jp+VMGeqMeGz5n0Y8V6mxDWe33Ras8r95vHhFUu63cSCjUTN51pZo5nidTLq/
alO5VmBU9of5bfbbGw5+DHuyJvR+QOgUGLtftyP/m4eAvjN6hov3c+l0sIeDwWi3oFLw8HCO7HHI
Fff0JPoW12oeCfr50uk9IOOdHMf0tIBXfFtPg2Vjx8TTdd7D9kd+wSpVYKCRrXFBhKxhNPaUE4Zr
JBInYJ/UHXw+ZAUcOB/8tmtWxUul7fukVKQCqoHFufAzJlmfsmpr6bRP0JIhuJy+8FbOGw6xkBv0
WBLN+cuHy/0fRapnW+mHcVHK1WcvllpVmAz1bobLgjsBMmeyht+evcdUgEcaIamf6pQ+yManNu3q
RohBHt6UXRGCvEO12rMIEVeKUFEBVLmQD/4Ng+bLFxyasVP595V8wz/mbI1Vl/odUv4RRcEcLzZx
RKvX/VECu1d2LHKyCwEa9P2OZDy9Qxi7enJDjqlQILYLvQxFunkiF5X7PV3Ej7y7LgG4KlvwBlxS
ZtbPYruLsiGNSKyurIkf7UrQlz2Ove71+3nOiCiwz5EAV+Ys9yzlqzMMHLxnxQpWAV2FPKAviLNy
wWmCJdM88YJXJTupdk/CBuDrDTRKFdWxaNKW6onjXGIIlJlBKmc9PsHleJFUCuvE6OUlt712K5dL
AKKLlLlyR1jYEPVNBPHmpc4QsyJMAi+EkgFiyQYpAuKoBaKz2DtxgamPnXMfB4gENkq0fwC0Q2Lt
wZMGcGZNnRLcPZ9XTTw4wm3pkoaqIDNyE3skECf1Xiqnpc6GC2BmWo7am1vsr4n9EFOWqz4TG7cT
WX5u0gIoTFlaFqUSHNAY0w6qUy4pRG89E8yah0jdn5Gg/BAt9wzv97IFQt3i1hBcaycFriNcUPdg
v98M6ZsPSgtB+s6jqUOrkWM655gYoPfOFBcEp14uu/IHLM6UqDymWQSAk4IdW1DiDzb8dBdKztN0
uoMRuqObafAPwCGJRWR4M1BQyANugI8gY2y/47pRQBGMiIA7i6wN7GZ4uTRYVQ6b8honYZhRohvL
p52ceulDbQpaYwhhdJX3xRuCtgckcv4fNfnjoKHIluhvXpSMeZYtrq/jYMwUw8WQgGponlEeuIpx
v60AnW1qtskJz0CYs7JdkJ+L2+VI0r/lF4lhGTKLtKjytFNKnZ/8KCFAGtAQY9jU5iTUCGLBrZMs
qr53G/IC2gXQLY/vdcJwlDMzrfSKrWhiJyWdZxevZcC6nziT6DUtDVwGUfDsFAZd55NmPvQsQlZl
KYCfP5AbMpSpCuJ+ENQXnNUzKhlRROFz6qfg/RGiC2TUx/REoOn4+4qATbp+rPTq4RAOPBrfsTxJ
yXbdQuIGfmFJFqVgrTpzUZ1sWyh/0+qMgu6zJiFtAyBNWcUI9vOt4c/w32buXjCCm1g8Y7AmyAuu
QUv7NiUiqet4x11lanVmuSWsMpqaquOqf4PLqPpxRgXEVsTg3BPoIv7PnQQ0kjSPMb+PVaGSWNU+
BHCVl2s/BM26VGdv6iocEfsnJO9UzLJA2VlDleKdTUIRjE4nFn0bvYAohgxl/VC00CbMZO4JzEdG
rtW5YTGjDo4sqfSUgHa2XJDMXp/Odd81CcL+8f2UjdR2lNs24wJ1uqJEq3HfJ9GQ1x8eZTjrJUpO
kLJPAVqdJWn5+SjGVFdkFiE59uILAeyXXLyrAGbmVNfdckNd9i0rQuzkAgZk1sqneY7jZMCgnBy7
yXPFv6ppA27bBPKdHad78dtrGFwVs6KzfzuYJlg/1px9iFg2XlcgIxhenkCaYsSphbN4cfUPNng/
i1CJeCff41DtHUGcb1XiJmBTNM7Hexkuk3ONFVEZCIZz81rLlyP2TovEQGaYGMFk88mmbvpNNExf
mxwmaLzhu+rR55at+Tjai0lzta85cMnOeEW0pJL+yJCJ+R9zgB27qbyZcDpFOor60XpG81BNlyPS
RdQMINb5slI1esQXOPp9cbBQO05hDXTX5cD8muoXuc/hO6cds62IWqosFPCJkDB5bNwaYhDKPz54
JmGTvUsJ0m21E92Zy2/9y88h0j3g1piCne0JMIn6NXWEZ+EzHKwDJUxLIsSaEzS9O35qEFiIFpAT
15KOzPES5/JTsp5D7jKgdg41zmq0z5MzmcjFMJ2ofptU05Uf17t5TRMBN/mSTq0tcJrZGSgNKTem
LEmOPKcCDBL5jfcDb8GEg8yryGnNqe6eckEYcjEhL/bbLcw65Pq5vBwYPaLugL6Kl2hvmlbg5nWV
CdBjFv36Pf52hjJhOoiXhHzpi+SqtIPXa5MNBPnd8RXKLRH2I4L8R2hkYGYNb0QUEYMrkJFsZB3P
w9lOOgdHQteFUZqWQmdKAlikJ0GnaTCWSe06GEL0TxPfx8Nvmv4JCgIfGS2+NHBHPxyACBqapaTC
Sqge60licOBvC/rNu52ibEO6qOge2jFo8a8fy6vDjcHxN5+sniAgCN3BjuTN6HXLu0YX89nXirri
qRjn9W+AcnuanbaL0X/P4aSlGyGisNYo6RxwuzO8Qs+oF5zerPAmi1I3p2AepV3lnP7cZT1h48SB
GsqNI85h12R+i1zZdUSQVo1tUFTkOUwEvHac/OE2fEdC/SxCUKgtG6hzRdIPPsKjTkziUOUJ55ri
O6ydAbcZRuEvurSZTj6TKO+lUvaXRwZq2tr6D/X8/5aeOQHNHSGb139cfuucOKDmU18U9ZsVBXh3
y0UticY9IgZW4JsZ/MEyudif1BnE1/UYjrKYiyy214uXlRmfHA+zontTnUlVtlILs4Z7HXxQ7MRd
mt4mXFXxb5U9qswSohT7ihnFWtRBAq50zwRQ7/2n1y/YqYVkrtfvEFucuas0PlOL0hZGST8bUEuY
1BllqKx9l08jDRhyG5DlW0Wq/uCdlqH7qeuBE/rCqS83Yw2MoR9/V8Fx/cE51WGlHk1mX177G4iE
gHEwS2Wtrh1+IUWzkYimQp9o8+hBdUhTod5/PZxZ9IP0/4rr2h1EuZqlR7oLSC4L+HOME+m3YMYn
RyygleSRqQl5xiFhioy0TKqQ2kIUSezG44bZxyo8UI52YUpvx81B4tinwttc7TaZZuyafAkvVk/h
jUZuwgZ08knPyLS6VRrtaRVs1pATTdNO27lIvzSIl3JOKqms9aSiRLX6IdD6RusN8CwaVIUit7zq
GTS1AyAZIW/kzQ/Vvp0jVEZQnsyYZYxVCSjTPxHzKSnFltcIZ7YBhxgA0wF5A21mntyZQ/8I/Otd
5KMxWcA3qJoWdSZevC+wYgIrgXZUsDn94y+cvRWWVamOVJ9VRN6YTapaZpKug3XpfR0RIAapLbzH
/93WADvSdhoD2Jw//j0ZCJZ8aNEQCAhHYaFzLvHY/HDlI4OlMu1VBoN6Y/3AlJauedmHwOKUnU9f
v7pchna5JGEMBlGRubZvYlBpc+7MMdKQzzmT2Ej31uTVK4Xle538q0Bl6ZAipZxVPVl3Hgn8+K2u
16ojnCrjJtBJCDrJuub+tUynwh9DnfBYNZDeDKv5NrJe8JLeGf/ms4RCFvA3jssve1Epqz+odued
91w5wKwpHLWDQYfEuySuTlrEaauVjQZKgRLlZ7z1FeYw2r5d/CkOJDQBpI2YSQVAJGLTOVaEiOzj
Kcyz9A69n0svZq5i+ocrWucSJwH3OggQbwVtHgHtOqNwNUhu5BAVgYgh4ps05kbxZuOSJCxTw0lD
EthROALIJYzu9t86t49Xi4UMThIID5lv3YbnIdakw1c0f/GNE9FiL00rYzuVdZzT9eu1+IHMgjrc
LdzJYLiPQhviUo8HN8tO89b764Ozg3r3aT8rKgBFema1anAET54n8UCsJLTieqx7JUyvIfDnp7Ur
29mSm+7HIDtkeng9Wp8LlI61GlrkYyPsI4cXQyigYFdaMhyqRKDCW/sS34Zxjz+IxqI31m3qvI75
/IH3MboWlIfEyRoGCfvNbmWOdDMbhpDBmCaRpZwDaf5X3Kp9z8JDRiQw/huLJ/wiEs9PMqEmFsBP
T224QsA3Gt5mGtQH65wM79/XO39Sz68DSy1/4HhHVYMWlBRmfPn4us7N+wjLSpv3Sfmj+EoqkdkU
nTAVYzwmFf7apHB4QkjhABQCaa2KO26IUi95tRAmaUjqYDW/Wj7q5bC5QNsQXYI9iHOGCbKZ4mOJ
USWhvqus89ciaj9wZuYcSPgcLdqDVbNMmmlzF6Y7/KmHsjXsMRElXoT89Eypz9eh6dvxeI16aWRG
pg82cImiHo2O5mxBckXc368usvew5xYFaF6FoUXg72srUXaicXX2Cg64/Fjywrsw3SEaAVvGrkkF
YCKuNNq3ddFb1xtDvM3TTp0nXBziJtqbsz55pLHEBeStb+6edKM9WyphTYzaOYqn0XfPmZx6NbMk
Seibo+Vu1ysFtLst3Ctg/CZA8Rek3p4Tfw2Dgd3IwzcNcJvIvJHs9Eur/pUZQB1A9rnj0WpKoJ3K
02gIe7AhZHUrjZrIjRZdnScPzEgwxNpiGobDngc4HsB4z4urLMGqr91hZ3mXC6zjxXyb0VtQeAE3
y/xr8EdLuO8Atno/BfY1hVPUwHf/e4Xuicx7+8MDHpcTT76K9XDziMswK2ZFGvqmVutxzgKwSoY3
d8IckgfP9DElSDBRs9ZWiRx899xsavjIcJsd04eu7SxzCFVIXeoDlTl62qYxC3NJF+k/7lwjpts8
sPFTMwXmrvDs08H+1NnzvG5ARfKl+7nI8qQDZBtSQZkz+1ycprgNPihVcZPzN561VpHEf+WR9fvf
o2tnsl9+DP95BYxtilLrOvIp/4cs8vryyB0I0BEkMYaL+ahpW8i+uaXkOCFaaQrdnsP7do2J7E5r
kU/NSueuKGicjgfp5LUt+f9jEqXm3W5bMzEcFISuw8OpbUpZHwsrTEsP/ZQSMWdViIQkMB0bKbfV
+d1zR4qxYsRiSsrHLAD0dAqs6XJVbZ9dFMsLsAruEjng4mhWB6p3LcV6ojcEM69UDLKeqR0vzz73
nexQ1LYPBes/jZOkhMrwdO2KxIvNGFesngXMmtkNtOw/ZmeCJcSvvVfVlKd8HueJIUYFKBvCem6M
mQ8JSiABxDFy5Cc+IBRkUn4DizgUwp60Y9U495KPXQAdFLdQ5/LocWq1YT3Uzx4ucqUF7iex0m2/
Y57FlSf1i54g9LDPIq0/rkCJS6Qn8KuMFa25JHZBLjPbLmBvupGRiyGAta0U59Ro/j6ZB32hOo+X
HaZxBq7hUrKFX5GWUZH8qMW+QuX2ASCJhnqth2knO83S41Vn6/rniw6HxKu0gXDTTO7UIvTpJhZe
HauboHDpUUfEeIc7axS5grGz71xaKip2anfm2U7ifMSxC4liasTqmWV6k5tGfEJq1ZOYbzU6JF9D
6wK1CckYTSjEQU3uDwxkRJ0iblC4XTeixXuYmDnuOtIUw/d9qqJqrnIPFJNInt0HPr64UrZgArIL
hLHNNaVXiQFlaTluwXnBneM9m6OqA2fpViQB3nRVcU2MUEz5Lu0wXct6h58nvn0qZ+qYBwe4Szgb
KCEtfHWVHEz8di3iLmGLJHbeDP2X0j1TAZGpm8ah7zO4emJ2Jc8SDbfLFJTmtqi7SbGiCJaJ4XVz
LrBtMob3yJVkTH+ndRKVSKJ7MO0mS8F41Qgp8XKbc+ZXnAApeHCfM2ykeKf7xiwJBxEQKgitm4bZ
veYPYy9ENCeNFtfNt/e/Hb3hDqGS8BrgeTyEagWN5xZDc6eIYFpsKBi0Gupi5J7EbrnJDR/fZs6n
A/293NxRoot3gW3Z2PKLggd8xgfCTdgCA9w9n2N5FYy6HPSlns89gfQuMTXTAdeGGC0syBTmlMLP
RJlVKD7lLzIbFvGD7ZZg/pLc7AqBe342qMlD2+przuCAOmI81Usp2Jfx7+UGHEXFVqRDMRvrnmQQ
GKx2CrNTLnO8qaQdHrG7L+MiTHHIudvkaYBJk4qBjVP8dnOjYGlBZJgJ9pqLbZvSqIShGOoRleZB
42XdMe2Ocpg2PCDUghaSoWWvTkn/H0nya42v/t14UXB+cKBHFAn1uxighPM1W+DAQgIAWN/iFxRS
MiyBqDYF9DY5zaQyXyaEdQP4C1M8JuBCajYipGVKfVsR6941r2rYABwqz4fCSahhQfy4S0n8ILXj
sr5o9ery2Ak773RE9gV/XZyqtghE/jWix7z065mZcyO8Agh3VvLdhO3a3qxVAUdflfTvBD+9qD76
QdRY+SdnS/+ENepoOGpwrcJdY+ehP/ZfPCREMxyDQ1SqrufzRn0LAhudKEOndSd0Q2Fk3+Z0I72q
96XGiIYIssaWtj7M82bLzWnPRUxmMIKav+IxCTrAzOFrsAM/cHJpWJrn3YsgE+7QzEQnj9MdjXnm
jaIOlu1EYAtCCDoNp51GSR6ue52Uqs4qoxOECcJj5wFx382Kfi/LmM61Lm12ILjB9HOael1Ut9i7
dO7o5ke2z4jHWWOOAGLh0dD+tGcBXKke9lta1mwcmRjV+uwL9u9Hy0VWT6DhyZ4olZK/7JNdQB3E
RPmbT4mu8wOB3psbBJrQKveJakbtka2Y99VZQUtGg0hn7Vpswoc8UsMdOooSaDl8hcRUX4h+1YRK
GpgpRaArgkGaoYLKMgsonbQ/EQbdwDOpt7kIrDvIZAxCrGcIqD0qRpvsfuGrA71xKBsE/Gr2m8U6
2PLmy1ASFPKCVTEznONEHUU7fQp1BM/Hemx60tlrsyuPJqTmCewiI5MG2FChf+Iahi3lQbjthZgA
z4bSQjUR+I/4mla/ZEDbP5ujSQm8o2gjdvd5fgFRcfsOhCjY5whKzYeIo40AJr21qM7FDkqmgJHT
PFFKfkNa3v/tGVOMAFMO2E6OtK3uyhPZdl+8FIUVFHjQK+m0t41zyS9rrlqPZkla/ydzRCQKCa37
NoJ6+IeuM/SaybEbWvQCLLjE8u3eoA+U8RI1GSf0yAaFjpHEWV5wRkCkSOWxsdho5s55sUFw5Oyw
raOdd/CeBPDNFbxJG5qlCPi3u0Tya2rNYHmuxO60fZ/zlkXFbeqZ7Cz0d5H2kyFe/h7c6+9CqFrf
baIfvdxURR2xx2hjHT6JeBl/3XwDbbaapxy/H3qMECc/+M35pioqjtvH2rnGgAZDtUYHjMDsCsf3
poWPNc+imd7H5X6o22a3M3Hvil4G/NW/ApAwmuojToZT9D0Nl6KEAoEBvwt1ap3g3wrPFAh0AZnR
+sZ+8+D0EhhG06HEWi5SOiz/bG6dGeNUIMgiiN2WhkfAwT2E2d17BufPxfFjQwcEixdBUG+b3U5H
+uzNVICHIVLcXjdj+6ydf3G+WoEO6ZyENft6/w5kioyfedvSEB/8EpKS3+mXRy4UKpUlbjhIzkyr
h4PeqOI8aEKMUzVRKFfQSAb8UR3oSyefuzzuaJ9CxtXxM4j2MDK09lLS09zuON2THaidHy2ULlv9
05S1iF2d53J8Q1R7O2dOsNylGG/KYFtzZJV+m/GpyeverVYminp6je5uyrq1zPY11QfYjyrM3LEN
H14fJ8isZaiXDmQACbXtIXgIzgoNezMY7NuU0kVGVYbVZnPK9iw2cLRMxcDIzP4VGBZVbdSQzMGw
36zICoGGHPm+qsPcXf5nv1uxkjLbyLBUfY5IfxPblpequS55izIcqxLkXyVIZ4oDfM4XkNoK5yGr
B8FXNIaz57yLL4SkTJMBAno4tS30+WbFwBlUxajy2gTtrXZPaP/1SSa5TflU4FRJqbrFiAIXP1ZP
zrYiAmN00AAYgmQH8hd8eLYz5S0DzBhV7j55yEGl9iwyp22748GpVWLLaUWZek3BeFqmZYIFPKmo
bQ5ufR3e1v4WX7GRYAxmDFwX5GeT26bi6MgJkhScHx8p/SBr3zlrOem6V8Zoi6EHTV2WdL98+3Vq
O6HfZ0pULtWPBV4uSUlKvRojNqB50aF8/ac4dSG9/aokQBLopvViwIIhkRyMFzfxpD4nccqsbDQa
867J4v2KVFv5u1ffr6Pl6ToGGzkbTOGOMW6H3lLYz9rMrxi/yJZ7S4iWvhHyTnUGgrPmMbXjQhgv
MfkY6sv2XyAMJg9WTzO1q/1bMXT/tjowCKLxeslQs002Dlvjo/mxOORlfB27qNBZQ5aSO7RPFv56
zp2kYbT94jGGE+4Ipl4Oeg+Z0EILV587Tx0S/2axtagj5AVnV+kROEiPlqNl3VZPRuYEEU06x+kv
fGqvCFmkWHoSW3/+0MK4rkzbEd+gsokuRKnrAvYSRNt3ZkFRfCb+Q3pHteqky/EeVslqabdJL0CF
2vRLEnmwWskA5YeNvjrih7dkO+0LOgPqjiAGFKSpysx+WD8NGHpLz7q6m1f6r8D5CGX3tjH0XhLD
MmB1NOvzuXZcr/jfsN6JLKT+/tKkxDXEb9rNpMBk5y5N+lgs99mvnjABirjGGtz64C92hfnmNTIn
wtxkcTtbYGX4KHM3n4M2AAUbsYGS+zEnyIDE4QpdPjTiNZHtljUiHc3GvnxyiyGf2+tylqpbZsXT
kwSmH2EzzOOg1fPrc+XAacYSGXpV/tqvbPoJO6tk9HWCgAOcytKWRUC4oMRLeU6IOIS4slGI4M++
TEGA8GcEBfaPKZmChn3d2xUKTAcTT64CpFcoKv4jrndB7UF0jgYcLdL1eKJ96HtEbBeefX215v+2
ThTJkQU/saeyIjYna9Y4MbntsrMV+R+HpzvWTqFTg8WaCg905L7N4cc3M0fLWiuT/ZggnEhB9EJt
lCLGOCu8xgUEW9lajZW+3Ch375U95YpZvP0Br758bOmBaao2/4mCV7EJuf2IZi3rnTPhslKsYlvT
XSbcC7tjohaDkBvhL66wYIGAcv7rvHMkAZL4jcj/U1vomcM9DJ4zr8qOHIgiLAymC4vnZX6CeWKI
1rwaM2nWxNzm4XJ6XvCEdDIkZskK78ygCldR/9GZzimgqg55zucJxyqDJPNeYD9ZIue+Okew9dgg
78ACnc2JUWJjEx0X2P1ihCOb+WrlNtA7hVbF+GJ9SuHjZnauftoRh4mYChkwJTYKO9qoEv4weFMp
pEqn21xBaWWZg/TnhsRqLwz6a6a9J7d3FhEr9/j4uugV1S+kolsJZkoE0TznhZtYf3RRUx7dUwiZ
vpBbQlOtMKHUeY1qQAbddlbIlGMRV2XTHUSebU20cTLLp2pjhYtxlMco7wZc5kE9EGiu0Xj2wkT4
AILRZRyQKGZzba7gTNmhI9AT71JPiNoUzh4Cyjzyy+Y4JkmP9uN/rSlWIrjqlQXvrWMRAUkd6pmU
01LyHKkiu/0qQ63ZI5+/C/f1tMAk6vcBmstdu+PWT61Ej5YGp7o0UFZIO9NhHqlhxFgOk3X9ocgD
oB8v/jwzVz8FhBogr56EFSPuctcMk9m3yi/D8Qst/ZjfChiDRwj29gdKEgk5xwRK2PSbm3Dsbp7b
9YKo1VPWik9HfVf2au0tbwcXizSkZtnTWpO16JogCapkz4YoK56LuuwfsGAYLBPo7BQelSsf6i5X
PhUseFxQ6iO7dfXm9KuKrJd4JUSAw0pcBVl60BCVlTePENSGvL0KHgfJJ/+vOuiNJLxsVW0YIw88
PkPKNffB/0sxSPdJYJb/IO/AoNF3pzVhr6xUzF0QZVvQc7xXLGb3EOXdxXzBAgdEYbily8WTIWSL
dHZp2/jxDr8p2bxcJFEf6GUgVQEJwSL8fAtqyuIT50DkMFAD+7PhNuGN8PHkoN6o0GiQFQR9BQu/
eXXWTK5Rtb4bmvReYMwarE48eBK2hR6pd8khfwE56StIjSsSqDdnm7VMuEbIs1LlwnY4bOoifq+1
vGsSSpU5mYKp4ai2p4OqgcgP+40j3yLu+NE6l4Hp+EfIZ/Y2tbanSivDnnbYMvb8U5lNfMBcpOD+
QjPFcqYON1vbqZpJn+B63cgtWKmZ68kRwJvsWZ5WO0/kUqPRwbOI9nvvxw0TNIVDdeivv3xmcnPE
N07djf8BmkIQQOmV4rfyYoyOEpDOR2OTIca8JFJ0udZ4hTE0MfnbZoURG+TCc1zzpAa1ozht4+BS
QwJR8HlXpw/OMQTA2LZ0ydM1nEtwPIv0Lf2AZQ1aFKvAdZ6EtLgpUlKwioCUdNWJNotP0iS9G2Gy
Usz9ctnkOStLtzRsb8/QJBDhKwRyss5W6q8muqAX4cyfPA2oXk4+lUBd4pS9+Wd2xqkIbXTWuous
IZJQn6519C4b+KhR8TKYa3wxiS/2ijKbnQccnFdZk93SMuUlF2pHgOeEsnPF/rNOIZ/lmOUeQnuF
QJvFaQ5ZCjbm+1H0A+IwUY7cPhrMexSOWlYK4Z80ohIiwXBW7BUJHODBjqi9/XppDbxDGqoMDEPE
iN7AaMN7fTylZKYbPAlyu7rZdTrHuoI95daqFAKlHS7L9J83JStO/6RWzL4LeXYlfT8yywzXKjKm
fqdsaqJTWS45Slt9IKFANrf2EZ4TBoOgzbVf3GiGAnxavSlSYwqscEjxhN3LPuYx3CgYMutLMlP0
yFwQQXwVSeRvJZyec/Y2voqZJYA8OqiB5zY5NyMdvDy5eShc5rUKx9xn2P0bdL+s6/jGK+i1VDnE
8exWx4CArsNycCJx2g4+aeFY82ABrs5kJfUDZP7piU0nlzzoKLUHv0QAuzNdfN61f241+XW1ViH1
XTTa47qJ7Je7aIguBYhAIuH7vTaBKoiVm+1bYnFH8oG9SaxQqj8uwg6zpr4Pxo/Yib97poJCRmqm
48H2I0pQdqBX5wv6sjzJ0vy7Cm1QVM0G/+OF4qyeu9+KgnBCr9hMzDQl54ctBLxeM8YtEq+S8UsJ
PCq1fsfAnjiWFj0AaYJnMg8hurAZGbi9gj4pLjMhDZuWc15ktaouS09HbIYRVj3xOQtQFWrF9dYQ
Il/RHqHbX0Pvryn9j/b1oFshBSjVvsSTwY8VCtoy6Db7eM+YlwykBMAPSC2g825yW2vIzXxil6a+
5CmsSnLWNpi/wvBtNJQLE5Og745aAV/Z8o38WBSnhkHPoTbRSzzyRs2TVxkiXwvCmc4JIAECLkwI
tOPCOVBnzyd6+lGmndfRugGHP69eEYhUpo03qrxZspip2scFaV+2yOzYhu5JUeaqVtlhLT/O9TDC
GKULk/8s18sNbhk8ax+3TtnuJArrlAMyWyqVjZOLUMVSOzdmXhSELVu14km8hHSOE7NaTr14EOi3
roSm0IWNM/e5HkXpLLVWUaF60QUI9Gt41RFJFKwKl352aMyM0KnmLkAuLdgr9BcA1iPBhUuhXcWa
O9SkRXjIrYon6So9JQmI7YMnPU2MNkC0Eh2wqgVGmRlrhxp1Ltzz+CUBNondIQ3RO8vIxz9RJDgY
4+2ReSG0YU/Z6xNnTv5zEVC4rcVz2p9k3IRru8ZOaMZbmB8GRHTpGpp5q9bCtkphYDHW09S6cbJ1
Vf7hyRFYG51NBGUE0bK3B6Ymhdvz0shlCRsEz+llUAeyyrF4u9QZbsWOnVdKudBklt12olMyHpl5
Vf48mYPX7I7g35YogxfQJTTNrzGdgLh62Zn29lob/zLWfJOIPG0yPWXROy5NO8GRrU+OO1uCjXTB
peq6qxfkroVcDOfUE4uzGeKfJDa17J510Yq1WA2JOprMoZl2S4otTF6CcS01jThPEt2pzO5l4BWP
2lu30jG4wq7nJDWLebymXZ14/FAu6KdIC0RZ7Zk/zMyKjGZ6OS5dI2k/sHI/yZM/g0wB5pwzqte+
G0Xl48ow/7iC5mGoeKQEuuV0Ez9sJR1d3iCV9BOkMSyR19BRDnTEk8Mt8wTZV1SzCxrvnBvOKMii
SNMnipPfmFxwy2Xx0SaymBLNliaWtBd/5L2WW6HYhZeSyHLpo09wdRBWCS9t1ToduWPX92L2fPRx
lgRk88uDZH6+0ASxWIpGGP5Gzki0gXkUv00uKH9pRf5Rn5LgjHqAvMcd9SZ+B4sKUHXiU8Kz+gBX
IE6lZOXyh3nA+C7++mkjAifss1kBbt9HsX0rG6W2SvUabn70kgWUE+t3owdRP/qHEvWkbgr1q7/0
WqAX4RZjs14oNjjWps+fny83mc2RVF5L0IklqELR8XZ02pNQ/700jEbNw1XauRdlIoqyHfoDmOXa
XJ1Kv8e2V4a7oUOmOjSBp+DZkjUg7C3234PLadIQ9nV9P7xPeqOGf/OvbhmnS/PEP3KB2r7kCyWQ
tEjIdA+uwdL9kRu4/XvnZ3emJEWk6dgEgZHKxCt9fH2w7XIYXUDXh0UjRXPp8gYD3DQJXcFtf5KA
NlWHXwhuw7p3di5plIYRYNAUZpXSmq4/ZWky/u/ZbR39M88goKvYTnCMIkBux3JDEyYjam8NRUfD
QudDSOk4ir6DvBg/Y0z4UHJZA+5afM0QtMYRuzq1AYySq3FkFOW3Bs8q6jVQeRTDritQIxyayk2b
c/73uJAsY2MRNHDU+atF6F/gVpeP19Ur8CWO5XhCNuH1O02pqQOClQqHRN179l2nEm+M+EJTKIdk
fpP9HNgdOKnaPHdHSYZWuDGjxzrwhxcpiJv8qj7xCD+DmbIxgKm4HngXjOODQb5Tmj/Mgx5Gte2J
vWYEovHayXxe3ODdpP2eLPcHR1DAADAJoS5YOF6eK4/NserMjY9Xt6hLu5gup+1ZhUOCBbVG3ZmO
M3jj1gbe014H96qtYcXIE8ZN9XsA2gMkG+AKEKMzB7fmDSaExjg63lXQ4iLxunkNcUvWupD2k1NP
xWo4LtGiFzsBxLnvWisiJTEMRSGCFunlO+n0WDPNq7B2jC1bZadAcCR3Q3Tep2caLr3FciDM4anl
Z7RrH4T0fn099x6LDnJDJLQ3+PpzKEHvKNGxkM5YW6GuStK91fdYrBO88xWlWUdywQ7QONehAtWV
U1HFCf+A7ysLXiFkpokvXzOO3ZSqx246hFrlH4LE1yQacuAyC04geL+OWGajdQnsHnQQsrb768DL
/2W7qo8qbDRZeRSz0HmaoWiR4md7VDtkzu/v4uNe53Rtaxf3EEkX/NwzJme2+o66ej2O/+BkQmHR
rd9+g9mZdx/oyWhdxWjt9etjuaz8YgvkFW7/izWvG0Us1RBlmkdv8QniRh/dq0ddrSqVYSW5Uo9V
RdjIicGpjHoBKI8n95/EoPGdUNZJF7Vlzcp+eM231hw0DRbT8Sp2vbdkv1/47Ek3Ht2sH+YfcodZ
Ydn5Ou96jjpivldofwrNEH3hQEkUaV2rvqbYzmRLUlnPBgFBvbBq6Z9ZbFHgEBWuCJowj92al72A
c4QMIttynvRMuEr+Z9fWHpz+5cxjWuvUxGyeyv7Kia4x3O491I1c7vVviV0E/8uEzc+ynz088Gr8
OnsLvfZtDo5r6eWL9cygAZm7VwEmzGKjzRLGas5ZthorlzgaMBm5qe16xEa5FD8FjtiDlggdmLTp
jy0cAwcSfNhVAeMHYFFYzg8od9cmUpgT/aaV0Ch+efpj4hbOdqiPfMMK6peToea2es0lJzkLmasy
tSmuseAZPBgaXTsMcizI+pHSi+5m0x3QP6eNESb4yBHwkls1PEcLuxRFsqHlVDRYk2GxYC0ZlLus
ToOj78WyvODZ5fbSofirvmX2v8CtXafFJl9B2ZfSgCxYBHeUlkJ9+G67njEXGLSj54CsQzSrwb9y
C73DRCmSteMmH2H7+lVSEckYvlAZuvgi0Kzp1d1cX4ea7LU1oRNDJndgEM5ebH+83CvTshjgmgdD
3ys4diI2Tdt6oH/b8++grwFBgs+B1JW+RNdCIN5G/aCkdP4g+lCf8sqnXttgLwozFPXBvIAylZPs
niHblEyVR2tXyCcfGG0rAZNXiJPcXlQNovRRbCAm4CZc80i1bvRWS7JmQ6lzWeHgpaNGQzokd7RA
oT0RIKPB/vvHO+u86MpWA13EPuCWTl9q6XXU6z6CAxyeF5xRzBRGlnmXewF7VW8ldJjWga1M4fby
7GJ5N/YUjOG4/mGmeqAVEAKtLtoUMxZaPrp91aWUJyQwEEQ1ErhYYCsXqjeWdXBi9d/XH3qRPknO
qScGnZeXpYHlXiENwX5tgmm0SJWdd64HvdcfSTFRmNso/riGNFut1N7qfoVMRcdo2JIbvV8FfRq1
y6hEEIbc8hIFl+1w5Eo4acMV49RPGZVNjh5oMZopNeHQwII6apZmoZ+JLRVFrgzyuYAyFnR+Lmmm
nbAUsUcE8OVXs2+vDoGGsdisnSuUP8clmxaCCPfQuHhJjoiWq3pcaI57P+xE+soLBEvc6c4b+v9i
K6CHYLDeTrLYO43+oCdGUNotR5VXHu02y7RFj+PDhZBzaCl3hUA8nhhUEVx5nWDtDgX70HKPwsnn
Ad+PNp8K7TcpHy67PeAWsgGBA+LBNRDlAElsYvCMwgvsNJlEQeQunGvWIJEpGebyJJXe1Hf8eqN6
xefmYNiOX+Bh59R3eFV4+U6jEC2udyrE9TJRIGa1+NhSvTKxYwIPycSb0UG4IN7TnJIrbzxY0y/i
2vqI4eHEyREAwBheS10Lb/nNfpriR6o30hBZOVez9VJ/pVjJGmZ45GXYw5tq7qEvvVoB1T32Tl7h
TTCRqOrB/+OhE4l+Z2JhMcgrnf+woG0kK/DeLPy2BSg7HsDFvhjbhoNxVabiktfC9aY2VXJk436I
4bEb57K/YNEU6KAKIlcVbwmVQTnOHXviRAE8L9L7MtPx6r9h22Xsl1dmpyDG4zAmjoWONpAmEf9n
R+0gU+3glR+OT/ZF4NwV/76MK6/I5W9DGyBqnw1CLt0C3+fC4S+UQYGjcHJnfzaLmLSMy1zSVIWm
StXmxf7qhU836xaKnWOZH7Oi2sc135oMzctg7gAjroHutoqdLfglvV8jTPrsUc2EM1tuJTV9P22j
3VTY3IQ3pTDXwtvZ+Lba8XH4eMLR5xt6mOzIgUSMz66Okx6N3O0DplaQ0vDlFQWYAVWZbWHazo6H
M0SCTiVilz1LXYlLLJooR4AmrBSCABQVyB1wGin0UkHGxh7bu3pLYiZAcEEEWrdV20No1YnCwWJe
j8/MlSCEMUQ+u9zofo9hr1dUidtOCC/LGvI9nvpRhd3IsscxUqWRkAQaNUe49Hd8ty0BgcLA0/W8
6S9SVs01+sRElWSYIBXJKqdePury/+jI8KM75jGwRWUBj5OY44fhWi9LcjFRoUGDB7Cnfdw1Gj9h
yUqGE57igNq1thUzKTIAQLAg054pCdRfvxe48zqcAudtK9oqI+xvpWtbJHCvZZ47aWZyZwhVOuos
AVP7ys7DHVmowjjG2ZnJKXU8jkdHQLSRdwUvAUFKums6RwKU4BovcHyJ81wGAkMuT5n5UYAlS1SX
cjLehewkIOwbJ7JGIeP3Yjbg+NrSQ3wRFd4n7031T8yMxYSPNYOmLpw+WN0iWIVYUFWDNJ1gN30X
56Ps/KfSHjkLZR0SBYXVKxRJoMuFqqcXzDId33VhDPiQXfh1cTtgAf+Ndm96QpKbPDjxxNnUo3fN
SLpYbfZBtVUA0vxBXjxlbzm3XsRyUocoailjjoGYdtmLtFyf7QXgUwtowxEm7yNudJt/WRsu6HwI
WAHYnhtah5y+mvREgTCxCDxWQLiNrd7tZKlL4Z0DCq2JCaWFT1iDHHPdMKtNQReRv04BWbqSPWJ+
6Ce3WdaoCLSPUJLcCuvqGnXXo8Zcl+YKrK4G+waFRoMfluKg8hwxOstj54qONuzio8PfpLvtTzre
HgNIVo9jLsgVLXw4a6cAalI3HAnFNZ0jJWLkk3XQE54JUa8CwdgY5E5bxDgWoA/q5/JwSxoVSAMp
3ghWsHinn6wBjRUQ0KWcraee6sAHzlQjbHUwzWfRLXKlOsFQ1d4wxUFnu8FNkPAQvtvWs4u1TOxE
uMxdjYuBr9Pfxyf/0U/8wOju5EegZ9RH2YIXeXl/u6YUGsRVv2Pe3N9ZCMjS2hOaI7LoXp4HBuBf
muby2c2p9HTZnimWbsZ3xCjOYxfAg97Xdc7y0p/j1aqDQZZpK6VXbCn3CuIKllNVi5uULDut12Q4
C3r768ZpOg/t+seHgflsWG0oNRvVPtRykF51MSfXPupMhWaVTtV2s45nAVbmfYBN3k0ohdwkAk5V
iprBL6ys4mHHLVY8gGWs0vtWKIaFZvYi7M8VqTtdeoru9GwPX/DVFl3cD8IGPGFxqHk0bYDdiJru
DP3M9R6M7/Oh+prcmtV89htt6MQgkgGZ28pIE/INLwweb2VeLrk1NdTdKvL/FJxQJrIB8tDkIozj
9c4El59YTwJ73SLIFP5xuDmNmWRLMrYv/jXHbV/e49C/GRroL3kp+ScIHJQpxMSLVT7W4aqQtywF
fqBZjhPp2tZa67IapvF8uFf3FJsKzqHcXHEGKj5COMWRnFHaGL/+XRy3ciCrOO0tcWsEVSFtCvpn
l61298vnMiofBIQcXop0sTj74ERlFG2BEBjXfYbI/JWnXo5nt1ukeSLpb5ZRWbxvUs4T9w3SNODm
XpaAlGsBx9sM6qDQwl4RFOYAVCKs+poU5UQkNRa2VdOvGzqHoSTxMCH9/SDom2eCdfCIGjtKQMYS
lQymazmXvohvDOoowOs4UlAjbCL0LaU6Z/9yqKFK7XTsg9G+XVmuj6sB0pnjdp2srrXKj9seZh9t
yqLoDtJyeBmfd2B5sd7RWNJ8pfkQjy6QR2QczE1Jq77+GvxWXvNcc/DXi0sLgNjyJg9kykUzzcam
CjpRMVfjRrEC58FYHosgK+CM3w2PWIRtgWG0bLBZGSiCluqNEZrv/WxXA8TLjkRcOWHj+2mjLA8z
i8LvuFiuwhRFKxZ1rjAuyoKgZGpEEbND/xsFdDbotc3mOCoABoh2VTeOBwhNKsMs0PJ1MijN7fPI
i0Mif3zSt1RAw3Jl0Nq32dhkbfcSWzcY+3i6FfwW3rGXTc3A4iKAJPHHHLfd577UOESCFqtSBx6+
K4OfUaXKydyq13ZYigVAJ3fxnl5VTudou6XdciHGM33+0stAsXJlfA6PSUw0IxIIcC3xBZN55jZS
fpPAjVuTOz2g9mvzqusCkUOluKy6c9DycBcmdlOk4zMUu0rgIut/J03vZuId++37c9l18h98Rp1t
P9NcB/R8Yw2+4hxOn7UY+0KvkGlzWzST8vXtIuMofRZt2GLf/FeSuPnlkoxAhML0h2dqt08mBrAr
lbSQ/oDJDc1STPGyPF0mKlLF2nd3NyPb4DVu+JJuY2hZZchnvggjIsdoHBi+yIrtb1rwvBMrXJeB
6vyhQxkXbBSR/FDE6vA75JTIYHNRIr7mSN3Q3XYqk5N9CKVSYJtDM/4Ama80kRlPc2j4nM1HD/Pi
n3j5WjPCIEjaHTGFZZU6VYdaQk0xYcUPld6pRU0gqnwYeU3VB3i5a1LRaHGQXHrpJ66Jkxu1Vnsm
UJ3jx1qd7jNNmUtcw5MBG4Ylh+32gni7X+PwIZo/SJJcU9ArIM8MlkWA+cBiO0wo+lEkjC0I1MqP
JIuIJhKCJvKr67S4roN4h+QVSAhS50XdY3jbyIGmuajwmpqrLDu5oJb/lyH+zdg6ii8ElJU9hNhq
6G8xT+rIcABXBzWQPXqhgoOsocbUUIvppQbnpF18WkyQbmjbCCVKj0Um/6XqyhRRAfUd115Cgb8G
YxbIPNW8bjr5CBgVhZoB8cyNjQ0wdT4l0vvkScsUa745MYA4NEQ79F0pmbckNGlvqOczyglDR89y
XpHOJT+w3/0pULfiJ/h1kj6oalMaZQHHxSFS3LJ96PtydltQSlpgt4VsNu8IRNeVSvQiy6jW9IXv
BNKqpjXgkE3IysziGKnJbCjHsUEdFznSwChLUHqLV3Yj3bTCfHozWK+w2JMcDkx3zy3G9Sc0YMnX
Z9KGjQrL6TUvFSrplz7PYELXqXHNna8MroLHiaHPrTUaw0G67LLcbEv1dmvJ1jqA+4EjY2waXY2P
DJrSsXVldL3M0vkDFhkkTbR4BSJCu2CdrYsigtGWt7SNMFXfaFUDhNE+Vp1lJRArzRziSVAhTs1e
fXzwY67qMhuj71X4Xfx6xpahyUrh5gCHiLD7vcLz9N7dPRFF0l5LLWxx2sK4pkJyc+O8KvkN0g3W
A1BH2KAIgJAF4mPn3TM7ik5FuVYNlt+MDIkKDVHN8StycSwlXlYQprzofB7YbtZIrnGkbTcgExc0
LnCc0JORxAt1PCdgnzTAvIKb1IuMPYRpZtl+0ZichzYA3xB5Czt3C4ojWyR5GpqmRbWHgyjVOvBa
FxFyxL3g3hyHEuZxcfDvUAnIIYZPTIlhEaXcrfG24brWp7d4vcbkfSkt4pfoYNGcfkQTNZ6lqV7D
28c8BwSXqTUllqB3R7oyMV780Uw7yW+cCpHtuJb2oIyElqLbgGBATyV14DQGAEqOq0jz0ZgdFXRR
sl5b6kk4Hz49lShv5Y36wibVpHxWEGB/sKQubXXC+nxO6ukTbWm7vGMCv5TqXtW9V2F09EVgi4KJ
52Be9dHjqttt85ooVEqyID356sJSm4ba7bz0orxWXCAeNUNgrBer3EKFkip9yN+jpbttNyUuZjqk
D++FPys2Mc591qlJ9N6kqmWM65Sns5vAyXnfoSJRRNLjdYS0+1gxUdNqiNanL7IGodQL0cE0xcwf
wU2Ga577SLk56/0Z4VhKhurjxO8fLuJCbCcbfmQ91fndDcs/GkebreCczOZeMHZG1rHMEFXqBOFM
/z0HVYkivCDRZnbsyCkNj4gtg7nQ+3hwgFecpvHiAe6FiAxnkZ2sF+hx+yl6mT0ZNDoXoE0efovs
WbNSlYGjIVeFv2OiIThRYdCZDW73yrTmBhh1WNsjD9yUbHhopfLub/vUwfe8xWkaoyPXiFNdZUP9
uqKGp7i5sYBvObWmbLMf018CM3CWG/FN8c0Z09q8kPdX6L+ZfQM5zRjvUxnkUdxbOe7bvD+zIA3O
VlIHjVTIoAMOkU7MKOOalEaEDrfP8yK7LcgHYyL0LLtS2dKrmB0kIutJ33PGRxEoU0HPiTNGJAC4
6ghAuS6n3NI+R3DPt3yI/Q9XCEk39tzjA7Dxb8Afwl9o1idVp2jL5ZWDET8rjR0/4H/hYEYwge57
jPsAbFmnJQb4TaehwcBW5IFMT92mHZkndcj7zedQ0ETklKzhs4/LXaU3eaXQygts4BKsM2OxjTH7
EyEIQomOrOSZs/vHValOPbmfdqlLzvk6ygOyp0yeVHuH6miBYesHQ/+eFAJLHhm3E92wH1ihRBhG
z9kP0i0hcvDo8n0yEAaAl19sWHUQa25ZVVYotO4M28NEsF6Qql7nSV98BqpblCQVnCiAH2eT91pN
CTn6hkLenWiZ7sQEBxQTJZGouHLbXHw65JYOe2l81r3Q2b9ByoyvRMs23OkaH58sLJWbGJjZ3eVL
mc83a5TVeF4DLQo4BgQCXYVNTByjxsEg1aeSiZx5ugSoRZB8o7kWEvB2vflbEiv2pfuDO4hTXilJ
u/j5JJSZzw10I6+PTLcUnhDlBwxFWE5Y21rz1awh6MFeTP6W6E1RtCdP4FmXTn1bwnGDk6h8rpWn
4W0RZ/J+s60KIC+f+lSvid/5dod+2ffz5TTkZA35v8VtpExI95rO3Hnc6fZ8YWfZ8DigL6WurRoK
hgdQqoTDJme+KQDfRGP7e3UI0zlFus5atA72LIJirjDVoaZ+gOtGCQVxw+Avfb7cG/BC5DO3leUI
HZxiqbbELpM03peGPXJmXYE8fIcWg7H7ea86pegNSr8rIhBZuDFnJqbpsf24RTt7ul4opLrQzkjx
BrnTyExKLhXYDosblvLYxo9A5Y0cidNdj3QAwLtN7ZQpIMjN+GnpwC57ty7G/G1RYuJjA2JLhmrM
A3r44itzF37wnRkU//MjBIsWGu9uE1Ssgg+UgNenoiVARroXotm0eSvHKcn5kcGiZqiHrqmNsQj6
JpsynHrCxzOwwazFXey8ErlvsYETJhI5jGzXKOK4EvB5+ACKjBZbo7GAfwaFIMcdMqDOBPnOCSpd
S1aD7080CmIZgHfOMOXZggXzGtq91Zay6gJ3hN6G5QoDGLTwm5j3I27KGhEX9zyVoivFyuX5I46o
EBBPH677QB4rPJe/r6MvWLaEaTLnEB+hYjl178DeHXuK5yqPTE+DAk0jn3Pd0gOoIk5izJF4ILEe
witP1tLWEaW0N+QLWvRx28F1Hp3FrBwMhezuMZn4jCxP/ZX+4G9N6XEd16WtO8vsX4aPSwcvAroh
U5VLSqjV6Eb8dnEve6oaVM1Jd6BRqMWl7iqHGBSdy5WUC72rNxGZPTysuXYm6jxpb4xKp4Qt4Nen
uLU49pFiXhllNr3dCxzipapiHPpujz5mm7JEw6TPabxmq4wLqRJB0ijoKP0WkzoFrjiYFNpJl8Ky
wlNbLlmfaKGFVkek/LX1QVM7RB7kPhE3qFJDow8jtisbx3fD3jY+7GqXwL+zY1zkYttiVqmLpWr6
kI/1gsLHunvyphyCRy+CxHqtixBqcF4/oC/zFGR0q49fzieUSu9pVhEgFfUN3FAucXCEe/G+eHu/
aFJXQcmH8yObo/Br59k6rT7yhl9FI2QXLpRjW0G0q1SrgqrRJZr6gABQB9wfU9kwW14nKP1/suuB
JVh7V03F0D9cHRTmqOvQiYBYfuX+uNFSH6Em4J6j7l/bqhrxZ/fCfagYYesMDolKXpMNiqgpqpkz
Ed4fz/xkSOQH9i+FME1b+KQ7frhNbnzKnKc4iZ09teQCrE/ucKFz4s4LLUyz1sSVdZXKMJxUkn1V
5R6q2U+WFoGg5nAAkwyCRfsEljyEcEGffAQNCuiy7+Rz6hr72szCD+Zqn8PhXZMrIr+Cu4DaxzFG
f9SuSFoHbFNWezG3UnV5AJQN/TyyTOJJfhj1onhup6i6FuUHdXwQOlQ9TNwFYgPbCsNVKn1kU5Rd
+qSTTHst9Wtq7tI3BhVx04HTt/qvN1HQ+cEg6YLl3mnKurkhRIrpePUstC1FNe8+tYkvKwHMsKdm
vcH6ShYW7QzQfWcRdL3fja3h4wBRunBHwg4R09rVShr3tdTEbmVYlpVNGYjVn4ywT+gzInIEXQdN
168JZUmpV9K/qfJ1tL6GguUPk30qPyGHAG9C1Ji97U89SEMFx3bn9QN2BG/mUk8GzwUci/HohFcr
LK9rCTxIsQcbplNJY6vNBzJzGdtn+2QA2PQd7cG0NmzkHztkyFbdrRJ2cjUDwof82gLaSeskvZzu
F7XLBhgdXV8Pz3xeRwLCveSC8w1YaSP/TyGEb/qPhj1m9Sq9Sk9exqsxvdviubRruefMLJYBD74t
mwuKrCJJmK3e2mp5bnz0+S6K5verJh0u7h77LmPfESSMTZAi1jK66IMKn6GG4l13+lMTz+7boLNe
HJ6k1h7g6E0zhIJKmSLSfx0hNTpndQeE+DQ4c5y7SzwHbVqun/LOxYqPRmZOrj0FsNSJ67ZpS+Ju
Lsp+Bb14iLAHBtjWEcLN9/6m9/etheT2GhRmPJ6vHm9HZsAtjPdpKate06G92/QaKonL0Bwp7JK3
rgc4+9zUtqyh0rO8EGD1VERKz43SMOv7N57KmEm89PTSczQpau2hOfv3nG4jGfu8Od3tr39AskYQ
fyLSWGFVbmvGEcxdKOGKczC16BjvrfLICa5/WN9+LEaYl2TlUXvvKaYCeldkhDAA9FZtMPJqXDPF
3hN/LG/zmtwnoRRtvprgZBcyAG+NWmcbVR7bB2x8gQyH5LE3CP2HEliZQfhkMv71lbn2ezKTbpqd
tifI5bSW7P8OaM/5AZydnDxKh+VBrW+wSiVKwf2AwDw8QGf07hu7gGEew3ViFB2X/DrUQCapuss+
hFe78nnWqOdCXlvqMmSnuUN6PZj0Y7o5py8xjWiNGIGFW1PrZIVEkyIHqP+urRJhyhU8ATbOdDCD
j8EEoIpWk9fjXbrRS3qDT5XYJAxbhRGFWVCJPnW0shoM59W6PEcrxZGetpmnSPeSHIHV9HlXcX3b
25K5pf9vO0N/GrdYZoc5kXwtqP7+9SHDibtaAWPSdE6s5E+3VjD6jafewLP3/mq2hzGsyy35Mf/U
7mMVykhcK6JPUvAdegiTqrpwoy5uLbptlsCKOERGKkTWrNZuRLdgWAg0I3i/TquoetFpw9IpEj7E
Op2DrJCIZBMPGkks5bs5zUAGJHgr2QDu4YD2MjzeUboX6XoPRWKkzcuAgckAJPrQkpls8akoeCQR
oK7vj2ly58XrVXnY7wk+o4JhyLid+5BbCYC7tKHU3m8No2X3VvYTIZrcIFl/E3M9uLnthPPzqSzG
suisRTcffBk3yDYrD1tgh57/myzFFjQM4SCpaCRr1sA7kYRoqdyE/cMGh0D3n/BPcgBaImSQktvg
pfMAhmqVTazPVfvLcBjAKmCzw4NtSNOWzQbbRHm77l+LsM/fO3N245rQ8c7XmXHy8ZGlAD4GqENE
DcOu7ttCUD0SMS9btr7cO4IEFOR9HJJjO/az5AxA3geOunH63Yv4+v0jqpyUFw9RB/TxsoBPnEIe
/ZRMVEe39QF8e/JAC+7MsUbsWhQJmD45NzcCG6c4sh7XCJY22bG5pwLFOWyqYRCbi7VJvHxJTGOR
Z6MIO24XMMaxMOOB8CU0uT/nBD0ET7b7laqU9D/pJnfAMUhztsqwUm7YZQH1VACht4GG/mOyu4LQ
2hKDZFHh3WBNo3BFoh9S9p1b254LFnofom3mRTCM6uHrvrRtBMlflm+UgxBxLHJB/cILuvzQOs8I
+5Xrnlqj7FTgJ6lsPxpTrIUsSC0Xz1maJ9yp4Zo6IAHg7iUBP3ZEjhJ84rULMr4T2g0Eu5qaujF4
W2xw5XjQ+U0kheWvJpwcceSkKe8F77SGtRh1UscTnpJk6EgyJjXVdXZnDR5wL5YtTs9tE+UB/lzR
YUM5NPPfxGFoXhxVKLCDV+AK8KlChrV7AUDgiexXqc+dBHpykwz7xb8csVDyVAu7AwZ0tdRi7byj
qP+j9VV7hbyljuUL3hN9TFNdO1DBaBCEqztw4uhZtQAlV0ikldv5Dn1BBQn49A/ha4bMHdqRjo+D
FEXdg6gcE/37RAnHBA7tgDjOG+tlixqyYURaWo4HVpR0M93THxLWwz/GagAk+pkBW70jDqam9FkD
r5u6MYAOYo3v/zH8eUsU4nhIQRMj84BrOnoZQbY/UrBXZrSnEZy22nSCbBtoV/anx3ChTggVt13K
67bl0hmscGjvjfqt/eNxD0siTTagadbL7sxsUoJPEQ2M+cLYPTrrqx5O/x5MKfghxHUBDAooZbHW
sxr5R3gGA2lDYIm5zH6pEXV0rnc5teN2D63ZsmCouuHrIMYxtd6OQO4JzKZqEyusV95z0pJtiMrf
LP1QMANHVSySBLttMJYP3/oY98uQdNLqfJvGqqnXuOY6MxadL+V0HCJCDVMkcP3z0pecU70RHkeM
8Hz8y3hena3Q894Qn8TfBdMl5iaNDylNUlpOEOQs8RjoGDsyY6ZUICpt1GkN96Lc2dgZaZGP8Vv7
4hj5vYg3SQ9RbXElcH2w7ls9dburTZe9Tb/ypsM2SRtBBsIR040yGhdumnssa1P8LO3dVIAJJMct
LEeSA8vDlGg8Xbb4aaN6bzUf4V5pRydiLnypey+/Bsjb7d30zw07XFV7h/HuiM68iik2gLPKasF6
LLoMBQeK5xzIjZhxnn90Vg9Id8o3oesImM0krd361CP3tGSsL2R8tz33WlzCDlvHApzFeyy7TAIe
MNBS+zLns4nj7Waq0luEYF+H7wClTA3OpsrLvCSGROFGghgmtkqlLIGRfF0zdajcOKVirZbsFdOC
XQ3pfeQip+tGJIt/r7La2sB3wZEIJ7cLhgUXxFyTu2IE0bvOfdxZ23U2ZK4UpKALX4KjeslR+/G0
AcQnIJ5ywd5wKM6OHoQwcjfArzVBIECp0SRhndoDxEXO3pmXEwFH4vCO2e+dhry1hq1RhPLtMNF8
iZ8cufGmNb1NfTQoi88EOb2Ungl8xU/NicISoF9oCM7o2yoPafXW4RLrO4vrnVsJusJKFB/NwFJz
3jsFfzrxyELLhhA2bNs+3uDppG052Du/AigP7BPFVY5+EwrTw6LMJw75EbpUA6nXCV87nv/5fC5d
kJmFWcRFH8qcNgfpJYNEk/l7L+A+mD74DdkKQFmSBShvbIp6zeXpZXcNfmMGLwltev5tu5KzLe/H
ZitE+cpD72J9aLL6ppyJBG4Bt3vUFs60UENCuSmEwyx3rkvyvYt5sBYoFo4uZVrizHtiZbTZSuTq
IcIkMFvxkYoEmdDi2ObBOCwz8DYtHc+HtCz48pa5lamVBStFuanafbKAsBKZUt9vchp0S+75MrsG
NXqTpZmuWhPJGJ56uoThQ656Zf14Yx4QolAkUIkH4Ry4tQ3K6iRcnC5rvND566bRR3K1hSAsgzla
vkkJCbP5xiwboNNjYvjwfZ1cCVWh0InDFUQXDneS5Jd/LuMxIEpnwIwKB4hOPoS5zMHyQbl2aWuF
X9i0DTXejJ3h1EDEEVHgdp7Z5Y9bSdHyISR1l2dbfvmMPq8Npeenn7IlzGCb8a06YBQMEwbtH1re
04fDJ/rms+reuUp9ipbgWY59PQSFIHLJ0X54e/wlmv2zgA8ifmaLIKipSSEErWMYdymJ3RUU8xDY
ZtA9oLq0UL0MOXv3jjlN1a74tUmEsvHyQWcITfB665SRI9NkH4iuv+FM+zE0o/D82ulcd4JKCUIJ
0/Vy0UC3l8e/tmKbjxzLgq92KbLrj2IE5ff1TvFyxTTkQxmo/46JHrX+Z64h5h8Tlt7tZRHCRYEc
Nc45XWSuZBn02ZOMd0dbCYL5+KxnIDQCYadz9Va9vmWFdX1xsS4LLmrFcmZdd/i8dx76QWT+GcfK
1Xg/pv0gTySoP9b42GGsyWdtKUleHArHBHbxJE/A4vzOB17WYa8SiKIDELNoFoNYRP6XlZsIsvp2
g8ci5vJnrJNNiUAE8Ox5HCs54/04H7hGHccLJSr4rRj+Xb0ESJSHfNJ2YaXtmmtK3c+b4yIdOtgQ
rq1fAEd1xFz0F9i0MTwQxVSznZTexd7S4ulZ4frlFgRuc0ui0va61d3nAjYB3W6XmAF1IZwFOGKa
AvTtu/hvLKkPe0TmoIjTKq7IpQolkOW9B0U6MyQdUBKV6qlTQBmuEd+JvOSpZs3RjHSwM5SHmJOq
YNmVXbm6RzifuO74q+7u8Dgq7RHvUbZO4WsQElyhxd9ke2YGg8uAuGu5My+4HWil0JSMPTtsME4p
MeMm9OM27e+oi2xuEicAnmJNpXPyhEJChY6qTTGUdB7CtXGq5FjuBS1efVAYbH1prQUiVn/C6HNv
Knvm4HzRb8p4xKf6vyT8fUJGBxvzPbWtNx8kRVFSU37VYnUwuPBQQKKR9glKC3fsSor5RgzV0pYA
nLqdc/WL6bEEHG9xEabTpQr1oyIROSHcyK6hKTwslmJD2sUm0Q4lDvSRsAzE0BVzWayPvV79ywWG
nNesiJ4zXnIAXSjJH2eDUMCc2dSlqN5jPV0pS/cfB27rv/utDfL9Y1U+t9fJ9vT/YwZHMbxz81Fy
/sA3mNvJoTlOAekrYhaFyMiLydBNJegl3lkTQG0Cf0/lTl3nSLvl8KDc411p5FCLWolgxbOm7s3n
+F7Rob7snIoe5MRMT1xSgXTM5mz3SKyQz3mdei3XKWMaJ6gar/TUoBlZnGibTRb1JIKFSPsE3e3H
CEUjxZjmfv7LXV2ZI+9nn6DfJ76cknvhq/dw4VZgbpJrF2bBprxOeeVYycnZRydcHbk88M2rp8Yy
S6eJ/nss4gSsFny5ZuU2kib09lthi59vZJk78377gAwRnyyv9PtXUbB/kxOHAa4IN4WxrE3AknMz
NvYHB1++Qc3loMTRWvFDSd7RV80rWh7DxizB6sl0g+fp6Jxgbw123au2F+JaZTaoJ5HnHxU7K31Q
FpJFQaW5IOrjtNuRJsGsZgYNC8KG7opjTgHeeSeQ3ZB0j9uMXPpmgTRMDKSODpN/v0fwHW3TyQZ3
KX4ZcyNZXcWZN9lzwCND1n6d8w0Y00JmFbcL5nIAr23c8/jm7T8f5Pt58vc7P5NiYXETRz9jD4bD
rDsVqLGUOOcbBtarLGEAmptLPkLuFS5l9Vv/FC63f0526xF9a2a7imFz46hOoXxHSViVbPRrwD2G
/LSKMgNYGzuoaKqxkVI63AARO5/Vx60JK14/E3zYBErRWhv3WT5lYJrO9AvABd3ExTVsnzzjqpEn
FUncaTPfrgUfw2fqRheinpAHC8MNCcfdHJsx4XUCmCQmDf71KKVgWsdLNNJXqYJCzcwCLrlfefYT
aKq8uEZ4+XA7vND+mLJ8dQB0+UD+2jMoCl/7NVAVjfOkrQErej90R0WIVsdOQEwrs2wbjGuSM/wj
+F9KOQrwgCcRHcqFxeUu80kT/wwSBkHKYIawmNY21Mntoe/JAdUBGf+T8jkFGutl7H+g5D3wVIzO
cPjnl2g/KPwTxYcbQow1ZGg+Ya1mxQQEPn4F6P0gqxQmmMgY/60WMcMzvjNsA1FG0whE/0qwmFGe
khlQim99nDOYB0NVSpCVdyc/wl4jh2eZYHVaHJzW0WNayvyLaw4lfnFE6ysSrnsV9y14gpEtbfev
2ioj72pWVglHOLlVQTGzHJ9/6BTPJRujRxDv+HX/PB8GubT1ooJcIbeSpLrSZwX1iGiRSs0fSwEF
/0SQzwq87ZVfRwqIcQ6BV38MlsdPfBnMqyuVwqNvoE4Imm7NNk6a+xHahmlgQQyki+iaqedB0aXD
FgWma2GGSCDn+GKfAy3ELXvRRJ2ajZDxDXEF9EJnN8gyuE6EcT+dP/HSbR2LUUkqkRVZmnFKMqnT
47vU1rFpQEoixosZWYkpANQI+LCmf2QoVy3vOrdVOjhF01sRv6GxkKS5aKqpo0ClPF+lUCZOiw2U
cBlQ1/1owwt1SI+lJ7F9uwhrT3cl+xehKIgDhe+B8141WpJyRrGWl0QGT0EKNqFOUwX+YA4gl4yZ
lL7ooh86LHGgt5OppNdglv6UbYiklcdureIcCjHjIr7RnBa5JFC1yrF/DzoqH899uOoaWpbF0OCy
nwFAPSWQTJ5pwxLJy0o7hIxFf4mYfDlR+YLX08Pb7L6V+c/0w9fHOSRjAiDTUEgorWBBbpIL9BP2
/ORghUx9Ede7bgGGw3ElZWTtrFwX6pSCYjQFh9IkERuXyWPX1IttZ6obWC3ZPwnV7LPt5hvBt45f
09pVsP+KTta4aQdSDI/PwVjbxkhgk6byLjL0lZLGda4fSwwooTD2SfGP/3Zl+6QurwhlIhX20b+F
vtwAyF3d623Ughc1cKUy2/K9oUlgXu4EUwW89MZY6W4Igx+EkN0Qd+U2hl5n6VDMN1VXNKz1A8Mn
bHRRbJ8EDeG9MXQ+SI8CRzMkZIGjmhBdSvzmxcsXvgZG1gI34vABO+8PbiskUitczAaGcCzYX9I6
Yw0CLofTdLUO/vUC6JQiW9S4jDAxTTxmK/39QJ/ganS1SpGviLKL4JrHveaBHOgcjs1TK2jryytX
6MehSm0a7IH97jhLUL96iu5KClRCVuO3oxLjYSBdPDkPtrA9DIjK9nFd4PQadLw91v0SY+mQRLy0
cE8eggzzKNBXbjQvWtZQbF0wtNwlUQY7b7jOGgsP+AOyUvKrChCRX86rmFnExB4+E7X7g33L8yPx
bxVDmaBCX+R48n42VKVQtho1gfz2315Qu2LpEPbbsWCUEZye2N6Yl9bN1XN0M9m5+nG0dzCO1w0A
4JRdN/BJcOUu/UnxxvpmYMVWxGDuqdreOWfNRsKC6HX4AmRNH8SIbjlhmfh0i4JMY1XcEcrqMrXU
FLepzZHeWawDMrJpm7HkGfjjf3Lv8h+BIlF5khvi6uepHiyZmmxV2mhuqUvmBSyBN2fDDQYuAWCb
upelfP9P0CaH4JmDuoLIDCIEFZRW6V4481xvQvMx6kegDqfsdwnHkpqsXu+fQ6xfnIUyJ9Rh+aN6
pqKz0crXnMb7/V+itZMpX2+QumtRIBPdOkog1DLCS09MFocO9rou0ZtnOogPsJxszTX8B2l79Foz
8zO3NdszCamdfAXymCDEsTZ0XDJLnJSYQApXgssLo91UPYio15+pIb+XrJvIiXTk8mT6cx1i8pgE
FRXRQn31ZcIXXXInQPVD0mab8WpSGxzhvjgb5UURF1Oi8RbRxDbIOuY/kIG8jc5maVNnJvXrGJYE
lZTOWBCrR88Cz89Ik/bvI8o5gin9wukIgAWp4VQ1/3JAlqREqrkxnhj9Du8gu7Mi/fDbhgJjZ4/t
Lcb84QQ5e8xLuoFxL7TqQSnSPzn1kD4xrSlC7mWqaBHP+PYGJgF+vJu6rRCvT1dy+u3l3d6JyDA3
lnWnD7HIPIWCkmpNIrrNR8L+/Lg4lEu+QBAjNu2dArWyKvAURVQ/ooqb88n6Aiw8tVz5kAUkEiK5
6bs6p3E2X4xtJW67TLgzSgsGt826z7686FAeG2kpsEeQw7dqT8Fay5jgf7+Nl1GTSsfhBeQ3VyYR
12kTlD4RebXdkQNcBfcBgmyznAvInSRBwpu0/LUOdYWoqFox9a9UTeRV7oy0lATLPuAFUhl4ttIe
0pW/+21y7FM/JyZzwSBe/clyXAwq0YwkCvcx1UqRM+OgInXikwH5nGq/nfC563xiNbwRnJQL9S27
0Xx0/MNcfdscM1N+Ng55pcJAp1LFE5zecMfZV6GYMXlN27+EihbZqCiOzRIZvCxfRacTUh5Dzevd
xujqFcP8PlxL3w59akM9cNO1kBJ7fhDqOxcsj+DZGSCqwQedkDDao9Bwm7UHfD6gUTtaskxlnNgE
9C2ahOM6wG/7K22YUsWhY+EC9GDIyYqzXxxoi55M5DOUE4OiZal/ZrH//Jtcg9rpuwq3TSxL0yt+
/trwtWcis+8jV/0SSrhPFi6r+33B/ArBsRAnXYbP83gDoTqLDyYkdYf4UnfXqJe/+gMgihrUGEBn
tdUxaEkTegocpJtwwahjVKpkVxmj72ftW9vhcKLHmIjU5iL7Sj3GzMD5R0KpRkx9Tc/2sPhMyXmJ
ufMDW/0aUqg0i3gHFg+8iGqNWJg8daMjIdzDGM/aloFzg8xfT/AYdSz5/WUXaadl2pjboqBJaOSH
v2NUJi5htCdfyZFY1chdQFyW4+ETRVGkYLVidmDa85yUGyavmsFHR9cJD1be+p265RD2JzT0dh0h
Wthb73ZZ8xibWAbZ8zuJW1rQJrzlQJmzTa1JBISzRyPDi9z4Bypeq8YyRRkv0wg3GBEfJqxuQWSJ
gUPCDoqKBgdPhTgkBMpEfl/kNEFqBleXWO3jUqC/1T0KiYRkuo02k82G2UcII5PsYlg01fpFM+8h
qLkbNMHXpiNwP4FnzGahBfAhMP4I+Q1U8ppza2FirGuAf6ddElEOmWP1no+6zNGuN1YPIEuPZBKf
nsVii9OUzz+jmZwDRBTSAySs77lt705uuglXdmok3eW1IZpeXuiUQskQMkDIV96RjE+dK3syQV/S
AsiiRW1OTKJDSZloMaNLIo21BrnOlH0piAVQOn+GgjVAQ/wiZcxp0JB7lBDkkpu3uU+Go9a/NgZD
vclfTdpibmKe5qiNJ9BFTylsqDeHFXHT5Ec44RCw04EYI0nZLk1CqELswSuQFyIcrbWkMl6zy0d1
9sKm4HYGhtRxOocW1DFD0p/zFqXE4fqrzp49tAwuiSZsaGG9a5yYNRpfiTthUBlZ8i3COamiKt1x
ZUaAQyAzpvOTLKiv4CT8v2w/SznUmA8ZXBjfEYkmc4WWKBH/q5BTwi/M256vNTABtEUqdxgN0doU
DUwAufjrU5XjX91z3WzmzuOlrnjb53MbEcv+0yeMbkFmzk5hHj3JESiNBwC0QridryF6n1jcIaZI
CxMiqWj6GyOLHwNUJo0NT1INehol2OHxyLEWl4sXP0rEKawkF1HNxVNxpODWP0KUn7zTAHIDq4Fy
8QAKEXN0nDPaxgkA8fS4wfDCQ5pDEGCd71EPhxUEOUz7lCqpWk1HvzayeY07nAdaM8k9JzqBX97m
tQyQGovuNtMccDhEWsNTf7UsLFW1nZqtyq/sFXA2iBoK9g9a6Yfn3bqeUxEdPDfXqLrBJH0hhKic
7awphoIQk0YpgiAayjehFvtJ/4lJJMo9XXA6maMgRmranQ8fi9jzPiH5Z0ZlY8jzb4tn/Dlm2YGY
9TMkUC9arh8I6hQycA6uLyn8eiHpvzcFToOJF0ZDwCI+g/3w3OEZ/hDRKuGc7VZny387tdTWgZhi
lbz4+rua8KwvtXBwO5U8i3J5+bwUqfz+Lk+/E7+Jgt3+XO9ld+DoRazMTclQh5AL5j4y3RUtRGsM
XRWP/i0YlYm2UiU8xHpreINZWs9szFzYuUIefoT23MjedxiPMV/NnNea+5PMOpQDujKHtf6Wacd9
GmVwWCQ0BQnwjxnOVQeFHiHNCY4MYEMRQzr8D76HRIbj24fWz1gNCWOk4tfNO69mJuVgzYSMxGz3
MCQzRo2TGEmRzUVtKuPXzAZKYBI3T37VD9MQn33CIgrZTPGlQ1G3WhgLa0KUH3cacgNxSLKJl2Q/
U/wzcOqh1iGhe8dDuJdWb/g7ixIKcOCqnVbT8yg+idZgBWfILUm6Do5X1BlP3+bDshm16fq/Lk31
W6B6FpJkHT4SqqVocTY7FgyWMW0dVGnTlJ/rYqsiE5sCEBjd5J5IPRQ+SfrsxsNisgwOfuDl5DGQ
98v5Sw9xhKcAh3DjbmOv3IvzccgUFdog2Rgey/yaaPur5kgldKfs1ChROv/CZTMqTijvD0tK/SyU
C4YfCZuQajSQk1KEk8Qd2mnsX5QocLauVDZw9ic/OcT1DIHWWnX6ej146miTMykTpqwy5KJmXf+7
4hUmhSPuPb2ie85KRPWCjpVJIuaN3DZASMf5G5ijV4xY62TDLYJnzJn4bnWMvxItqIRY9kcNEy9J
6bSp0bIqR/t2adrCqQygd6NOrBgP+dslEGNhMLjCo3sRHSYQyw8x0NykvUX6DxEhlsalbPIJ9EAO
zhTIiZ3A4KJ7DoHBGUm0Q2uyGOYlDGDwBYWlhiFtMO6qZZGIRUa5ueaEqD1V+A4ysfueWKbRwtLM
lEpGCBIdiyOq0xZtvsgH8Amw0ffDH0tAyjgutfPXcMEllOd3X/1ZQ2IVs3x5hsbucgZrUzM6PWZn
VUeTXqeRctnE5jgSgvnzGZoZqzhcV5cjh5mZavCIsbyxfTPB+89ZCBZIhc+YI2KvAqNdVtAPcRda
E2OF6tEZCNB3cM6+vFsU+kWoKpXFf4sMsXFoFoU4binCS7iUQtwWi5bwVtiQAKesYgLmHfZHLKtX
1nVne8ZCwDpSoaIYRDkNiQcpDQBLZAbCYsIJzSz1DUKnpbsIolZboLJqNzAjKXL4eGCtRqUOo7rj
da8Zf6LSl1x2oGu6teoFRBAXkCKtMpoI0eJUEEevtCE/VnqXft/78hivPvsSXBFr9gR6jeUWFnF9
sS8SM8qAZHzynLCPzomNPWkQ3/d/vCNzKZOhJPYZrfCMnW05aHNNN2mk/cp6s09TixFVIRYuGJ5L
icbMQlhQO3sz/qo0vRbbBiguD+UL6emb2WEEKdd6m1lzqWwqi7w+PrW9DH+fQ8Ry3WAvDmqMKDH0
BQaCU5IcWorqPD2sHdaleOBMiAAKQsOoKcfKfVJEL7Gum+pyNUe2VAX5Va17k1+5qXE07nNxuYpY
gzamqHsQ8LtQc4GGxybQWD1sLSlyCZaXt/DM2nUpazGk1BYRdNpMiZSZDxlPCJEDIx3f80JsySOD
PdKque024Jhe6ugv2HuCcA/OL+SkQaGa/WPRCAYDUzWvK26724A72jhophkQ5A+bAsibXJM9unGt
3303keGcvScKyFaHEEBMrwQMNWY9jYlg226zki6p2Dgv8aYoJWf9zlyb2aYHak1/HEJMh9wM5ieT
IfSPnaoefvxsyzn4dR5fRk46vazauzjD33dkTi4dwrZuDSjjDZ/3IhwOUMjVwtrXmII1WqmNhGhk
a9AXW9qw2KxRlx/tnlXPsumq9NgPyOxj0qhe9wpsaM6/YfE943RvnK172EC1GXufS6O9RcBnH4h3
WNJjw5A1ZyPwSRg+WmrlBY6Kkeg4X9mKkt8vGUSrH2yXbjuLtj4txQXa07aGG3OQJS+7A3ZPTHgr
sq0+ko0bqMHAX+FXBk/MXsl50e3/DVqSgKzEbqlpC5ZD/C5etheI0r1AA4kqxskVRVf9xNuL9CTh
aCjA0g3L4okWrVkV9eWTEIJ8rLD7wojdmx7eh16jjCxkRo97loWaMC/U9xsMtfTCqffAQzsuafFq
6p19rbRkB9x5zOubis41wedT1OrL76gzzsusstIFWKZYlrB6h6NyNmrmkcaFtb8DJwTJ/8CftEBa
B9TLkYKOW6GU3ZFflwPaxwll4UwZ3hqeui5Hwigee5ruJLRdWt3PRZASsc0yZy4iXBYU7A1oP5rM
BCUFp1f6r41pHhiSRyLOmTFgKVKXsXhUPvVXexIJSyJTLNA7Bt03NjHYSwhwoR730/V2jqHpthMR
+kpzuuYZqlwFYgUk4lOZBBCpUszxd9vqLnD66cleYgCk/86y5UQpATDgRb9/Rcm8/vBGUe/8PLc2
YYkS9ALWH43FXzSU48umP45RPSZvB4l3FyLgeeM+ZzVfneeoM8CR0IbL8wY1KbrHaYnremjN9rr8
xhcKxFXIX7NHYnGSxqfKGC1iUgvBPJ0U78XTtIPLU6Ep2o4MWvwfelpguAfClAD9urLkyzM+eWlv
QF2KnM458/pcXpPU260FzdZgdjCvPJ/KaiLXfQLpAYn/HG8v+ThFHpdjnMT2B5XkpdK+aS5YsyTY
FYjowzjZrkmY7fSR6vJ9fSTNenWmMLzOvcdrqLgDttg23tXAjImotI+ScKcJpA8ZhTCYGR9kF3Wh
mNGnD1/TvvV5RashBGGyfsTAHlDUJDH/ESUScJbm0YUCzijde14iAFqnxV/2U95l+GoNePYo4yCS
P4njO+SkaU+OuIgk31w4DiJj4bQ5cnNQsVLDPJBGHA1ywoEbeyxL2vG21/QvM0TVWmii+58z8Rtj
ZrABJ5vXYtKpCahxQIFLWT98NKRXx5OgcpyOvNdBkMlIx7TozvOv9Qz1+fNw5b6eAoigZJqru5Yb
C1ZY3nldApGx77CSh4fvER5whplFW+ppg4xuz6d07FpnJZwjHDGcJSSky06DG4exQ1dGTDgagaQP
lKXI52esScGY/mzMEpDKixANRK//Mkko6+VvFrQ6uzhMINrne/ef6bmsNh9Wdz9lAsgvGEo/D5QG
yN2R+vbDXWB3mLW1qsx0qp3zi7w2biQpBeTr9tjilFXG0uspPYE1tbJw3QMkRayU0Rg3c0AU9ajZ
KIzdo51fTCdliqQe3/oSP7XRlt7vfiJJiatDFqOTE7mR7N2U6mgbMBktLCaBX0BmUSj7abLRlDbL
64pNhQ8ixG62HhL60SJEUhsvW0uV1XMo3ZzGQGMkxCH965AzbVOH8zZ/PQ2wt2UDcYIVccyZu5P7
3m9S2bu++9Kh7VtFT3QCfKfmvmWzc2UgQYL7eQ6AXTeng4oAxqDvr7t6hONZEmnLSvH5jW8XkkiG
Eioa+PI6sdf0dWqLqOir2rcHFom/PaTFuD2gtDypAzMJ0aks5tUgxev413A2hJX7U6zlj3kAVuL+
AIA4bO2ZLsqE8jwZ+na91qMIrJlmz2f19tRnvh5SOx0DV32jlBfDEm5Iyf2HWyqWG/p6ELEhACX/
t8gRLr18sTPQq/aiIZa5jl0YNOz5OFwWJELiFYVjHuNxOq8N1GrNXQWE/u29TlU+fnptb/hEj7Kn
jFDOJ215B5gOe+JyDDXlMTf1S9xnE7HhI9p1Uv4F6aTfHiNgoKewwci72MYXPW3XF9kwP52ROKh+
5SMHBQrYjR62Xsa6Ikit5Oefrftq80yov1ndTDwl2NdbX4htwckqp5cHmCpSbMPXz5nv3pUkvAeJ
BBhaTqF3zDY2QPIM8dMI836hSDa6a5+SsJfjGFLz9hYYlo921qghbZ+O5K+hIeky4PDpz/yiLSvG
uqFqug1jDvuWMqzLNJH/Lr/41waBzoejVLl06kNdKm+BKs1T7KUmmn/MevwMQYeRCzqPPfdCvdEB
XuCxruDzwA8oZDcVoiQToJwrZUXmLziSb0PPN4S+NMTP8adpL5o142uX4iNjxYRckNmPzfed+rdR
gXkc890/Y7ZUijKzFl3TpgMD1eOMhUNCVhXfsm5Hj+E7djLUzOpL40iOG/+DTvGYl+isAcZpf1YT
bSP7X0U3vAkOy0rOZVXjfdTCHUWRczxnfPqo4CXOcQ9K07qntxBo+W4IqWB8B5WCHpB1Vrzg/xET
IgeI62sQ29wkvPGfoCiFeUfBhT93TafuOqZj0wcdBxYCCU+Gha2oxDxb7M7fjv3Jd12lSLjNztn2
COGYbb/y/1MFpsFDc4PYPzRet+Dn1cd8rM7ng/VBivAFsmtJ42xOigCcCEl28BOeeYcvzVeYLH7j
4OzFSYQPDuvFXBrE5ojQdgsXGm5AaKM9tJYZMT4bfkXp3iol6nBcz3EOVvm+ziDSTZ1nDFCCAKya
W1jBinbAoodC2O9Y6ESC3bvCGb/uJ23ETawjBVBk9bzYhG3zAxu9qrwwsxeMcSjSlZpi1RU6nXKN
k6sbln927AMAleeJjzCwLaYarXFtFSKVoQBcbwLlcJQTPoMdnkKdrIe16Qorg2BwC76Yxj6mNNZB
genTSMgdyMz7cCoeyI1weBGxCJSV3+wEos85jjIJrVY4nLatUTO2dHcovd+I9/So5UBq5eOEtAW/
8cbbb2mBYUF+66ecbtd1i3EufLUEasIcbGEDEUX2T6NNg+kx1aVUIc4tyaPAl4ig/r1jc+hA6cN2
36r2HIY9UW0g6UAc8OyvwnCUHXApaQSgCZUdh7wXi92PUOAfmxqOuVjkRdzfi/Tfm/kyeuuX4e6C
t25WreS88MUKhngAe7Tf1Vfv/d5TzzpyXJ0d2u0itBitv3g0qOfvj8QbbkNpHMPvpLDhlUmM3aa2
AS3/vJ6aJP6IWlPm67XKJNmeZU1WwtS6gAjFhk4/0xqc+Z6kLS6aUEy6145oK++BhWuJS3pxgD91
CV1j/1CezA/hVj7NXzi3I1o8S3C0CJqYM6uI1KDZSHjpYNK4U4m4M/EeY1rcDM4qFh5gMW1rygOv
cNIMG2FSbphVBXthy/BAOicishfG99BjEaF2v2F/wasBzaK/8g2FCrNLvbsBsR37+4UgOO85xMjh
IC0s9xAJGLX9HNXYnjawA5qiwOIk2rZbEONOcIWWUijfro4OfYd83mQE4ZtuM0hu5axBaVxBkltF
tBWr2j3t1z8tTWPWI3dCVcWzU9L1pUeIhCocZD/3PujSxKbl7cvpnct6SeLH1cCtr/OikWTlZeR9
r6ELDrN/qLWXBHCE9aCpkMuQXFxSGRd9nLYMclq4JY/rF8IpSGEZP5AOVhwYv2geZVa6TxFWhYcF
0jO7UruPTwIAQyEFRTGDU/+AW1N1tRPFzOJaJfmQSND7lr00CZA92iao7ziqqyMSbf3P7oJsHpN4
54L53UjH1sHaVDaHUgDm93NqES+jsOin2O93fx5rcldvCZtIlI1/ZDlwXW8UezEfwKMNDBcuU0uJ
yVXcBM5xXShNb38oX85fh/4QhSGSbWHX6l3r5M53BKb+Ov+NP/oCRmXH9qknMyerzpodj9ISPojL
vBaxCWmo4L4k6EuL6LKPGB6Oy2MpK5qDiQyOK+7mVqRXS9UanAi9rz5qjKO2WxZ1b+MFDBTz/LW8
yV1JgwMhUrrqOfqHHO0A+liq96fFBJU5XK0ZS/X+pXXGKJTwLyc/1ZBDvM/ob6UTppjGDvOEof9q
jaWsMK9ZMn66MlGgJFibMr9CojY331DqUO99DsPfvLGgv+6quhvfOeRGAdcJBHDGfkciKIjttpDf
Nw6vhE1f783otpM+vX57SdiLDGlSmBhgt/VSCTEcoPf0K8U/4cUm70bDYchf3RZn+n6NTYqIjekh
VOPNYcYzrQPajETREJ5h8IKJS3OFHeSMMRUizzvBs37gZS6eMc7uM3trBAAzK5XMjfeHTc1CQuTt
VPPgSjfT6+bRbrP79XgwbDSUojROKmBq/nsv1ak0kNVm7F5OYJrOJXRpKVSLA7vJgWrP1bys3M3q
rpUap5n8rXhjA834EeL8wOjRHqJzhJrHQKj1QgMl4xo31Gz60iGQNYLejqxgSeJHv9bCOCh7DIjB
TubhhgaiEADIWbVa+G5JVaUxFtRn7Vqlo0Yt3XNw2hwFWLWVBouuFmCCSPQsHv5w8zqvwwcc6CUw
9TGuSujX/3j+frUFq8lQFRdGHfeFhlKYnA+nQvlJX2NtJk1Y9IvKits6DOsPRaxMd0gy01s23Kto
NTe59Ki956kXwaMXjLj7QykNmtviEseyrq8raIxcCd0O0xfKOnRsg90GtFEQJCzsP5IuH7Lmvjl1
qBvmkc/0rGYjJB20EAqtqz4RontSDZ9yAeiXWDAi3xdd6yCMKXJ5Zxg+soq6Fk26eiU72TdNBHvb
JZXu4u/J/cNDLNRQMJr//rmwVfLwBh96eUdtS39VOZ0LGm3alioehyNiunIOFYcmjZ2VsieKRg7z
n7VhScEfZ1c8XNxUX4X0uWddUR9RFx6b3WGKmAt7x7gwQ0kgCJ9etoIAeRVBL8B/6k+WjuK4Pv53
Jrp1CTSaOtTKl3yJOYEL7bI6+8ehcIaRUXbX++4RG/OeYzMMgSesPmEZKgptuUlOI9jsPPtz9QRb
jojGjM9x0UJoMmxTWB8x+L3/78qo9SDaOdZf7pwhW0ld1twgZ0tevDDtDr+7nmJl3OGr5k09oaVB
YTVf+U/iYnmaX7inaMoH23SgX9i73TEs4w9OSOZJgNbSkBgw4xbBqd8F3QJPL4GhcL8DgzmHBOmC
ShAYysit41LklQBgFbNs/7FsFb5SdAgM5hYA+LtM3wgEGn1p2zCmJSAqEVpKwJOTzek4wxZp5ztk
AnkM3UZmVQ781Eo8/ZBghw4FiuJjD+mdS6jebPelM5ubRJx2KqlgTCMexWdKdbt5g2yFdS1+7Cf5
TnlBnBBKbhviKWq+uWxQJKKmaGGPGeUXJVQHnffvV1ffGNhG66vrrLqRnohw4SpkOoyfu7dM+8zG
c28riA0lvwVB3orgpnzAmsLxna5MEPEk8yqwLBSs3VbymCd5vbWBZcdDMxFBKuB3c4xnKM9K6nXK
Bh6Y4KchuuqLs2GyGn5oyA3guMHH0gFKIKyhx+qowGe4s0Fheh4IBnYD2GaMKMXLqE8CbjD3YOZM
aXs4grA5tmzzof6Vxuf6ydhCKwQ+QxNI1lpSvBcA/CymR9SWj/SRahWqlaYdS4cjEjQdi0wqkY65
ctOR4KFH5eY7gakOhC685mF9omO9XoPywqBAxPmgdE9CMfbsocrF6IarEXLdaQLXO6htDPqkdCrs
WEGtzESy68UBW6wG0l2FcpXH5i+RMM0sHSSg6icvbvJ9LL9a9kgzsAzwTciDLNTu8To9TMH+YoFB
iLhBwDOsoDQB7r8nEuUc0LCnAwqig5Lv2JtGnIp9gdRQJWDSC/j8qNNbXes58dtSJzE+T8uHNAXt
NQ6dJ+1+t+7tXpxwad7Wh+W03N+hWIeOJHs7tvHpay/dw0E05xcw96VIwrKyVC+uvmUA69Jfdu0F
bUB1G13GQzW/AMdAK7iQhF8qTmf60b0pUMGHt5aE71GtNrkXGPgW1JqA4MVm0HJRcUvL/khJPTks
tYca3+G01qeiXpIHBssJmrfL9iTyI5FtUSb9fEPfsby2VyRa31fGgdR5NgTEO1cCnmHrgEOuS4pd
i400rwngIWkSZYJrxVZYvKLehDrdlkMH5gToKtWUEHJExup7fBsk1awZYp1+nF75heSLqp85+zn4
+NPEf8+RwYsWMhK7OdooravAh0fitfCDlnWlm2u0ZtREKb0gTza42fwvc6WoP8DlnRTolx+7Sgzy
3a4OriXv32N+qHjf5P8zaRIzvgRTHBY55JZyobIfUEBEmhrKmgshzpGI4LQp/vh9hyjA4AngjkL0
+iWcXDcK7UEnnCn9Cuv2qZokpfv82H9OHWO/s3AGw+lTnM4q/xIFzoVNOVQSyrCOrln0oXsg0lqy
vN86ZLHdn7WWoTnhj2NS5LpsZ2qVJKKyTN+AXRu0QTdgraELbv40O4HUs0lngGp76JRYWBm8Llkl
WSpXeA+gpAZKpg1eGeB8FysM7KyMTELnbmH/cypnRnYVnyVRGCNaKhaw6RiL9yUJiFvQLfN9lhH8
Z8J0iKiaHvG8LPmSAohdlivQE8BtUPAsGN/sD9Yjs5Z99TL4VQ4xaKzOnB52Gm+rb57sq3xOuZDR
vyv+9mZiF3Td/dIggBU2Y1qYkdx1AgSys83cE8ynD/a1hyofKtYIckX5OgDHsCJpsTjr0r42+Qn+
XV+eGEq5kyIq9r8IzgU1tJJkWGxAj6KSm0kfRpk5IJKz43SbSHQm20qQsNH+LMJ9jg+aN3BZoGwJ
RPHal6S+f5N/Sob4qQ5gAd23zdHPsLTOyglGhFKDcaXdsngRWkLufMm83dd6q18ymG3q3Pm3PHBj
F92WZkzYFA0D8XS35/22H+Wwm4BPipmv71IJEZIqqaX6Nvuy4/251D6rp5Ot6GOt9h85IB+lGYOD
Rfe5f++gGGcI6EQMwa8W5PL5fP56S/5+9dXzJbDIzzDjT0Ay6RKJOVeCQ7xVYyI/HLXqdn9vaXEo
cd4s5Z8HmUu/u4rdSI15fZ0JlVm1z8UzmpSet68z5qoEiBA2M7jafE5eBWkj939i4eO6LhGI5/MW
4igqKZDuWtqI6k159gZFLOqBOAL0m1yZW6c6HhUa8HKgYgEtUFhLvaxNLR7efg9uBgnLbr1vu9Wn
1VyPyM3u6ck73D0ODj8r95JTuGwAqeloDGnscUn7BI2uZ5T8m26U48F/un2Z6mtSnae6t8t8/Ub7
BCMz56hda4CGV0RtZcHhdO0u4czbxB/S3EDOqnZX6fyP4cB11YHzxDbNvvLvo53//Tz74N+3WunE
JfJqhiC1kZJJCKluu2c/3pRyuY1hkV/r23QSK4uKyExglIl6qix1FunpP2skj1UROYd2XIs6sXWq
xwNuGBFV/NY24T33y5HstG64lNor2dk/j3ls37+rht3A/yNkGfv1D7Injik+pP3pLAnI1YblJVmn
SIROvNaV+Er3KDt2Xs80EM6eZHmHQ0+m8oy5vwvCVvx73VeXH0LE8hj73hX3aluOzS/JxUbsNfMW
Y/dOlW8icB83Upl83PfjtaVAf7fwxN9k9R9OQDVKsEFhtJY+Bz/dYFBjxkm4KLZfbDIzp0iDeAwE
8oAE1KTQp6tUk12u3l1jwJSdIJLPjfdWjPjw4+w9fYk1YCGmWKQGhnYUVdVfKv4jb01EM0TEILcH
3J5nEPXbLbcfuhDIjkyBxAcDsFReBdW+0gb631OhAblbtmOzTw43yfmlLEl7+xIhCKF4LzLn6ntm
PHnvAhEHi5mINSyPi8MTdtcZOp3PmUc+GNxXhFuZ+KesRaHEZGKKKcd/nGOJZwwr7zl5HfLGup9z
mLv7ZwWRmJHbgYcHP5hNlXq6uj20tAZHEOJbWDyL+Era2oWNPn6oxVGkI+yPBu41yWKgWIoGgmof
Y0viFfkyctDx6sdJr3kJaqGkBOv3Zyez9NIizffFugByZehsJwkPV0axni8RWD+rJ0Lr/nrYv44B
4BSLYvz9eV3bYlF9fzHYkz59V9WMAmN36qFvQFXfjzQFo3nwWyvBVNwkEkZh78fGQmQdtQA+dP2L
7WgkJeZCMnlypVuk9BG8PoWgDmOuEGcbrjF+Ru64Ywp0fGPu2g52aY4J2vMY+fqEKkS2hijhQT1C
7tgc+EWGhuD4SuxFwjTN3rfbw2fSRpbxgfMbgD7p64vCrATQGdKqYEmyoldAjUmXeNE2/oShudp6
SPFeYD5B4Bt6LyR9mjxwnF/qj9FiqjKjDOc7bJuTLlRULK6g9D1TDC0jaRnZyAmp4Sb66mYrDtC6
gQXx8b/iV9irGsTO8cQP3fcYTfbyEsWHT3mw583zOQGV8uBqjxIySAzjhSzwnU60nUOee3CqygfB
UgPWO9a0g3zb7Q/asKJHZRY7DUsW33FNPHmHBf7dojYA8fGb3QWtqoqA6BTvPfA0UA2qY4H+rn35
N7CEuoT6EjCXIOGz0k2VS7I12JKBZV7F21rgarKxixCn1zYxKy8VS0s/42u53AV/viiUHGhG5Hxn
XWwZMrOGw6D20a7f8aNzeUZrePNP+N3K7kS14HB3cfACKGH5mLiiwslIq1bWGPDFpal+ilwoVxBW
EaHuk+SF5mME2e6x6Jil/1chBH1cmWZZx1Ttp3u7okAcDvhmFqA4oKE+rZrpxA2bBqDCTlFqUd99
BMoYgaU42cJrrjn3HWI7Ov/ptkLBzThfoeCS8F6tH80N0ofhrHk6Aa0TFcz4M26++tLcYgi71zwH
8Dr7QHxA6mqa2MU0PkSPTOAn2VaJ8DyHpULP40xHDiuP2StHRPKPP28F51nXjR1POXGYHmaSZ97O
ha0JB0Bq/x/M0KrbXvL1lX7y16pMbyeszXUwOYHug/43zOaFIOFP7hgpP0Bi9vr5sf1/eCxUbxCf
QU0730ERuwp3LafoLtPn9gamYFa7cn/zJ+ecFkTYhS7+4fCCaPlZxj3lTLAFMUCpnMEm4lRYSOXG
k4NhH+LPtmqdLDEORrh+8kPoom6zufm4wN45wVfrV5X/yOcGakeDX9C3u/iEUsZj3NkO1KAvPDBA
Ckr5zDmz5PtVfL043i15e80hKQIBvlsYaTYCAvevYigK7WcuEuoaFaXJmaZsWGtR1k3fZWC/VHOZ
zsZvhYso2/JokbS/ooJzqlmechVLuodzXZ70ZlaohEZ43UhcWssi2on+NFjMqim3uQqW9J3LoL5T
GGGGgqm9RmMj/Qwe49b0wpaul4Pw8yUeGdMC7mloEFyjstoBdVAch4htuy7ouQIJHVclUYtTtj9m
/uxy2J3+6GGdHPvKF9cpLbZEHO6Htt5x0UJ3by2j+6fHpKvLGZQe3uevCxZ9eH/DtfelGBed8Fch
IRW70QaTIYIkK5BXHfEWvmW4133s3n6zAWbBL8Rw83dqlu1AwQkt7sVNrAaeLhj/DWuyIVirKVs2
G1dFOFlv0ZZNoGDk1oOS+Fw1HFwKacy6Vycl5/J3xo9c4N1RLlRSxsHJpcapvDyQT9a6pgN2GjNE
QnDlPSmGNI4BabwDvW4MiblpoTUpw8BeVSC2vI9KvUvzAEPKIag+aXpylPPw0ybo5mcqXsO/xxY7
DyBky65qF05N86M+zDkyOEAhZf62RHwDaA/9ET3hkFhRM5PF+XfO5TuXJjI2EQWWIdr3emlsYzNC
bQrhMQcblAERwpp71n2FJZxcxUBuB0aadtR81GXsruEkoOtOfSZnf8aF+TYzfDC7ys4nkX4XNfCQ
6Wlmo9TWY8rvRAfX+ywQle3nZ0hDKCzBIxAxELXOGClRDaxQxpV3ch8imGhlT3Z7r7C3tn+cCzRk
eMXEUr0uAkcCQXWgeRd4I8W6Bxbt4PgRwe5eKDEViJeHcAbjsRFEB7zYyWIyViMqtW/WJThAYOJ0
c6NzXfJA8RqoCB1BgYY/32tm/MYwOKvojqAiFv6wZv92JCrlrjvi2ZcM3x62L9EWgZjtzoh6pXNA
X4YGMPcV8A+b9wPj2ElTBNGXdKBndW+gWrZc4yCN++3N2y2xYqxEIyLY6z/1/WoJd7bOl2Qx7R5j
JWentpEZSUXcz8W2VRHnmlVFktzGwie+ZelnkvDD9qyqkz2XHbIDtutqMEgWZpGX0q/+7XvaMf5D
xS8yWoOuyMPfW+I2JL92FrhOJ9GH6wn9N2LA32BgK64sUn8K73NpfUQRqsuklDv/qJPMII6y0cqF
GqAVrG+CpvxZGUbELOj7mZry4LUJqUvPopRnQd82Diso/XOHmfxv2m4WruFWfZSqEeq+Hx4za1Bq
BvZLhFtZpSb18uXLPn54RAmiCj/LEGaYD4yaeGAa9HCFsbhGEZqRP5MBWoiq/ygYxqsgHt7iDFbb
fY9QP5a/bUW4LBnmHCWM1cBWXNXanSN7P8O5KXKTklfJ4hoVsfGgDPlTAzdDx40gT8al2NS51cxM
5WV8M30ehBgGIm72Gp/mQNPzFp7GfvkqM28cnVvp6OXGChmqNeaTBvT9ZXbCbt5IEph12oYBsCh5
fxXgoZpKcXnOKVjNcWSjED25ieCthKnUtOJT2sf9jORrWpSK6y4cKK3FRjbJFQNBbNXb7eBKYZE2
p1KuCt1XsnEYXAniNrB4vUibq8P7gdsIktrqRLakvrZhQNkGKLlNrmxZVvj6tyxTUdjqr0Goxe+t
tdqzdhYCwRO5FkNhguDgeU+OLfx9TRGzFfj8t0QzZRunWPVe3Poqm7O/8HsKsYQJUimWZV6TPG2o
quQAZynaj2F5qx8XMmrm4oEYEUR2YSMQaGnpNRT0g04TZ4JR1huRoSJ6SstGgOTGBbM/S9Il9dPB
Sbuq+/Ma9Q10OSxbhdXAqEYanM4b+zCr1vSVeWCZKLGfJ8nPWPjowPUxKvcVDHt1CZYQnZLQNGJa
JIURQUsLNnZ7pfFk1KMcmO98/HS0hzdOFvqbHCgv6wW+4eOLdavJOGvmllKvNf35emaZ53W/Nq1Q
trQXe4YEJnL6rs7dLWlIA8BhAV6+1sn+OQwTCD5Y+Eew+ivSw4s1LgipQyytKGiUtPB6blGMeZnD
bVum9rlqs/6P+Tx5HlTIYXH/o5PMSb/+czfnIK5w9ePGdgLBxoomWFvLg6XBnK7L6qvqFK/fYoR/
EQoQ9dOTAMfj0wfd686uTM7B6bBXTqyEWEJU7gvOnl3sSbXZnu1Wa5edvn+7hZBlxhb/N2mjbG6o
NCGRqfrr34HaL9e0pfApQYCKWk6lkiyLrj0QKAPiMKqyZ9lvf2Evad3T17JAxnMWJs4jofgIwMMb
sUYnSZ6Ue/0bVztbiylmVVpzX5TlGteJnSixHbzf/Lm7LPzdwfXio3Kyy3bs3cBQy7wHMbmh1dJX
SLjXhZbYTxfrm7QRoj1MXy4w8LvHz3CNv9jHcqMma1hodJsglL8xLGhHQa6OTIcMCMtl63umX/8V
h1UQjqYwcte7u6b9KpCrSyztRKbDwZuAH2HxUM84L1IPAhy2o+oyM25+FWq+DRR1XP2ijIuYigpG
mTaVGyGrobWG2qOAVcmYFFndTqEhyq+ej/mn1dJccoTfZdaMPI6wl2YaCeVx8rp8WXm7XQa98FW+
i1FiOV10sy7NohluhDl9EK72uIn33Vqr2IOmiTAivAhYhCedqZ7pdYhb3DiXLW7xFJLdiYlTk/vy
ayq3MOcw2rczcT4uCRBl7Oyt3fPY7FQpQ0ynkLczIWDqndh9FtnybJ6+2njW6+ZoAyVwYpqvUmeJ
LYhRqS0yaMHFWLNv86JAfFLvRoSAnZ9bX4ZHsTbbeBq35IDeyYDfpkX17EFuk+3/pxfgpd5NHctr
b8iCaz/w6L/MUxMo27iVDV9oNAvcYJtbiQcTL4jPL7aKgkNxVcJ6oKExznWMRUYR+Z99sf6tcXdw
2eWZ0xR9hmX0mObjKI4Tmu9lmHAzlPK6zEbBonhStnftu9Wss6uiTiZM+MCKz5/d0OUpWd0+Fl14
aO3A2PK9GfdGR2s4bphN8hUBHhmgkbPGBPhoVcsYdqn7zVc7MqtSHhH81sN29BRyUIyW8jHOgEX5
hbFlxETRAVk7PB6yNN2YtuOg0+vGicrluzOOoeig4oUslWJIv+pznBswjGTHrHbuoh8VKIi08lwK
KkP4L7XktKfH6NUteJk5cxrZ8VlpC6/ydkIN5u585n+MD4er2C7VvtKNOEEDURw9f4o34pxUA7Yp
YAen+AAxRmYC9emILNf09Uz7vYmJ2kC0xIoEA/+couvM97Sb5l1bfb3uqkCmYyhIzQhR8YVEliH2
vq3SUakZ200EYmxXmMLi56dsWe3CTxPmtqTR9ioLps+E29fBTrUn44SZFrRpBnydPH8D1aV6zUov
dmnNma8saxc8uKelMyVDFFgPjjwahayB8uzyzrnDfimwhf9XKPLpCAdpXp6dEReqZFpA+GrjNwDe
kvPHLdFfQhzZcKnJIpggu2DBmpM1K9c7aSIBXtC3OJtjz2wJzO9h2OaLcMjzD0Ktqf1cr1yAJ0eD
Zrq5cwpkCYqy1ke83p2NuloU/1OoEODrOwV94KlYbXc46nZ+yy51HiUokxrIxbbkkzedyNn3h5Lv
j5j14TcqN6fteBplcLkrDlCCJ7SvCvmDZhdVkXJlzvlbWH7pWMznppOFCfuJh1ZaIFNx8VN/bkwz
GdY6MBRAb467uJ8RK3E+8hgXI5gddVuWxymcwrDAu5fMbYyN3NRfj6A9TU8hYF4ubaingAKbUyGZ
iYyD9UTez0TEEyQOsg/SvHVHLTkzfNva4Q0Q6oYcA3O6ra7/rFuElr7kGVA57SOPEW2DGfi2PhZF
XQsxKB4VhB55MZNO1BQ8nqlVJ+mV4jE5xdGMoMsGd8o7hFXfhcPQZc0GmVOuIWtS5hp3yrBwWXXk
kA/OqL8WNTXOipENVxEOKdqM0sicMjfonoIEAubJFTLcINO8wHgpJ3vezf7yAqIZvOLhBw1KRVb/
erv1/tpCTqP6S6tqlz923F0U5XVm4MJjOynnSyt0Ef52L9iGd84g77ZG0UbQ4NrnNnQmZHM+KRPG
NfZrJRp5kGEZ/Z5ge9MXFgLYqKIDRJUf7HSqJQ6dKlf4b8sGyBcrSesJk1HrwiBU+cMnORbl8B28
KO4qZwYcystqrgGRuqWBcSsBb2AOWOqU2tNj8Eb8GY7mytS3HQ0OvWgJrm4gn/P9V4t4En4mcS+N
+KGr9gzhWjeLPn83++qXF8aoU3Cv8aFbFblYBEGFV5+Y9jEQK5VyrgHdVb9ugzvWYANkSMunYtV+
ZGjkeu+NBGaE1s7EGmZJCqvcoA3loJ8L7lSjdpT7V8CGEc5A57N3s91z48xzsZwoyxNWpzhBXTOE
df74g9q7VNn5TVyitYYumLqp+XFCbO7wpxnmlLRF/9ywDFbGVPqjC6oGmAF8Dtjl2gU/iOqAuREt
1J2iJeijDnvMEYeHZs3iLQzIc0cO0hMWu4OfwhSTgYKGeqgNu/gbWXF/onqHq8icdYQlqrHmIoeG
5iGB7klcYHgYwb6y5IldSvhv3j72qBPRFLbTbX5P7ePC3A/KzRhCXjrXxUHZJZXswiRFnJwkn4pN
siHeVc40n0xjUiHXe7C0FVfH1nbAf2Td+sK8IXiW8rVhpglx8STLJS+/gJ6+AYbPZo1Koc5ZScdw
RxtO6Hjpy+VYFysWFWh1o5nislzOO5wAdTvHW87Ys0moqCoDTViD++bGJDP65Anm1ZheVcabrAJy
N7BlVLBLqSPyZrjH7bs/kzjEs3wLKxHQSeU2vKZMv/Fod+pYdxxmx55DP9cyEdf63JlIW/l1RcB4
su9QJmzv4qs49DVMe1vhgFnwB4DJhdkujLIqlmM2Mp2EF4QJ6x4QehZHDxJ7oLRuzs/qH+z1dmS4
TIusNJS3957G15KjRzCw/rhNtKbb6e3t452zfR/OJjW/HWKLmP4hvZlWaubggievENVEJx8WIABa
Wk1jIvZ69f2S6T+9ZQnBd0uYeJG7Y/QzNVowwxddhPjdmTANazX06K+PCs+/DpElMtVpcvSEOPeH
Da+9Ov4T+w2dMS5d8+a5S4cSKMSPbXb96D1snp4PVt+kB0vv0TGwY6oX7YUisPDxDiXfjoXgJTGK
+pOgo6tH8EnMSSVJX4YuP4Zyma/KZFyPXUCqMzhoeRrR9Gdg+uMrFqj/QN3UxTQRWMF6f+Iv9a0E
fqzSLR4VDgDF4ASlRB+SSRMQPpjnYy2PikuFryHOVk2PgyKXwpDQZz+QHPZ7t8JALr/1U0KcdUoi
U5jcFJ/Nf5fWLqNVgNUqifDlZLPeeCdDNPYFGOFnfXhCqhq4YnW++jfirJZ4hYGYeFkI19S3pOIg
viWDDxt0Aic/mo3qGl1iBxb8LWqwukCpcjYFOi0aJv2m7Xk/9ltbQxnCYgWkmtE+11/ElimP6LfU
TiYZKxn0OpDGMGEng+pr74a8gT3wOGVKJaAAZJgDy9H+viJMpsFb9D0dsbjxi/6Exiw0IYeifyMW
Ieon7opUwHrUEWkPUdVNhIu17xcY0oO5aytvDKIC+SBHk0plDpvHvzqybiENpZ/tnkEgrwnJtUxo
X8/v2e47O8pEGrg/A+rbia9ZXMrlL54CyIELjGXxTUkP91wMuuV3xKuCBBUh99PF6Wr1mLkHTbAl
lpoYGv0EcsfXJTCAMPhOQWHjm7zzk1hUWoHQVf3piZIfX9kPsJ73RBrO8DDqRcdmjI/MW+uOUp4F
cb3SkGQne5oLcA09B1nX02xrSZ/mS4+s5qiDTMyiBjuluX8tpz9xkcIu+AZrtsP0vPlpqyuOifLg
qo932aW3YhAt+FMj+L30z9ZlXkatYk219B2d/CfQzGrUsEQkWRaI3SBWEQjR4ibztzGYULvwc1iq
lka8Oq7geXgd1pYDEUzQhLBqV5eCep4VQnojAabnVTPnKFIO2do8miINWWGvUyIPDgP93Fh5Hlf8
VvyXCys0H2GjLmiyXNU46T82P/MP0yMZw7uKmBX7hAa0YkyfvuiGePXrmvtUr6BZTvbTuY4LwjgL
e19lWHjJPO2w7N1BaJOUtDPvWrDqkKOEcfelAgeYXgUyJN2Rjr0W9Mjjo/0NYGEqiwDIInzRdZfh
xjmYQeFC2J1rQkxuQq9F4wxIICeoduUrIfwq9hRznF3lrM3WaHwDbJieJ+xioGCozBNdkfGVaNHH
EWRROPWLVVR6QHMeTFEB4/IoqQ3fxdyhIjU8ohVnoHmktoSP2OoaoQqEBlnwIzl0XIaL8NAYu9Aq
d44ixfcy5UsEhwgaV3EFF6IDzFbeKFF19T7O5qJX6jUA4J0TwzSP257yVnPcMV3yzJzI4DBrncz3
y7ekXbtqB964lbFoTXDREMagd6vSl6STE1Yo+JeDcuqjWyW2akKGfQ8B/r2MplIu67c25R4PSbSJ
7qJL6O17eJ9U4lhbXF0Umpp8qxUFiNE8oMUtvipa5jKElOfm9hHnWSmr1TcVqFKa+DvxvxrcLzya
/rvS+35mx2NN0+0dFZEkPYDGXgzwo6UPKrwO+608zkm24GJw1AAcxK4ZZX3DjgLD67+XOyMh8BcK
ILg46ajPpLLBh7XNupe6qToUZ+Rv+WNrJ1BcixY9lARHvIXUnNubv6r4yU9FtPGNDTL5bh2Mxyje
RQ7ACYRuLLMW0/2T+9UNh1HDdrWltE2a7CcD/eKimDSz+id8M8f1qspIBeIIPs+x/axPPP8Rr8Mj
C9WaH85s5AS7772CIC2LZOM3y+QxybuISxwlnUXrVhBZ+ji/r2Jj6a3Tp0n7iUMbiVCK/6X1nGEZ
/xCk7TqQaIGr9MU1FKbHGKmt500nzoenZfOIP7ZQawFMa/rNwzngK69qRcbPddkDYB6BDqHXThk2
7iKeu+FCLo3TO+a+N3dhwDlFu00nCbKAyXriqgBZJn32YkAipk2JvAd4lPWSyN9laxIhhbtRKgpF
hpQqaRifS8wwF49WYJejgsxvlXxLvxfH14+qTDZBG+8sxzKZToUa/DtX5pRUT0KoHYU+i0/SKj83
TCny6xuLcdFTk8ggA933/MDwi7p+G/OC6Ht4VG1Jp1f1W2092YDJqaFlbYQSgpCKmtYCJa5f+K9q
gs3ogAWQ8CEW3hDT2ixUVRaw2J61Z694xYZkDzcWi74fIRVqkaBEWOPq8ip3+UHObQICuao4ieeO
+8h/p9BXU5FMrC278aRo0oLWk0jxdsnshZSxDg+GvK0Srun47UafOccWn6fiotZE+7jw1X+AK1Ml
TZpGRC20zuJHYYwc6kGTQtxwwAc5XTsDAdV2wbdco20FHqPbdUdPg4BTPew57E931KDr9RRcZM7a
xkzs6DbcuqqvUQry2fLPNSuBvp83bwgI04SJxik5iJ85OPkZTUQAf4FZk7JKC3IfoitpQ0HHFviY
VaHH5VGEQpNs+yvsUvXMtubZ9roW942h4rhX7cTyhh+6E+lalZNo6k9nDFr4zUIvXuhPRFBRhBL/
CG1eMgl8nIN/ZD70IC2Hm9uF+1H/aKTejNvlkd6DXdsKU1y2VNRANZ7YL2LcUv1/1l2II9Lr9MfC
2GsFOPAYdybgwNyeYBEACDY3W528cmUD+eOeASyk2L8sGvdyOkvdaIeMPbbNdq420GciEsqmqMNX
PGwr94ilLViwMniywiLYsEXdlaMOEepIKrCjCoWCVThNagJ7CNVUBASrzVm0/HmhE5hmVR66Cw1S
zSx9jsD0IsfoBqDYucgSnAmMtwcUsJqvJCVPyHA5P9LY7RmR+AsC0uvzPmG6dJbr2GE+p58ZJrpS
95IdJqkMtsKGlDI1mB6vTOHlWXh37KHTcFqmb+ELw0LSN0Bcu2Xlospd3yksrKIzsoDUF0H8SiD6
gRFgyZDP6XqkGg7QktVnsfBjpSsWSdkBaNfdx9p8I6E101bbKaaudb+HZRIR4mTNYNZPvCJ4bLKe
UyI+7+g7W9oKMWbFZi6wEnvv1Bdk+weewCVZ3mK/GKPmfT06W5Cgl9Qvq+4fOLvZbZaCrg49ouDj
pGamLMwqlKm9HjEQuJ7DZY4/TjE9rBubn37rFNRv/JKYa2yVv55G7RG2rAXNnEFl+BRI7C4CP82g
Fqq37LEVOhuJIyoJQpizcT6PYoUbhQvNr/aaMttkXyvHFxm9QJFI2jFK5mtlzjtg5AqIDRLtEutW
EA8k3G64BHTuJI/yVC/WeJD6o4TkPYSDygAXO5ETgmeo2YUvutxSigHKp8JHP5drJk/UKjhrE5HC
4Krj2XCmdKlwPvHqcngDBdZXJdXKHGkdjwB3sOlAAZBp4/ha6T5VXF6UsEuYquuGsFEEPS2k3IdL
+V8a0KmE+r1OwTTtbaNJB3ZMk+owAXRuvcg3zNOAmkAT1KEcRTIq6CJEPyEAaIU2Db8ktiEHjzTZ
ttTGRNhSiknyFUL7FVnp8WCvDJgUeRXLV8kmQj8VDYOD1b0+YhArwXrpc6i94n/kqxnkzWaw48R1
TrEaf80lrKmOAB69C4a6rwyIil5EkvvpP/0G8vM86ur9a+W9Ef2Ou9Vhu75m3ej3rMPlAusMTXYs
UL83hzdbnpnkkF3AJiQ2/xVMkfM7fRd4yAogTwriUCD1SOp5X+lNHn8xK3A9Y0BLBrU0l5JGpSVQ
Id37n1VFJJS8ZW380ia0OXVxwmqjgetUhFSM/JU28jQJ1GkR7z9NUnAtepuJBVCwbC+2kWjMk8v/
U+TW78IJywB1k6H5Z9kmcMakraL4c6QTT1M1Ab4ecQTPbA5eCrotKmdb9Xd6j6nRo/x2DQXwTy/f
+n4uDlz9WeRHtY8RSLUim2doyidMIVCb2hSIKq5XMf4XjJANRDd1wwLxtrn+rkbjiiAcC3Tirk2V
hNdkMjj5j5AHv/7fN6JZlkvT6dKehpaPpttjsi65xvQNY1rMU56vwSIojfzLsE8O1JeN4GLDrlnF
+r/JgXqD9sOckww52CAtbmCb5eXkTNxiEE7Q9xl1os3i1t/KWFgXFqUqKOJJo4jrcl0CZNjgNCNl
7VtZm4AA9fZGzIi1Vy+5v6ksUNQn/nDaLhhaVmudKIp3y5H9ZvuTK1GDSVn/mdAULKvkHBFvfWyz
xXkgle+OpjEzFrISCdG83B0mnFRxJb84e2TUL/ROmIMitHpbqaA3oE18Qgu1ZbiB9KR+HeBgTTqF
f7ZCuw6akP6lJtGWRLobWEa96M6Eu0oUBJ46zAX6n/nb0OYf2njaJp0N08rqW7ceIZLZ8tv0rEsN
M1NR0iRvmllsi9rYx0V4eG7rrlRD3r2yVh8D98c3PSUEMmeolXY9BmuwCu6yZsrsKLaqqVCo78/4
u8OIKmfnV/zUQnILr8cuhwDbn+pV/TT/BoTjPsWytfHVEKmMnfky3rnGz5MvhA3qEEMNd+VXRtPe
I9YPyNzHnjyrbFSU5suKFhnOoCVFm9n0OYbPzptpVKzLO/CFE54zJCBAlmE2qPq/1nmpTZLWE0Lz
U1HaCfwSD4kDTFZanA0Clq8XAxbt7jwqn46qYiOxewAxPpNOJzNW12XkXRKS6H+ln5kVqvvDSbWF
BGaGjEkijjFxOhiCE2YKDvoKvrIZ1v0OwJXiqy1UKb0TZ1GcbhQ0vtdcP1vH7OqWtQSUmkJ/beHz
xYsshzgzle4QQt4hRPPBOtuXl5g1fWr7Tx1G8c31DCNhVywnsjRV+P1HIor5+ZXlyXJ5Dwgw5Fyu
qoqPGqTwJWoU/m7+uHMjtlTY6H1+eRcYcpv6BS6NYmClzMrIRXqXCxWLgtsKEzZcx5VzHDna7KwY
qg0u/IJtDEaPuJHPKty8WsCD350Rl+/It7MuAECHbxgKN4/uO7T8xplhtPnLSA566X7/KfcitLSU
RGJ7+5nb8UWm67SkFq8in0YN4LWs8y/rr1Q2KbOlcSq2Qpzmf86pN0GTkBpy4AxNW3ubLtvxcnfg
/z0j3tXDDoRf9nYnjHm7Xec45L15nyFWA+60YLTcC5FVnPTiUW8x6y4IIfqyvt7KwmgyOwt9s4MY
LAueLs7qHFTYqsX+R/W+2AObEnerBsbxy2jTyCl3yDN9VQwohCV7l5hRg74u5yxMIZpexAiczmtc
9T379YMNvtKXmDcVt+A093/CUCC6Gv/RLYsrcP2ypdN0QPYkKVkHQI2lJlhYC2bPy0V8u7AnDYVa
GePPDDIbD4rUiWJuDBf2nT0N/mfDLcRNJ9Y9l8nugIZzhDRwqGjzuLTluh0ZstfIT6y50ZFU4Bhu
zsma8qFxOEwmQq8FHJGv9LN+gHPgs4Fs/IZIwiOM66xQLhBBQKpO27FgxoCUPTtuoqVMd9ZiOcdn
KP4Bu5Ubze9fnRMf/34T6Vb4CBNhzXMv9/YsFcHqV923i2r2UFDQAroVehDLWCkniJyTQCoBVS1C
lVaADfLv/bslg8McS3kXjamIkg8ICvAyPuz3vHD++pzXGJFwksfh9OyTAjXUScUapAhBtVZsG8cM
Ng3J1OIhB5VvOV3EtmfGdOE6FoBLz77o7QLAkX5G6MFBjqXo7e9ZPt8YyztR3mELLB5i8/As6PpG
1gOgs+QJ4OPfelWw06G03oMnbu23oQb1f7iHHwC67OOrFJY3ixYss5+LuZiK892WQSkuUggHnRjh
f7xxltT7yTQUb1jmfXs9q5MjZm7rmuVUidEi4yK1QuBgt1f4lxnP7RMgkF7go6CbGhAanOw3GwNP
mQlgsDbyS/BwvcAdexDGJS6p6ykLbQhfRyrtf1ozAcUjSqtDTomKaWy7rQFGFFrzTue17j8WG4CA
B3BcDjZSGq9m+EZxlw8hqGX9HA//qlsM5vqbTQrdbD3/5Ynliz72TdwHbAaXUL8m3J/5mRX05nVV
mUJVqCjnTjHrnNca5ecvJigl1JN7/aHx1JEWdBwvrNRx7fLUIxY0k2UyHgyep9RyEJIr69rIJCNp
HBvz3t8baqg6uca2cnFJNq+ZxTD70EQYNQwOelXYYijEgl6dm5BnkGOueaATB+eOe9jXOKAxiCr+
D3esxVt0/bkpZvdXPS23YpNwCdAfiiibdgFtSpgy5MOiM4ocmyNU2yyGlWePRtHsNwQdP2bkzII5
t0Inteyre2iUkM83T+qwK+w0fTI1vpMfdwgxthn7u9XmKswtZU74mG/wLzO5gdazt6SQmUETW3LP
Q9OxSdSXnR2asZHhiWTljHbqFSvZBhUpbOtEXr/pT7RiWamWp+4IDtagE7MDGYg1aHpCpcNCXC1G
ladLXiqwEpR53u7zag7IDs/duytZcMpFaYti/cLcO0H3DnSyj1/C7c/ruddQWi6iGM1wxRLF2DXf
Y9NEmagjeQALqHPseJfQHgmQd/dbayNrZd+1ZcjVGUizGjgxXtkniZP8PONfmJQ36ojjx8DB5IVw
RAqpAAruq96wrOWdshCqkh9GUG/M3dL8prfoNur6JFwf1Wg2hVulOIc4A+8Tr+jBac907hc3YP5T
MGgo+HgMIFTz8aWzemznTrKV0dfYhTT9e6y3PuzbSz02ytHNRCb8wyokt+u+mRXNxKQVQDnp5VPX
4Zzub6Z8rhI/r+g/Lis5KuiA46TId6wt3EnhKZtrQA0EQil7M73Cek4iAX0A1rpETpSI2XZ/wxI8
MEwmkJeNi965ekWZf+5bwt1VjSSCxrQ31CaR5HkMsdAem6R61YWwK+84/EdPgay4BqDR/4MO+jMO
Gm5Uibp6J03yl6djWw0QChQn3VQtdvOoZMQhjrAqnE5DuODqI0qdJ9W1QGIsFStdyLoChkDhjK6M
jtah1+1h0Bjw+us2IZEy/WYFYACOyEBojaVHct+aIsn6MLn3VgX7gIPXxukYaDR4inIPyTw06PQn
tpz2rVZYJTtUvvV0ar1UfH5A+OSZw5WxBa8yH/4EL9gVs+Jf9Bx2SUMKGPDyiOGTRLm6bu/kN+FK
alK0qBbh23NiKQ5P2IUtuS3Dmwf0rF2oYYJboEOU5gJqPZE3Sgvskahkp/tD8a0Vs88AqO9rG98T
B4xrLr/oHmsPhuBvEc2JeOLcLzcdIh+PRg1fqJZjBnzmgvVyCgmXz41ldIRJjMO4mmLZZMS0PQ4u
qgDHrBOoPYDDomciAeaJk3ukbTCJjqDGkiH/u4UfvVgE5r+Rs0CJyQ+di0HqXRTtXk73LlSVSfwK
Khu6nBj5MS9TCPKcfDfiiHnJctO1Us4MLZfCmx6iRqJYdqFuaS1zkcZny9ljR+uTa0XQ1kOfcE5M
jPbc8MpOXar+bJiAX1ewd9EkspKQoFsmn5Zg2ygMz9mfbBevyt3kdaByJMI39KM4uXDnsDO1CvSO
ZTrwnsjpMrRpttbSyzagBU/OPLqp8uhSURyntbs/l6KzLTVU6tsv+Ep/SJaYQ1jSimjKVCMZdC+P
Uh2NI95Jnh63Y4D5ATB5pdWU2zTThdU89HH6TETwgxCLAQKVCx2gHV+KKSPS0L/wDpXvjcwGYZ99
+MPlxt+5YSY9Zu7kzI7516t4SJvu36XV5YQTrw6fjytLetM/kEel6RlOegl5qefsqMSnzpmrZZUo
o1iuhIi6C/U8G2MnJm+7+ZRe8DXXHaDpIgc6JBd7wei1GZqPmbUmq1sJyhmhyaSPUYWOgfcVFiQa
xDGIy/DttcC+W/Hk+z9qAbcyak7ZeepOpCIDlMTcfDaw8qPS3KM8RUdnbxD5nY9PC/0HRi9hAo+r
OL5l2srk0FTY33EzvDAxCvK9P0XjHljC/uPtNTxxVzpyMJU9Rl4IcLXfvhsFoDE1sENH7+Kp+LQR
D+AsH++6Baw2BHyG4/Vgf7/vOR0lJpWbZnNUoiFHZTVpjuPtzZTbC+lczeuqa8VAX04fl+ILqLsW
BiYzLvzLD0R6rxdWWDsM/vaPY3gjbq/LH/Z84wg/sZOh1HxT2R1TDRm/Qv5Rng9RZSidY+NWYLhb
tKZk0WrcMkNx9cf3r9u3RTe4otNbo9FUiSDhZWm4g64BoytJln2rnytltVgvjywrGqxC4O6Ki6Hm
NnKuMrH2SyoFg81VB+X2bi5GqFV3oso05tMYu74VcfSxucsrMNtAQ24ybjqb4j9IPdXb7Sd5XFnL
lrQ/MwJCyMigTtPx5tI/FwOlDaU/oUYsQlIzrh7gQvaAsYKns9USe7tcWBhkyA+7gVOx2Ky/CezH
eZ9ZY0utGWyW3t6kqYQFa36JVyoWNcEQn4R1cUkresddUrIsa1ud2sDyy2/bFPqPnOe3T0HR/ll+
jJedrCtqOvE6zJCefPE2zI5lurcTG5hdH0Dz0FcUjFZPcZM1B2BzbMiKugNhwMJw9GvTd7CS0vGZ
BnDoiB0bjsiM/KkI3lJx8DJaLLhWerCstWDgxlPzU3spDQDyr4CkExGG4ybhlBc1meAt38C9rjsT
gNP5jjLaC7Psblcz/Xr66RkwGeNLle7LrGX8Npt1FHBZUNAPrCSXKAO5OkeNe4lYnesO+2gMwtSu
mz8GcRKq6J/2DH4erAIBTHMbYNgCUqHLY9zN1+C0a/55lwDLO6hyEQdg71nfRnwkbGVNcWrCdrFp
4QXe34zLrGhJrPbv4OcyFwAptu8FwoW03L+C3c5HoMi2eSIkiUzfZn8RwaxSZQ0VMPzzD8mMjrsl
EkQcCdcSV7/nXqnFufznoMLBe5ZDDA0rbLvZA2IW47FqdLn77sN46lRqLimUZwBDIoRfFpZMGh6o
q+nLz+OEs0IXv77Xo9cbFc2Cy99D0EG2qO6TF4DbnnQuW/tRppSzNWvDvu2kO403JKAIHrzlqecg
Xjvv/UbTFJ/CkgHEO77tf1g77N8ZRAewm795WA+huZYT+LW3qXxVNINkIyKK2bQrX/oD+bkegkOq
gpwlJRS9YGJtxfdiqC6Do8FBBu0wmNIvYrNz7qJAnTYYaVu2ODIP8ybORNcsWNvAJQyyf0487x2C
BHkS5uhelC8F/vnFEcnLsaZt2iE4RygHH8s1TbT5mLhEVy7OBPChxZEa6EPQTKhAiVgpQYUCBqKv
y6OMc30dp8f1MUY7dFLjzj/bGDOvIBzLHVtRwdXoZiDuvEFEwu8o+UEiPyDZ/uQHfki0M31V8ASr
tNRySfabxtHyRnvFnqUNh3S5ZTpgT6mEdQLysB0dbSM3Wf4IGB/kCDcjTUpJ1h2ERVL+3KIs+aZz
RFRdK8x/73nNxGiK6Y+ho+BKUXQDnoz6+ip6IaXGWUPoakFkualUDMbnnzlJuHxCeezN+bZZnEqg
aimAtrFF7pmWXkcexDOX7/cr9bTXMzyhkR2tWLJkPcJpYhLUHa1VATXbFrj6oTY34cf6lNttOCHq
f01tRmIfDHc/ld0ccqrJmz32ckZOCe2VOWNoDgfeKn4yvAiLgZlTaAxAzmMNJ6BBFXDThFDk2DO8
fKfcjZhFU8GwBbdUdhqygLMBEtmF24b1RFQchnOz/B2XaELroJaSqlaxHOPNM/X7EURyEtACtAaA
4/W9ybluKJ4xXsMAnNfBb2/ZTSMVkKKM83V76J57mqBwE2mygZfaVOXRw/1Iq796itDlvt5i/sxM
21q3yRYs5IFOeUhAWehm7vD+A4Ecn3aLIOcUHp03PW5egDvuqdurXswNgtMld0/CBgrNVEE7ubr7
s/Wn4SeXmeDnkDX8HZgN0xN1JxX0WWdBZBZqD/hc7NrrogsF9Lr24JiMJlG/AvahzrvrRY+b2mSq
PdbSrtJiv0lk/jcig71ScSCpJAoXsH2QgJJuiG5wC8ZvbfpVSqVqT3j0qPFArc2gqo2XpVnps8lr
Olqn39Perfkgp4zTodV3LViajFPLpcQRtEPVO9JJd+ykHTbS4dcwUL3DgGbHcR4waMYewXVA2sVZ
xQfjjRsVQpDGZewDtvKZ+3A2LrUS/izSpVDtHyWVkDtDeKADvEk3IeLnaFlWgUCQ3fc2GGQKY2wi
RFP1wzwqhwoi2Qa3j6l7oLk7/ZfsXghTmCtq5istgP1s7ON6Te2Rg0dTqT5evNyDvQeoMOOIAImR
C2t6SZTjOnE1i2PSjW5M0jfRBRUswTqe+4DwPIx7Qfnf+mvvjvGabL3V+/YBh4FbnmNC9LQAtkxk
fZW+Pdv/z/4kbcNkVY7YFRTpuLABUaxjb9HtgabYEcZdcWL6ABf56cfrtl+4r+VBOdz3E0LRYTdX
hCmsTycghmjMyIB14egjVpBykCfti3laUNmFHmqtKRUKcHIgwu63DuAtm3bq23xZm+sjXGCcti5S
Zx/vsQd5N7PbwwvWeQGzYAIVl5Tqlz1OF+xrZvDRZgtgcT+84ZakeNuGgtv71MUKuCly9P0+OgGG
0RnFzeE5n5FuY5B9RVZ/yzY6SqymTdwI2/yI0RjdkLSINDEWg32gkqnHkPqnfMIIacRcWyH36H83
QSmF5aBGq3dkt0Dy38vMiUnAw4+R+tkdvOWhmmqNnh+O1BkWM9YhIAW8Upt4IcwKTOFozk4mqoqd
/GKQVvX73sTbg3NuGi4hFNoIQZQ4evyhswHIFR29Dja5b8TJfoFaesvsfZS8FeuBSbK9Y4CqCbH+
G7w4RAU6VtuWORssVQ2r6zCN5W8g3hwX/8gadONSkQNNfslfJD1kK8mJhQgcb7IX728aD5fA3Q29
v2FGSuji0bTsJLnKU90RpQ5k0y3+tvb6SKLXOmUe/4Dv09CCDhGsv24UFtYHvifwez/eDhjNxJOI
aqAbS4VOkKbEuLY6aSW8TWpGJ/ku+deflX6RdKMIkemPA7xglQ1Jey7vbqUb6PJulkcVToGxuAzp
3yZ4ZF9jUF2AQ8AnCl19gVWE7mPBiRze/zUxXfolGUPyug2eQA+WzbSTT1BD7ldf3g6mUhKG6Z8h
V4jAqy18RR1n5U6ogX7E/vh3aVthsQIwlUYw1/m8sS8CmvzpC0vM+3/OGZTGR67QQDmHb5a9HQoe
EZVGV2jUo/O4HzfTRZ6sTeJMXQ45gwMH5HsTpV0SSquHQO9PyemRkhOwKqnYayFME6CYDWlzBnkC
nH3TVtpnUkrDW+RzhlH7uHUxLtM8Mpba3BUV0eTXDmJwPtlmodG98I4Ec6A+RdvbnmpRnytThZ1H
xQTvMaGPOfRGd1+lUgh87Foy/qAFzpRgVNFxKZR0/vEtMFie2WlK7HPUz71rZ8/AfcIUvP6PCkrE
Pr1LptlH997TnFuKsWOlMhVMc6pts305g9ZNwOEJ8VAevwwqTLyHCijUvljFjjMPk6YFIqiKMYiW
1TNEgxxRCLeVuGeDaBM2+9uufNeoUBqodMffvBcnTIC7/jhJocCzVLiLDH2YWPELE/xABMvdXYdG
X5atMTF/fTj0Q0OEzZIuapKx4uE/vBuEy1ryUp1izzsPpJZ35OonIJrmafKggNKA37/5H10a4vOI
qWVNgEC+8R/8L/eZDh8b/2NpNxccJH62cqQkZ1pMaBLRaiqJ5eRQdPbjZxOb7tqUuGFVKpu0t/fq
/EDuvlK9unMHYb9Ezjh8apAwQWKXoRBd1HVYEHxSrJI/TCNenqiFNZjEaJLextmOoYxAcB9o4Qet
WRVT2twjMrhm3/IDOfBF+ACxWMj3ByS8TwapjT+613POoHShuRdlBWmP7SStrh/VYJm4zZYrRSFm
2x0uEbHE0md0TvvHxvYJzqQ+otxh069PHqPSdT5lx7k6NVUKAa7Hdy43kEFfsxKRoOOh06cDoyar
Ip5wovrsixNqRhpc8y1UvcUhgfwkJ0oQ0l64OTeKijX87rmb+OVvpZuWeEc0muKYkvlG9jNyFHwk
Bb9Dxf+XVtQ4ithni+zeM0nvfVEMN4w23SKMswZvpS6kU5Kh2o+T26oMIyUoOkruKqElwMW67xKP
sO7asrJSiIeb2/FfdV7pdma2lBDA5IZv839RO5VkF63eZ4mZ4EsIcY3XxCg4HM2VCnhC3Pt0icLg
AwqhBubxbLybx4HVc5auU+aN3/3tkplJpyK5CgHtTK6Dv3Ca+kWwoXG6h76deDu6MuNfv9vOLzOg
WXfE3HftWjCsB4bqOaMqOsdXyHmyWgMhLN9nvThU3aHfGAvLuMr0PL5wcbCSiZa2UtEP+ivqA2ES
27NBylAwjSu/iNV/AwoEAyZnyW8bYuNLAlXyBBLGJYoU3jdbDRQOMBoVwokXcUzZm/s4sqcydKVx
dPEdvjCF2tNrYjYilbjZAx0XxiNPLlIomnmsn/hbF9W4KcD7/TZjmYKdojNAIY0loUvDCkymUYm7
v9eYRZEqGAswLU3hfJv5rj42rXpArFKY/fBVrorC+a8hHValH+mx1nDB7S5KCO5e+lcI3a72f5lH
9+HmjHiv2IAeufZqK2Pe6XwjlzaXtCsq86aCEIOtBD6uUV7DbsryQAn7YTNv1q33vfp4X9268yRf
6yV0riJb2M6OKBHwolFKLLDuyVlIZ8iKfFfHOhWBFkFHO+/s8+ALaY1rD4Eo5EyHUFtS2/fPO9Qm
jpiKcnQ0DiIJbPVqVHbDBSsiLJBkxYd55gyE0eLRSbyD/MIImGeauOKi2mdBTTGergpGQZm7X4Ej
K1UW72Hi0BCNRHQ8EYavwnXPhaS1ftI0O66omckwUDspF5kQUGJTAAUdPPvRwx0pQCwKxw6L64KK
j2iHjAeAFElAvZzzR9ijc2jD7kz2F5HbKluBETunSVyMbKIiKUgRcBBnFD47Hzye9UFl2AhGQ618
6IQrOiWtBZEnOIZwOI9TzWMbwctjqWJZBf0R+YeF6xTsMtfqz4cBP/GqEsjKKkpodrCrRZyPr8QL
bhNS9ra21Sa9ODStwFlqPu1L8VZW7vHtUm1R7U/tsbh1uCdLJcaeeMg0fXNSfU5+wjWNQawd2WLR
xY0Z1N85G0cNFk5uL3DO7ehbKm+G5AjOeE5BEDyWk3Ezs8ieXQRcmdMp8bV1o8cBNndVfSGXq8IC
zXKWnnxKtlIN83fZI5LPyIBEVEWCECCNRgX0daxyMY76v1Tr3/OidGPQ1P5Rl6T2nK1ZSZ8sD2c4
fhjGFUI0WTT19hYX4Hh6ZOBX8hgJ90kkGJ8ofeg0UUyeqCz3chkdJbTtetmVCVNWN4FGav1AFC0U
YzPjqQTdjKB9m6Kn8YKjzvTFXAVEqolnLyYKT2oe7iSrelnwFecMTy1hihImMMKAJzhquV//wYof
E6O4hDLfB00guE7SWaZwQMPDue+jQRWPuHuw8s9wKb3eX9H1MfFXyVXN0TaXvAAuOYndPHVBLrUs
rZc9VJ/Nsk3K4sEhEnjQGH2OB3FMtlNHvUgg7idltpuRpvMb0itsp0+76uKHFCY5AG6jtNaPY5sa
XnAkvaFa925XdIJIGWz88lQDi+5lvRWrJlHSqr5qXQa9xz9L8+tu5PYcf2zEjJxPrv7BfXoWcVyT
Q27b/y2KOms4fD4T/WfFcehzeGSngRHeU+HVvylBUe8ENPqUg9ToIY7DA10t/bppKxfqDbMIJ01t
7rHIbfRklCCx7cfMSnpPDR4mN4LP+Wp7hBKzBumjtXVejjiUo/+qbTv4KGNog/MhL/kff4WGtgb1
Po9EIhUy+3z12mAuZ3YyZcSX6d46gpEyTWW9ntVYnf09lKRVz8xjf0gziKXaUP5sGeRg98hj7KJp
mAzzJJrwX3nc+m0glUyVA+BL6Edj/76TW+JS4i2QaVj8H5756yPsofHot+GHz5GCiJ44DRj02gPp
0JKfYicwgqaVFX4L+uGuSKOkRCX+hjcLMTVt9t0Jf++UQyvUGFTuwcSeNEAiAXdxVx1wYSh0Lr7R
rNhBCiMZtn82qVB2zTdQXLM+Z3PKMvDBsaedkEEMs/iT4lU0T0G+KlYLARPS3QPj/rVi+gRSuAzp
/R3XM0IepzAOmqV9ZS9dz7XtzZSaT3bbTnwCf2X7zPboFr00KDD/IfOBO38TRsFYh/bGWH40xUAj
w4txs+oEQKCdSX65lzX7cP35HLwgkzzpct9THnN5xsJBQaFFSQ5ixvPGtDGXrGayjmsLpR1czdvL
bl3JsovHM87miLOezrngWLY+0JJ1MUZhdLq7WEonUoIfyQNWWGZXeVUnXu/WE8u8ifoiPZ9xuW2R
W8lPe1ORMtj6xao6T31/efYwCWZiGL9c2mROQ1uUd1qv3xHtmfAd6t134H4vTxxF9tJDVgFZrbiT
fNf+AYGv1h0UlQInqD5b9Zc2zCurDCMU8RsQy6jPY2vmNmCv0qgyrPFQIJsLB/puedbSzRWUhJpf
fLLNS4Kr3q0ZDT2OJsWj0O615ihIs/gV5qIfjfsavlGgvcQ4FNz9hXXffgLwsCYpT2Pv9CIr1LJI
eHbsDjt2TdRz5rJPYM9Ijdnq/ymrTa+OEoFNmBTxKX1OXM7nguAZ6xc50dxJFiXoveLbBpO7j1wH
NkS23j4CfCQsC0GSSvWYaBzcGYgfvv52VAdfy+2EmI0eZOJXepwtXIFQcIYw41HJ554tUwFs1HZ0
2fOR9AUcZsP/ZCW85Ex0MHr1t+0N5shQrZ99+xLyEo9wof//d/rBcQNB/lFpm/w4z8Oks0PjLF6m
hcQhIdB/Yo2xhR4KVJ7ubZhKkJOs4dhGbnUZx0KVOk3lXg5bWsVcDsRvpGf0RAZAIYh5pmlfTSnO
vqcg9u6vmOS6v+cOa3LDPvUgE6/qkgeGGy07vPzlpH9cV0qSSgRfkqkdcfaRfjp8x94BEZsaHkqj
BnvxsbuADODLMJFsdqS8r1vCrS+p7z42MNqnQpfaZAWab2hWaGuZjNvDafM5j1pQl7M0A5wM8r4C
v4SdEhbgRHukpp1RoipJc/KlP0UoNzPb/HCA3ayS+74GqjFBnbtK+FYW5v6o8OAcqPUUv/rFNs63
VifjPDxzERTM5Wna6bInp/o5NJiRugLboszolWKBxBt1cL3v91MAi+doAnowfnwUvujQVSAKftCt
mKL9MiR7QFnKhEYPOYtQTmUveQ9mBH3zymEiFk5oOwsPXsfwzS1/X9U2KrBOq4VP2YTr5dVs0TbF
0dS7+zN4YoP/hYOxctT5wr14wpZNmBLpznicUc3x1zHlegl2YSSwpTe1Rbrcq6Al1+1pYkAxCoxY
4KZdMtQTCzhQvIVVJkEGTgj8YzGjr+mEDhU11g19+Gm1+TIoBFPw5AuGwnooi8b7/t5+T1ZLvhTR
FfZIscVwpBf0tO+l2/v9KWQa8QgtCgTiivxv5CtOo+6sp5PrpI8TOdwK0FvzfE8JlKdHpzxrf+q5
Mgn6frQF6lB4CO09GbXJA6K8A89XGEH5kcRTCab58tkH3sO/BdkjDKNZy7o3l3wTfpKsmH2yWnev
aEZtMngxzKkj8CyVDMC2t6ToWp8aplTKGLBenkHUFjJ8l1c9IND5u//iE62x3dX6EdGsvLF29jS9
l8FmXLWMSJ5a8f4mgvCzS94cHlBwXb9IuAsuzOmcSqLik03+nm/etRRM3DhbHInPkNlehRvwcCkj
ZCNtAE+VSNXv8gy0QQql5JO8suy5GN48ZDkECzu6Bx3YH2JvUUNVFzagb6IdZN6TkEwb0gV8SU5J
jSaSWsT4Fh/yifPvKy+nI8idzvyS842r1DSv1Ge3Gdp77wGuaPsT2eTn8Pvv2gerHqbl5+sg52OG
sv41ysW2IC5U97LnA+qx452//XnWpmdybBkU55e9M4mclLm+2pp+7mI6vQF4jmHwGqZYhHGzCae/
XWLAnD++v82jQl48rcrx57Kh8ZPfkubq4TEyNiiplT2zmQQ8gX2yOpsLVcc1BxzKC0rKhS6y+TqI
WRe7R2NnrLLvuvxQUacFddZmZbZA7rbuvykeuCNTgnpm3Jw1bmjBIjTzv8RqDk+Yqb2NYGGIH4ps
1xjpPCh7/ahxjhEyZuERvq9TkuabE6oasE+RhsKnoxRUEYmGlMiAamwXnvhgmgKc2XYm9hx7Bsp6
nvunmuwGULZ7DD6uebrWUuPmjTrw3K09tpi4v2oScV2Ojvp2nws2R+F4KeM3czIYCeHK0QgqiDap
xsIj7fAuVrhEbKxTdjfga1YwVgkPjQq6+j7EhP3PowLItNuzY9HtqMt96JnVitP97flVHgI8fqI2
TKYMvqUjCNNkFkAM4r1aJpznEzBNCygiMhs27wMTXrrU62BacxLENeus/DkSsVzyjEeU9h1EgGDB
lipwyXsir+omExoxmpRGA8HS/ubRM9IoGBA+BNlRYmu/ujsYsAaj7JHvkyjMWvRoUBonDt4eCvJR
6ESvBADI5b6fsWlywmQLj7ePPu27nYgMGBSGT8lpr0eAcBx/nVtxT1YOEHD7JDOYwwl+3yHewrXa
xlUWEXNAUAlNOl7X2Fl+LW3HXT9cablY1mwpabT1znWGKniVNlskpkWDsRonLSv6YoUcgca0hWh2
1I1W+1/1vnhyGXqyDp01u3McBc4sQ4VCrhbdK3TWaCLqmHNU+Gn/Sz4A2xbODQ+LEjzYdiP3FiNF
fjPDw7rcwhAvvqTbmNrB0MUwJNWm0ioW2/Re/13Fz4sH8KH5q6Dh84yE6HbWKrD+q0yUN/gtyapi
BIfn88jMPE+i1/fD5TSzlXJx9wUYKHl6WTeb5jxVDHn/zQ3jBD/jll3JOncV4aA6wb5QpkmUK/Rr
1nL1nD/9wiQQZLp5EJTyN8iANvHMJh/jwuvNgmd5fnRPx70yH3KPfPtFt7zWbcQ5jhwg6g3LypJ3
8RfEoZ/xFB9FXomuTMdy8iZcQqu7UunemWVg2V580A0VJitF/0NVz5eeKLSaBuU6uSWydaI7988M
VyXb2/5UXquVwTgd/cdDxyj99ErUyVgyM3CDS5cHP2ltjDCnKeqjc1N8VLK3xK5Dvd0OVvI9yOgi
34R7SLj/MbgjSgkMyrYiPsFXgKKuIHqWuV7nwbNSntOWqUQho76C9GAjrLNlFjbhTDkT/mdVoUHT
TAWzCWxkyuUfHPYcOIuIimE5NG27gDNKOAzqSQSOe+uxCSS1GiNXXdpQNqxZJss0s6ntJna0f/yO
iAseHM0n/ZWQXtaOyrb+rtuDmGGP++zAjP1SBTdCabtxrZiTr2KOHR8UM5wEz+SeCHU1OXz+2h3e
KT4mVWiVici4mHFUEJ1qitZWfzerTEvmqDKIW5ePGE6YgMKFhReD0e03U67Fb55hi/Of8LO5rCC+
3B5y7QfqLYc0O+fQZMpiXKORU8U59lxvGml28S2PbAkTd3zfptoSeEd/IaDHKtE4pxWc5jBoUuYH
5uVzslXlv4AIztFPJusEZtNn4pqrrqMDzfSpZaZSAkQH2kpmmhWarfSJ74T/4Sc1dSFUp0Czp3Uh
vzSctJoK4C/LxATecdQorOwi2JH3HVZmFHn3awlhYUic5xzDR7lKU17GGvv0iaTDeNjzCtb7fYp7
MBkXQCTcEoADyZ03XUHnbeMZNtvJeK6QLseIJk0vJGG+n6Yj5drvUZyDWe9ADVdvNF3VIzlYgj8X
+fyJGLSiKPQn9hWE48fRdZkF50GXGTCuL59Pi2W3NgBVr1fdrSQDTTzrundgoX2XNuJwnciyx/j+
oc6fVF2jwXl5JAapf/ctqkYAJkM7xOv+hJgNdhU1/ybx9N7MhXQ9mGaJAg3TRP4a9K5BE8oPb+rt
nHapySTGlvOENnhe34KVc8eoTs0VXQVNOnjpEZk5XBArI+LYxq/iTKKPI92X8KuQ0GhQVk5NIxIT
8hMv+n4uUH/k8a1QJg+5uFWh/d3MqjR31wRjWbM5VrF14vR8AQ6lME2geL/jIRfPJen+Gllp+bDp
m+jmASTLcGmby78ik3V585A+o5SfBqP/awzMQeqaGvpkC4vsNjxatYNLvrjXwvKS1P/VtBltgluD
k0MGsly85j1Ve01qRNF92GaAqdEqPwT0XotRjg+ux0LvkC1sJPoAZ7186nCM2vC2YSg4hPY8+Lt9
7T7lXLcuWS0xoDZ5ALyvAnv2J3Bm6zIIHp9QI3Jg8bPRXJKG0Oy//0JSnMZ1kVCMc7gKo5U7p4Bd
a5HqO2Pz/W8CBZA47EsDrmVKBWWkBWWIZaWfAV/RpNJ0g/HpRRgdckg4Mtx35ImxQIj6BPAtAiEE
ytxXkPPNhsQonhDaSZ6QcO8Kq6emp6xNGrNdKfkBafkgUCfVnrR/WnWcZjrZjh2+hv4lg1BLdl8Z
aCkCgKog5Wmp2P+ivWTc1IKf8UUY72ojcz91y7FyejNULBR1dT+JPtiuzZvG1QvjSaHteVe7+uCq
LYKhWXMVc6Rlg97rKiWnbgZPfsTXe0vYctGEMq0CAfEzsKJ8UWkEjKnxqS0VvwZem7QMJQHCGf4j
WIHTsUfBoTxyEF83sqZfZ9IHDydAbzEXReKrvhh7Lrwl0Oi02K/YY5dd9vhqMd0puxX7e1s4QLIB
HplXvKui3UKei34YHt4VLE6HYMz6yU+MJslMMxrwffzcO9yDC7dbtwj3yuvD8Sihq9659eu0Dedx
ZM5WNrObcwJiaANs4sZOS/5Pimcw8klDPCStAyH7vnct4WmXR071HnN8fNANbR76/uVbwAjC6Zs3
yPJqa2lt6QkNBFCjwfWkRqEDz52+MUyL+P4FpVE4XdX8zfSdPI0vdB7w+D3FxL3bPu7qU6qfs9yi
rVav9TKH9sin6IWc3uChvqni/JjjOtkTXaeNxiw7HF21kpp5SIwLkwur4mKQhpvl2FU8jFPnbkky
89ru533cgq4NAvA57SQ/Ob1g7lCjbo/PmRkJiVc5MF2L+a/UWQ/gzCyVQ+oHeUCjLuKJ/qFbDMUy
5Z1nR1hjMCD2y5NltFEB72A/l0Tf54bYdoKTF3ZVgHjtDM2Kk4Y4SjuT1gP8lmkszJ9jk38IXV8F
indcXpKHBe3wLObc2v6iispapJsvfUMKZtVo19uHzlh95HGbu4IsanoiPk7r7Lw4SyBikvWSpn9X
Gz+cZMcVsD3rKRTyN17W0CRNwLBf6efBLSKXgFDOI7g2ts3vd8GXYv+YRHEybCQK+hKyMtWECMFh
M22EnBph9OOgCQZV2NBEx5+5CxuEFmm1hsT1HvcacpzR89gKBFGUHiAd4cP5J7ZmYC9kmuwubugO
xoOphDpvq9zHvhkrmUoZqlqtlvcCeq8OYb1K/ZMtzqjc3UJ+KcdjIJtZFD32g+PZFinW0mp7A/MJ
4XLJYaHfVTjnHw8GOxV5o9kajnNpT2x8cyF02kyWjQWKcD185qjL6BQfiVVQUQaqrFs+R5Yr8l17
ogN6hwhoNrVZwd+9KUwd33NehABl0yQHCiIGPQIrKuOo1VAmm2IW4GVgAyl3LeOV8XP7CyvuSssS
texB4lTBn1DALz+HUBDFi+bYuXtZsKLRsGbF8y47/3MgamQkhbV0dzHxaDJH/DRIdhhSUPwYrS3v
9sv8D3L9qp7zQ7OgoBQjCqT1IQLZwFkGq8D6wIuK3wnORxqRk4rUeOdBjUTkqbcgMkkC3DL92xG8
RJyPxBnH9Zy53OPZwZ0AEQfqPCUhjQJcLsIudLJtALLysHFZLJj0XNqRUIF02oDQo5SilNfqzinT
wDN9b27ZXBhMbMJFMFu58L+xBY4Tg3Q7DW74pLNWUPUgz59K5Ta9ps/Px3xM1Dp3hyYzFopzM/81
fHZf7ijbkdSwFOPI2deMaQa3HkReizSHK2bgQK/nZkB7wxwDfIDUSTI436RVSj/s0veg2QoRWiF4
vUOwmS618fC6h8HhSEZzrBD8iiGvd4Y8+a/3uwL+DxnGAETNhqNTu8Fq5fNvBYgGSXlRZmkkonMG
OMYBxoFiXl1Lv8VNMm2gh55uRTEqyQ8YEqREHZB7ilmcAqBVy58wDj1GC+4jCzlLjY0Sby8k7VHd
ZH9r2Kk4ZX9lMPRzx0BlRu9fSfx6fnc+y/6CASqfR2NegUWDcdtDLKoCd1Vo6Q7x+tGJHtwSHOQ2
S6gsoODe5mHt/w4Eq178aRmSPF9tRmu6Jwf8OP3qgLdCrJ1nBSOg5ZBXEZpJRyN7mFTjWROi/1jh
pAe9LDZ3B5NDFQhfAsmySSogz7DjPFl4gPvYJs2yf4cGHEwGtRI0YCCnpaEahwYqtd9cJ9bEF4V3
HaEkNC557xoRQyi+tVtRfB0kDy9NPotIAz1DyfDG0YI2SiaUVA/1u4mYSIO6ZLVFwcnLiHU9CUqQ
XMbXQ3V0snMLzhQzfLGueysvrZaJfLxZbg+GNW2HhaaER3wQPPMfzKxB3Ydx2kAt/Y0ZosYFvd62
zTRbRIS9HGZO3vLsK1lmtUWQnSQkY9VVnJwvrGCYvCqlkto/HVJG9VdIoUCVLyJQAKIUQiU1+URu
8eGRQKAJHsSsc1epqdRWAvrV1WxH/LwFMjOb4wMOZdx8d+/S2dj7Z2U6nUuN2EqKaIFOKkanA0C5
u/ViQweTrB5Gtit99XsIdg167pdepxyFbxapLeuCdiLIS086D7zZZNspUpWWUAUMrvGy0B1DDW/p
ZCEv0wbt1ysC6450+GEgychdpLMO/E2HlUZ9hfwwb7oGNtFK7GMfnMamOdGktS+b4c0hCvcg4Xyr
zsoicZ8nPvqDn0a00zfls8mY+dq/j8zls67wmKRcPQXMZWqFoqd+e7/lqY/ueBlrkblcPQSRYNAt
3TGxJAbY7WfamySt5PBG8GwZSg8vJcbpK2oIowh+VkXZNSuGrUuByP+qalPdoSdvy80XbOngSNyM
KBPy/1Q08qQ/AJbqwRAjK8+6p3m+jdtKaYqf2BgdI/a5il22P6XVq2ZWGdSGKnWiwqkuNMtAfnb9
SoYj2QxyA021POmTMaWTlmiyksC0sSZnKvnpmaNUEP42AwZMJgfCfvG/NeRngqOGpAlRbtCCofce
wawpemMu8ZssBwcusB5K9qIuVA8UkE/e1XvEMJYbHrkuGPsCsCi751DZpFvpYaz19znceyb5t+2r
U4g32rUANdA89+LhIti0nSa5w4LVAJjN6NRGcFIEJ/ZNierS9JA/JSw8ch7Y8QcoefGfBzDTGCJn
h/Y/xhQba/zhZEw5oYfRkwovKxX56PzFi+6b4w14BunF4Vb8LqO3LNyqquiNNAWe9m5xeT4YuwdB
t7cRaY8xWdmd/PmHKsvtJeSvwT4I7d889TKXkvqI5NdWGh0Q15w+NJqclRwfF8QOr5s6l/63hmF2
kfOAuHZIZIrFBIhFDAkEw7y7hopuLS89vL77omRl4tWImeUIq2UpFEF5MJtbpt2J+8tEBJlUjMpi
wFCKPSITyyR/0PhaOJCYIbh1aeqmx25zwxFpr0MbQvPlRNgkSGhD0yTOggF1REGlzIGa7kCgs9LW
6gFcKZvbMgtpMzMyed+W7tzJf7K3OKKNmqKBCY3cFZrNVYLis5mXzKcAWa+31bVpiuEYDmBVqR4y
/5Kv/IjO2L2bxxX+7hwYt+N015tSabWKXLGAN4s9yBSjw5YrHv0RMgH/Ij8CA2Q9QDPtO7TfJAME
kzOk6zeDI+5pn6JVoQcY2toGXi7YZJhwRj7soLLgM5QtMfMfSzeRlsZAkVX3flxxasuPBDAleQo5
J2xywFEgHbPHmLXgCNMbGVkH23cYgRFju17opMzUuES1DTLwBllSSSaaYPhu25cIKuilVGfKBgY+
h6acauZ2vfzjmh1Q+Z62WxgMBHmlPGLpkROzN2j48JBZTwaxVEFsKAGo5YS+renCBgFdmeMn3iRq
U0VyJhnpTavhV7Qm3egBuA21tKO18uz/v/fgOJfCYdIvn4E+z4xVmkF7Ouz9jBpUy4wsU+Diqf+c
WN4Zqph0xMgOn/U8OlLTNWec/mkwq9HuqSK7esTyfveLKHc9+vhX2ALeRJ8loBvS9XdC/+vlsq0+
aG+8/3jlBukmM5xq/m1iPsgwO/s0+7E//VKq0B6TxsXFczJUU9tmPAc5w3uHBB3l1pMMF48rsbwn
2BjhmVaimmgUVQoBWbg2i4Pz2e5TVvgf0FOMdc7M1F4oCOpjDY1eSb775Aw7lm7jxXiEeQIM2iqf
5Ne6LQECj4xmRyE+n/E4ifHRSEdJ2mQaOf8AdS6KYzD/5DqnjU5+qOgLa3oHU5VdYdb44z5DxNv4
0wmqvlcTDnWEvHByPsow3ktUOQ/Hm48QDN3Ycq1rSKCPpwym7QQJMQyXLbHa4HY8df5Ib7FSWgnm
52jb++kOSeKdYFPSK75C0AfABnMf8Ym7QYiAgURNFScyiQ9/tP8/oq6JshBbqueHgPcazIPmfSjI
gh29v6efvv2OdXkorKWiLNcazY9aJysRtq0obr7QVVoeGQsZmnx2maWkQHgRRO1Z0ANvsU6uuR7o
PVF/K0tsnt4bky0xB3QNg1prJX9o6XrqqjxEYF2tmvulufq4gEZRxO99pN6XmoEFSfBpwvgeqKt7
lz829P0ENkG791TaLmJ+b7DkiEXZDtmdimkhfNBEyUSAYu9pWEeAViWBjL9te7/9tQYWJY0dLmPz
kzBpFQnRN55so0ooADAIzZnaXjQEw6J0EGBCSId/sELnIL9hLFz97k5fha2AC/uFBKGv2YwvAqdW
zC9D4+nmmTEDNNi2xMbaHFQowJQRrwGkWmNKSS4n/VfKE5AoI9cPh4VvQTYjkDnEeoqsE3uoiJED
E/qmq3DLx34mQmfx4W1ZAz/rsNxIwxCH78tFC31H7S++lZWKwBKAQengl6TNP++WPIwXGhL1dzED
S4w3+RjwnHvL3Jo/MVmmNr1OVMrC54jrJ/ALTbHkU3k33WtFLTo9WGBnO09XX4+QB5YPNO6zrUFg
aD3UW3/iJ47XTLKnQvEJBg9m4Nb9XU31tCrgrGZYDriJF6VzMhsDKd5uq02ByZusrc14Nfj/3mBZ
7WDbp1P0CFcp3Nm7fpjnpnjwHLLqHIgB8m2+wsRCxjYUqAC+axNxPG36l2pfWXz9AQ6ndABap0s8
YFNnikQC5gI0rnpKRJJ35sATOJRUjZy42kAw+3TrX0I4WVYOjj5z2mQ61cpTNThX7RBBIkFKPsJ2
FcqLg60llDJxAYP3XoQVvkH9dNFLPtfhd8UcUeMUD4zutlDhSnpUZ6u0gilbzvd5EjFkVyDcSrbt
OZ07DdgvnjoAUngY5VaQ03jG1Nzg8x5vKA8yKlp1ZqBfD4VE2KwSCUPaCJpgkL5YaSgXZb3o4Hf/
2l9JBQ0Zn/uyI9SP9LN3wncbaPBiY2ywtHjWljWAe1Fc1Tl5S7GB5UExKrX0jVDZNFJhkcx47Mij
Uq7mfcuQxb3S1J3KQ8EmoCiYJhavwRA111kh1vqnn2X37zv0D87ewulIEGMpxJozTD1bAFRlbJcg
78zck8TPKD1CjANJIJn2qJe+qnoGiStwJ+b6iUMEF7zIJud9ec2nSf8WM0MjZR13z2HkV+6FrILk
tNEZt5EbtX9I3oXATEs92zzn+bVJfH+XcUIog/FzkxA2kAm3yGccYSmZ8K1XSbL28Aqd1KSs+FXl
efyR642Tulcbshb5brwclGi6XOeO25Bp1Qb5zvwDwg7OfmREbaU5E7kHv7dQuZ8Fjyg+Hnj7uaB/
TZf2meZskHC6+ayzD1CRdsu9Pu97dTULrQ1f2WkLEwS8E8iQowLMtSVfWUXfa05PCawv+925lUsI
VhdOb9AITMJvK+PSLXAPmtBF2ohQg1/kb7hTvAqsGJ+Ohj9tFmiX6ib16wfKzMQYVajy5mnuiYgH
wGif887P+9LFenONFdFBLEj6iV1DiluWQz4XkVfmw5HtZ1BSo8y91zn3+6gkNXLvsay5Z1tR5ADO
6xWQq+b57RINm7PV5QCgiN+E9r5BxdPstkY/u/oOu9jUNF/3ihyvF8BG5Oio/26xWmFve4MCg+QZ
DOx8wD8TlKphaQf66yxOVPPenqfZMJoysnMzJVG9U8zYTD9KOrPKlvUgjAzJ5FDOsb/2XHHgX3aD
DgPAlCfvgVQV/t4nDzFD3aVLUTe8LT/Y2jtP9bqkQqnX494WMMeOfMbvgFiLvYv0YCEiEGsiQm11
TwngFN1kjMr5WeKy7CWIfn96P+BzISBbJp0NYSiGnSBF+QQcgJHomQJpKvmaKabbduvc7lzUA5OS
C6l29b+bg8VHujyj7kCa7DUYOgyjIaphLuaH7F1223s/IqUugtujq2494EAjFcvDw49WjMuaHVWh
F4O6XbNa+MxcJOW2GwnqRZt7eUqYYployr8bwSKFuoKzMdkzXG9fwaNm2HWYjqgd01/kR7KvhNxN
3+EIvI6UZv5vgcQKU0hP6qyevqFlaTbmETwZ3kDtLkj8fhxtTJLV5njgVi76vdvW/fc8NDU+7gHP
QVlRidAeIevtIcnyPC9gw04RDS4fP/GvANSSfI6hNkbS0XODQn6bZTk4ELPXlzhaR3McflCoDJ3y
gzUOccdDhETDTgRosulGLs2HBe+ePpE+Nn2/CzVmdZ0wIlLFNuHhb61f1BP1OZj7boTUwzi28jfl
5DK9XV0kvbZE/wNVGo0/H9tqO9z4DFaBGFReZ88Iya02JMjnQBrupnYa5TUgYSzndg3rXJWkUC7F
sfqQ6DFU6gP9tQm5Z9RwW+WT8zGGBowyLd+fMxjJ3hM/UXmF26zZaJoiqV2meVnNxP89I1q+ChGF
YzdYVnOtWciczX03GRZMiLjLJkwyBOXTM2k/MAYdxzesmq+UKb5lMtNibqz1IMjw/BTcKJXoKLCx
RgvpTudi0uEsKWlXAYPdCVsyk30OWyuZxUaYzx2crnGm/QuuWaVVOQiLSm/xP4s3VXFsXKx4qrvf
MKtv56I4KtIfoZEcGgjtTyV4a0T0VNMggjVxA2qY/SHf8Jlu/YyATVuyZJPk0Xoe5YGWOp2yFCVH
gXaNptKRYCKAcnZ0a+7LkuX+zQwmO8Ur98/cEGrgsbhg5uERA3NuCPkb1ORIkcnz70zfiHV5hMHg
n3PJO8kxw4mcjucMa+JL1cAH++apHQZzQB4UOzexD+MvM+EpC9T6Ek9s0tzD1VIeUmkZhfdHaUUd
xj73ma2esUIlA81bLwkkIaPYDjy6+alsZG0cozNfZiWKtWZ+aKzafAbJUwoJDQBX1VwOUGnNPNsK
J89qd8MRSGjzwZgXJUaDn539yYAQf8BGr2uFwTqRGTrH88RrDbEyOZWfNeVfULku+3ZDg3pxfAnd
viZ9/CePp8XTUOpMEYDJzBDPBQN1dyCUerax4aZZOdMCXOtJMPy/bscUIdaBOkXCMLI0AMq81JJW
56g1b7UN5E6yFtcH2IWRba7Du+C7SZwZ/MkpTnzoL0wNc7IReYSmuesnG7M39KhCN1rDxOgmSNB2
m9dVaejKIqzN8dn4grV3VYeZUTm0avqUXv/+1tY4fu2AikZA1ds5pm+iCCDH0hYgyl+9xBlxh/Vm
ruAN1dN8mdgtrk/fDYDBpt/Jmfd1eB2bVz1jeoIpV8k9I/ZIr9q5v8JE9LV4QYeKAku17m8lZEsu
0R9CKwfcLkMbBYR6gw4952xufZCt49K1ZyX8MnNk5j5W1HiD3e+IW92AWu//geIMW7iEZIRMa7nO
03vtKbM4RwipJszCSyrL78p2DNBIqWfgXFKXqizNPzVReVlMM1TXfh5blhi72oOGfzGKnB8jemv1
jh/ZBiwya4n8Gto2O2rXQ4b47EqikjoRRPbJAbSyiF9zkfDkw7TTh7U4bOiJ9w347dI0ByD7vl7R
Kwef8xnaoGnWlW04NV4ZT+fFHMnzEkATRFXnoRkZZMoQG/tT2Hymeqohvt0Of+nzp8qeIV6Zy62P
Vd2NlmOrujZ0sjNdVRRj1wrS6bFpNekoyvetyq3HLIzPDyhIKjQErMRLBPmSwhi0aVKn+Xq0r6Os
wVIUrpN/T1WJxi8xshPiGCWvRTYOTOMZfPdiGn7LB4DDhE6fiEOloTgCFJiyBh1OYkK6hJ0iaBxy
ON1Vt7Q6sVF0zf+F5hggPs8P/pZlduOyvol5Flqi9zBcm48m3kjuoCQqinMQ3PmpI4H7r26w0EBt
eXiX3P+oWdXwRVkCFZjs/pYlrzeDvsymlMnRHot+ui355vNg/hmzxDYMkgskTg0wJjI8Cv7LfAJe
KZ2K7HR/RrkU4Luf8cdqBHSxXr+1OZlA0m+xKgiIypzf6W932hb7fhDPhs3t0pSwOosDtSAn2rCq
GX6vdwPYbpchZ9wFe/Y+P5C8ibHT5SmS8kDtbMp3Sdpl0QP4W+auHMglZIKuOt1LC1nwbH6U6Xj+
7mp1YXcQlUP0oC7wINXH2/f8DUZwBhGPg/AKBoi+rCGz4Sq54xOeCOx9dhbW4l7At0s9euqsigfL
hvdvUUnS1oYhYvMbNTw1SiBK6o/cmQogEkbYna35DwJ1JwRThsmMn42WLyKQ4aXtGSozWhJp2Jdm
YaM8e8BN6q7OzKUBbnINYetqxOwzWhBj/gQeWExWMItWKZL6MbBVAcRbvQvwAupputRuOuRRJGqR
blJ0hFPhVpXtzWvhcfhmu6vOG3jZsEvx0l4+f9vziNB2+nI44KkjDx4uFIo/ZjDG9GUzsBUJzjsm
gAaek0eCssSwjYCBmKzhEmpvdfBTxn7pZJnoQ2NFhjq7BSatcliOtG2SH287VdBXHOn5Ff1INksF
HZaTdZLhdqlSCL0g5vSRfm6LuPHBovaiOWqoVb8G9fyEcmgOaes7S1DN+z23EOv2ArUmTYSj5fLu
44IOdzZM2a5WGAFgZ2ydJRIvNqMfyjkbq6zZG49iUs3iWYYjFHVovMNdAsqYgIKlHg/MMgAE8UXA
vRSjXo+e9pvqwlMV0JfWJNB85/yH0huNdDyNbR657kaAgZnDWVdepwY/DHty4B4xGoDVJud9tdaK
PKDfgqXTHRpRP/hBsPCmOruGndN5c/Gt2eeOvkEql9KNzgA5GXNaR95hHDSbY9COB89g/+9NEHpl
vO7M1OKpVGow0bFwwT+yqYKEY0U/57xj3YRLJq8jtdvUAX3p/TfOvgaafwXW8/QCZYhG2IxfgOBw
T6hFQTwoz94O/H+nkBl354YINZSVkpv6PX9l5SvcDtOlciXl2TTz2liBGXbjbNVugrhKqM7ME39g
sooFfgSIZsIPL2hOMywa4pQ1OX7Rwsp/m4SS9BpRu8KxFDdJ5t5jxFaArqI9Q3J4BeJ8MIAIkuFh
57239q4fc4ytrDxXhgQtGOcgtvMXr0di5y7drOhY6m7L1U17xMEbsrv1N7L72n7Uozf/0cZmQps7
oLQGNa8cXqf2jjYOILWVnWfoGfhWlK26OehB3oiqBMcGL8IJtmZP8FrL/tjHJdA/xY/QRwmeYmnn
+AXgsE7GynPpLfbbiB+SIQK344fNywMiyq8o3+ZFYZNrAiDct1L8+UnfpffmMSYVruMg0EMJFbP0
Vkztk3vl/s8/DEWrXXuW/x13ggiAJopawsnb2Tpovus61CNMlfX5Y9sVI5kySH5S5HBpy6RK36vp
TTOqtkVbhIxX4w21plmNGgKdl8azfUtsi6XQqZrmVZOgfpxRRDkBzABjU9stvx1yG6jMDJ7fq3/o
uD78PJx9AZ6oAXi/8BuAfL9u7+rjmw8Z6Y0tKJbYb2x986VP77p6bwttFaRvBQqfmkFIhWCMNB4u
fgihdWcYUtovPEvB0sX3CXl5InvRM6u6IkFUqzqov7TFl/y3VFw7Vf2ekxRMgafHgz30Y7MOjCTG
9TvKgH+zvzxcTHHLXzaD/R3fR9Ej/3/WWc0HYpadWaxvoDQdN/A+ibrZTq72kWrZYkog3d3C3GnU
iKxdQ18Te+dVk/6mxg2RXzF8KxwmzON3C6EqwGsjiBWQpMlcdbtRU4LBH7SETp44jdfhik48HKCx
9VRFmZwb/hdIcr5zppdOFxCG1nKPFasuz6Ol3Xxp9TnAjLRgRpMowSF9uB8sa+fg9h2Opc/K37L+
7cHG6q3gy/u7YMdsHdms+yao58laDTiB7M1VKC/NWd5pzX4gre0DyMF/FkmtDsD/vQBPc0nlLBM1
kIthHYZyqBFobghp8rEAey2l7H+OvoRdwvyNj3VLuwEeikbO0Ns0zY2aRUQ5aFpfmZCU/jBLpAbB
8AblXUL0jbc0slWSPi4Mg4XpxKAeN+gex1yHQgrD0MM6HVSl+LL9CVb6Ygo3zJoZ3YZYfxBT2wcF
udMdXXWW4lvsKXloip4V9RD/Sc6uvix84kAElki7KP5tlktRPNJiXKXCfXZdBBJToxvN1qV8Mr9Y
jbrMHd2NRWovTTSSJiyCYImTGMxNmjSPpT4psMmF6JI3xG5KM6Exv/7SAPnKJTkojd/xBw7yAIxX
0IUZIwHX9rxUzE0LJ1MrN14KAszum9YXEad5yhYAyvSPmE5UaTEaWx9SOWumPZXnh56Ug0Wn2vCA
/i2d1N9COOCgc9PZNBbQ6WQItA6O0sltk1ZqlNpxUEkgWMhOFYHBlpbpiAsqD3BBNTWpKN3hi/am
HlEtYYoorJ8BD9fdbjfbHobbyADit2DmZDPJST7uOLYqw/L798UNfxMencK8ZWzHJbkQFrnPFpVQ
I7EQHstYo+fvZ4UQd+zXARBUdSQ42aiOZl9awVR2jpWA5DaCoeD46pwV3zkq4heUmYiUkW89sdTs
xxx+XRZBP030zZQs+FR7CLY4NTuY+P6MOd/Acy3fqtU3RvdPgGNkdF/+5FnLi9ppXbCKmTJocHIB
aQltnSjW3YV6p5om5uYUa4MZwkUIr8kzN1IAyxZyZ9B65LwI8hP9Bf4RNC0MdAhc08yXX79DfLeN
yFYzQdDRw6Ozr20Biu8jiVkCw2CUjq/a7kDrQGn7DSyub1rVU2RtD8DzF5a3R7EbTpvnSWuZCsob
aFOzQlhYJ7dLDawa6hA/4JhqDXWhK85c9YlRrGB7U4ajjCXiuZSHlrYH308bYcHD4+7LXSdmbk+O
urCyf7FWHQi5T17EYfHBsCEbHKljkNE6AWItMu3HsXZS2goV9Hq1SA6YRYtL89+LlUASIfDm27UG
3djiBtEzDnKhpSVmP/DkuyGRputsKP7Xpt/zyV7z2JBF/MG17J9gv1CcKHsLqTKGhzHs5lnlKf6c
qzpf55mOukPh4gLHHVXxrtJsPr5d5EPHZLl5MNpLybuNhAQr611nn/dKsYGafMBbAltuQNAEBLaO
GePOOfrB1+QnxMXyjTTiz+/L1UXVNT05mnOq6kiarVuV7l7WAZLBPBrtHXGJuK8GXgx8c/FWQ9Gw
d3WG+ZAlbhtsz+WrlcBGywErpy05lMd8J7ey1KQ7a4cdtjcRVM5/iRPUqBzFKgEMZ5mShv8diiUD
pMDOVUXSuHDsJF2Aqp0ZJil1ZvEHXVGfJcJmo5bgqL80phpRdMzxdzX9073SX1vlh/bHO46dm8mU
odnbCovvE/pT089gkPRiWmjn5ATrhc5oRDdNs8DYjUZztXVRg89BAsk8UCoCizM+WyShf5UBAV7z
nsISixOzVM/TscyIgfKPOqBVMiSMcJhqJxmGkOt8C1nugM3HKDW8mfFIDyJ0nHutbxq42zHz19BX
jPDqp0ItDIRLHtjES+1BJ6ANSb9iOFAa/mAM4KvD1qhCM2MDacnTwIt7U9Od8cjfNjWZVrTEJ1ZL
V1eG26IN4WjJLTHPYQJXv4iXSsxWSvyBCK5kBqsUhwZHYukOkZ3NdZv8TQtcKU6Bs2vigGhSR+Km
/oQW4wn+JkpcpUL1xPDOp1hEuAs1ALRxzI5Jna6La63/5haD4PSzaukiayL/QSnIPRElQnDv6JCV
6j7BIrJkn22CaP7fLqWHGZYc5T9mcAYcUIpLT3CoOvbHa8Q/05koBnOVT0P9JXYDA3UhdUhFX3jx
8IY5YgDMhBHAPERh4c9ngXWQV8X6fTcg10xEWVulWlcxXj1igSyzmSW/dFR24z/qqmeCQdv1w/y3
8jvQRr1q+VuSoPgiB7oxZtXl99Q9sXiy6tYP/EIyF8rwiycuBKB4Pt3N5IRtC83AGE/Nl+uKL+vY
cdG3a54PNtxqwbdimaDdZqUOJbp9/UiDZs298b9icjExXhmdGrurhwv3g3FwxV9BQ+5j8WOber62
6PPWRSp8huhsMhPuhEblXtqp3j8OhkXJ/BZlVMseC6gA0Cwy4/cknaSdZoIULKdZV4rkXyyIxaIa
2Mj9oyh9vIIo8v/MZZYsWgR2eEBBAwBW7Yb2Wz00ENLdiN+TtaUG6szDssF040k9L9s/nPBEpZl5
SYRCklrHcDTb3OXEpOHHTOVoMODFQos6/t3+0LTlzTp8yZcKy2j9LL67di8++iFMTLWjYrwYk5so
yugDWFdmZf1Uuy6VKf4FBgXvtVyD27aqxhMdX2Gk6CN9a+hJr6cpt7HKQ7od6uWkmhBHMuuIqZeH
s5+l9pb/aKnNzXg0CPEdjJ+E9ieTowcwFZ5bqWPS+b9uEix0zFuYfXYJ815QJKSpI1m2C2/iXMb/
QG3Y9ivGJxyJxwAXnYE3EOimJ4BdD7d2cNl0Kprzqk7r/j95nL+FnpezpoqkTidyKqUPqQ0PGZ8Y
EQVtfMW2QyzWEHxMt/c1dVeDBvQPdYCnZz5Gc+0vGlSlHmgBy08w9OvL+dy+C99J6DDoS4nRR1lz
fGgp227xlBJAGHg+OOqQW4a24ShM1VNUtTrH8i8J8kD2j/bN5a/ldLEdeyZn8P0SCghEJmqZzfkq
0U8dvQtWK1/qIApmsHS7HLjEXSCy9oZyHG7qN8Onx3tOzzqor5ayqyzGMuA9btsZaHXZh2/ky8Vw
GsAVqvebznXHQOkJgjanMLLotxwzc5CNZg1ULaiA7LxXXzbhbUuVy6SNg343o1zEPyHVZsDc286f
Q2pManvgshUeZZ+oXBQAAqaqIwYsd0SbFDFNpNWgaOkC/wjt8+z3GSZ1hF5RXFaY+6KQe+nJ59+T
beqkWVubWm2cXbg1IYWQwDgZbF2F1i69F/5reFTgOgyNf6xhLQtiupY4KsdZ8Vk6dgn//6excU6r
Ha2uzxdYV2PSr7EcKX4JSig9H2Qm0Xy5Ub3mOIouMXCYXvvXNB4vNcRSrc40CNVSgdyijChze0pc
dRvRloE7jLVyZ7z3c2mKO4bQhwJyMbHI/qWLN0z7raS58uFFRXA1oyJaNtGpHBN9HSIM6i2DHWvO
O517JEDjoLUO8prv4W0b8j4xdy+BIZeImIaXtnIguV+YKSqhAvRjUmEyJXU1HO0JmpeLEV9igQAX
MaY1EezOOaoiCJJq75+svhmytfDszIuBa9Mp3d+XdNqMze/7/Kw9n7F4yoaifffC1EJRNJUtSuLt
qc4ijt0j+e3d33zQRtJpc+MkKtmxv/bOZCoTcFDrMZic8zqV5d5Z9CG8gdxCkh3X2PtjSV/FwEhm
1Qm9k6Xu559ztAE/rmyc8+mkgdWWalOvkS4XyaAJD28ry+10C/ybNq/QZgXytrfo0/rbHELslOeP
xHZDDm1yTZ4u2YoonZCfYQmZcUFudrpjiSqn1i1906CLYjfjNescYry6/1ZWTyAGYU96Dru7XPgK
zgwTW4k35t0/Gx7KxKo4jQk93lhDiUIsg3ddCg0bECqe8Pd/aJ4coqH6LT7Vn6UcqlfW2kiETbBm
ATMbFbfY/ABbUQMi86Jd/xGEc+qXEo3VXDDrc2dT1lnwqvORBPGVwO4admaRRQ6Wm5uaW658LWN4
y3VJR7c1nYoHPCPGIm8WEtSGrIBSZXZ0f6xGVBaJ4+bbIVnDRtR2e4VNFhmv8BGM2BAUxvn07o/9
E6grKWs2+Ot6MV/jl7RxCZNUbVhc+Z3p4HqIowDpX0qk9pquyhXEBw/uOWmgrjNVyzxwvbS+mNp7
LHW44F/4N2imyMDAFAearW5SKAfXCv0xwglSmBoi5JDVLOoIxg6ZtmobeAhFjyyPv1V7f7ULgIno
mjoA/7O1h333zQ0Ax6PM42S6bkVx7/OzfB/P67xAE0acpg0bs4Zu/uc8+Vc6VKp4pmD7e7rZ0oKj
/z2QcfEI2jk3wZ1ej3BckMrvU65E3b+3RP9+vemRmTOkvCHmGSL3aPaNFwte1ukzn/JgikYYaaku
ED3HQ3UdX5nX27h7DTMZS008Dj+K3oprjN130d2O5KtsQyAnuJNV7UKNeZ+w5nN80rt4DjQJcbtG
ao8RDQYqtYZfpHR/z/zCI33PFXX0/9RbicR1cDwR5UkpJaUNmx2rjJH/FPDSUU1OqjVYOaqixPhq
MPhdK6wT7SJ4UC22b5TZxsRrHJds3f0t7wLKBCjq5qBuhJYJBOIRULcFvwsHeSpTeexam2vg5iqT
fOsmQWxAQnWc97FeA8gHhgdHrBvsKxiCOc6jrvfAVjgsbg0TsXk1gqlhkxt0pwhkYLKSd9bk20wj
gQ05y/LqGzoe6Raws77xZvcr4Erdj63KaPqUuBCBqgPo4oUefuZ9LS8sRnUByrv2P8is855MsaLs
g7+TOxle6Ik/ANuR5KEcf7rYI6CFlzgSu2eyXBWoaQ1EC7cq2jmalHkj1ZafFN5gccxRnICJrp97
irhj8C9VqSQnYtIRSLyBwBkuka/YVUZvTAbTQXtixEYyB9/yqMrTpCuzP5HSBLoqyANv0jKorWRo
gB+Uzd5BXRpxUO0ut5fCmLHJDRMtGeWc3LgyUXR/oIC8Rawmoq410LUN+BBACWx1/oaMz5+QdkT4
ZMWbOZHz+ebR1SwD2ArywMnS0fofsUSJvXQxDIsiY36MHC9OrIMgPV5pbGamlYkO5aFISV57EfRd
VkuL9nhq5GcHUfvXLq4+n8MAph3FmVYLBY5BYovJae/cVU2mSzeURvFC0XXEXdjht9UkuebWZiL4
jswDXj1sqDMcSbLcu7VJ9hvcSlW6txkJiJww3UcDhZry2OAdai62uNZ0JgOqzmEdo/8RU2+KpzjM
xD5eBarMBp5K0DjGbq5MMjVht7xEM8GR2jZTO/kG7uz42xn05Sl5zWGOcgr2UJr715/8qemYoFaZ
9+D5cLXgCg+LhRem7dtL4j221cLvKNmcrdmvJWeH4iAksklN8nQN3iPCdt0Pk61UFcTVgio97Omy
ulgovwTBUjwDN9jSDVjapyUe1pX+ApHjZdQZw31UgzSE08FKyHsRdUHCpi7s24SOM2dAQ+0ZHxV+
z8f/2DlvQBQzqP507oqv+5KmNmbXq7FDxJ2l4S0k++W+m+tNTnippR57Uy3B3Qnn9qkJpUjo7Fd2
znhGgml4IJ0Y2bfUEtXX0USx+MXxf7Fb43SdcfwOeyTT4YGcX9sQrT48JHjeALQRZeijsWrJB8Eu
LDc8wlTYXOz5N+hzkQ7YE7pWODDEkGv1jkCadqJLw8zH64UZ/iBNZjz21HbUVsOgzJAl7bOZinx8
JzRlahk2OX8jcy36FfZV7yLsQ5G2T9PfH4G4rSMnj2/+zgpCuobiBAaY0yvMu9QeIegFkrqM1W0f
BwAw4TxeQSs9FEiZ5w/Fq7wepR86zHAg/jVodd3Ll1IjFfo37ahpKmsU/s42u0ydZOoLOVtOfQF3
U7hxthLJCDFRD5wH8vsuI6Py6CSTY65cdGiNXI2S9idzA6UCB5wl3OdBXQeLq4VguwsUhiWpczt5
YaQ7BdB4P6Lm93wRDfA4ABWr1irlyMnhES/tdChJKyq0jVwtJuh7K8FpesTaVN13gIz+kN77z7GE
XixBYhK4wd7aXYXrt6BosT6v67M32ounF5PhSuW3l4pfsnFCXV/AOtOR8ZIkG+43ciW+XSK9X4Pr
fu3tkKMTup0rQUjFznwDle3tJoJVdCUx7PguWJFtu7QPGyJduh6wwOuKBeEcj32T3jBIzOd4MztZ
2urN7l+dVETSiYdllkvm60kicJ2Cb++ClaOkSPIdt39le8o01lwmd55JB1KkUzGI0eXwE0NTDxod
BDG8Oa5DhTZOF1Bo51qThvnbDANuo1XT/uN6mBGYcfKMF13iUceni1rD77RYLns4g6zXfi4TFbW+
uY0FSpK7zw1yUGnuj75ZWhUOtglqYroTsUx5gjZPTiXD8RJXbkpGzEObPIsPsDSeEbAme0xlo6Uz
Fpgbge9AWh+ErHwsjNL1CIvyy765aMJKHXPM2gWbyG4DjMqS8f5NU1apAsEtLnnZrQfowI0FGaZe
GGa/el6HEgwad9veRK4QFxldmtpGPxhmb3iBw6Qux9fRVeNUVz1PvTyA2vHuHPJktQ+lOO+Tkqy8
vDklJnrLyHe5oy+0RkHi2ucKAoC7fA8unB0wYi8WuEdn+xhdgG4rZwBFaEuaYQhGLngqFrhMsXg+
c6TrA8tE3mBd8VEKs/owNiCEpguy49HBLZrTvLmD3iaDvR/O6Zccg75P47FzImkKmIwYvIlK9ljn
mX+CvM6T6eUHnYFVUiLBVtgTPbNpMPwQuW3K5brW2rz2l8yHzsFExcq0+b2KmlXAXPrRwUX/4c+X
4KOk/z0kB75AGcFbmGv9VRIXrEUbxM7OfI4VY75PqepGQZIC0jwSvmXiGG/j+Wi5C5Z/FK1+qdVZ
0qVDJas/cBHG5itID+fhqmaxeKrTA5JP3nAjz1Aqt50mqwHa0M/Z8Puv8sN2fY7JUzDCLUj+GaM2
qdKyYdLd0cYip79HJxydkamVavxEzSvpRPShxK9hpi4L1OcWXna/wAXx1iD2kssylHhprifY50VU
SYvv0upFJtaXltfO+93MfXo7JmPcliwKq82/cgm5bEu9eXASuEJYWShQx1zZaHo6yn8cJrx4xiAv
O/LVa8ADcFuQ5WrNtSd1iddB0uQwgOp1boGwVm5VM3nTGz0ubd4wcbbYPndvcosLiCmFrSkctwkl
OgiuvGgDWq8QxsKoGXC0Uf2bmdjTum7DxvW8sUkpMXOgtevOiE4ADEskx1FiOAjwNtRAsTBLdoRC
0Hw3zJJaiVIHRlqEFuwIerxGCS4I2CVXROC7CP2SUo4aW8YgiIIBeSsRdAnZu4ZYIgc3oO6z2hk9
Pqpxjnen/tmBfd3VG1IX9eguY7FpofmKGqSui9LatFps1qeLUfXKZB3Giq2JxxXHL6aI4N0pIRos
qHj1bH21sdI0i7jRShNY7HMW2UHsEB/waFMqn9eitvt89vpI8Z/IpJgC9dXZ6o7dJ4rNun3uruxw
4JN14K84mB4nww57oe16tT0ZyTRFFm1OiuG77COgMReIPwfjy2G29nkg+WJ8n267d0Z9TFtucShL
rJCa9CLkD1GfUW61TTZ8/c6p2cYwHUhxsjvIbx7KlULdP37deQMi4afaHsObpqKLC5yKWBexRKtF
3MHpbvrGEyyE5yOdgl3d+rOfwAArsfK4qpA1TY8us6jHiXroO4Qt3tkuNDn4t0+p2VVMkQwQHG21
pFUwfzrEOWjkGLWkqe/BoAly3DcQDK6ZI69gVmQVnliactvb/Lvwk/2gdgGpWtTrXcA6MQGxl9Us
yV85Q76e/YoRWWT+pmjat2xfbuFDSXy79GNJngN9hD1pt4nzdPSKE+a3RxR4SNuruKp4JGYb0MQ0
OmUzICwfWwZly+YPkuxiCm9OOuzyij+5vF9Zc71eQKb/yttTA4+H/l2SuO2Usbh/YXkSOq8Gn7kf
1G1GjC+fD3tMHiB03nbk1iSkAfoQ5VBWWUGWg88Y2iFNWv8OjAt+mk7EbX8U/cqjiIHYKe2/O+yL
stOjXKsk/Z6maFvGuqHiUi/vEakvU9Li1nnKPw/XjoSM8BZM+Iob4hHYaJu4Ls0XO2nfucr2yoPH
P1Gq+UGHSa37uKiCfKSrKQogL/cY28UiRoHlLHynISiVMv/ndhQot2w6VLo9snSNEgHfqM5ZDtAj
K66FmK62CkwiQD0+Ae+KENeGt0lpuD3WmfA0VROtumL4OGIAIxnRjuaqUoAQrUvy5HM0a1ACGfF4
m+wNnx2YszI9yph1JwtWV8xYp8HDl6J+lUhMuGcBuh0WE+NYqToBg14xJEaLQyXhpt2ohDiUBRvB
PeqE11M2RTRhjcQ+WUN+pEVzHQ9UYA262t7IHpCUYtEX1sXgnrtuW4THMG2iS2WbzlrJwV2FSIqZ
NJiDHunAK8kuL9iE5j3KhTvr0GErE4qU9Hih6XUrUze3K0+3pEoeWtB+Bb+1vj7/3LQzbMmEpIr4
Fq4t6mXGiHIYWjLnDVkB0chl/B54LzXVn4rvJJ32NawpNv3IUUWoX+NsdDgPeS/uKrIqxYqk4OBf
+pCUfEfXIKCwR/azqBguS7j2HW2vjpHGFSceqejnXve+dvIBIANQm1XBhRoJD14CPKExbVcBAyIt
y4LExCMQu+vLCu3gnc4h2nxmdjr1BYBhaP5JzNjOp2RW202BdHhx84nxpiuvierGegABSZ5FZW5o
BiTY7C7kHvv09qS+9DXQaiB2oRZngJz3qqW+MQc6CnHKMhe5R9P2xd5iN9qqRhlFAY0U8CCb8OEY
n/1wDzCJP2CMdKdndYJpbNUGXTChIsTKkah82EMAPMk+a3h48auyVuMbEInxIY8nHhFrYiEWQk3Q
vFmEt1+bX9dDpMKKOOdlv36ufqvvapQ54YYwdI4jmqU23+u3+M4AWpp27wMlRXXpLnCTgYFVJ1F9
jAx+mPu+hVQMDpdaxH+a2NBnkXC3SW9pv6vbMOne/wu/xAC16XaGb8vh/rZ/U/elWsWd6GlEKkOr
j9foky93x83vD7FtL2tvcc2i1nk6JWLbqBpU6ryCL0MIX3Ukpwn8l8XUc9amOqMhXRdjK2tDW1xa
S4a0bXtWS8/Qchb2/v/kK7NPL4tS/ZRb9pp5v8vpiZVbHKjO5puLa+EH1mwbudEo6872eQDjsmpR
B91Ix8tCIwp4cQ4NtLfwJjn82ohvpdMiUlNq38OoGUTNXSfwaHqAJToQpbyHZ3nieY/dRZ88truS
22pQyddEV13bJxQJ0VaNPOILzAG13lTOWztA7s/At576Xp0oUa4FWs7n/YMPKEsDRpRTjMT0li04
//WBMPPFXl15L2y9lAZ/zZSGEy5XJz8ZBueRQpRipINWNaxmVKicVXscAEpB1kjDt9mbn11Spbl2
MSWv5masN1IJv4/qvg2nPXhfk+oa0c5YdOWpsjT6gnqJt/l1W46xG+/cmzeBcV0SbBbLYvj6iZRF
eoLhkL3dArKqEWjh9PoDI4+1EkfFUcWbhqa6W00+pMrLyBeOQje8+oZsFc+pbZaah5aGfIC6y4Z1
YHfJgGX4nDjY2IJNqlikKbG0AtHVYygkLAcwqDX6qQO0dHNY/FArILcGs5qZSz6DLDnzFFDrI7A7
P+DpjZJUTXqCWbRSSlWIlNEna+yeOQMl6+rDRnji5bXTfdyrDqHWsy5Q0KE5J1cTvEhAyW03Qxe8
KnB1/xh2NlGMGewappHrooQywnvSSdBbY8Xa5NGZ4AqnqnEM6a24M9tPSADvGx+QMsoCipJFIQFn
ICwF4Powj6vK0V3JRh5v59hfgetpOqwQfIeDUCi/ZFIeD4ituyoav2OYYAA+hPYfiHI6UavhojKy
dHcOTqh5ym+XXbssdiTLNQnSvKXztrdWrKzd73IQFmDlguo9hDfz9mq0VJ3DjQ1EsLs6bqnD4val
o05kO9d8vON8oovfd6lAJkhqghT9a3BRU45IMwvFQ7MJ2QtTQEfyXI2pvWyKfFhwqNdYoARYzT79
+D28c/XMnLYUpII5t1E9tSXkuA/ZZJtz91NJv2QFdHDAJKnWMyRwkTMBDKhZ5x9a2LIKX5Qpp3tT
cDJ5rIHMynUlF5F+Kq9wn/V6MC3xYhmiWAcbznyxusK2aZvC8wYZQV/EOfpsfPj3S364rnrbN/Gi
IcxLnoCFMXewKRppfd0RlCIPni8VaYmAibZa0UhOSu/z6MGLc5sICAQIv7G5rWXVdeRq4rO6QQpm
vfBhxWxX1ZtzypjcJVO2ZfwxhlaKK2LdC+pzj3JXDPgM5aWer/x7iPD6tSdeUYHEiHNDsKlz5LaH
yZw65X08LQfvGmVYF9xvbC3fN1AaY9TIa3NgKBjb59KZQd9D0ph4MTkax3DmU06kJ3STyXjF76QB
nCd2DJbk6YccQdx/b586mG27kO64eT5ltPyAN56N83nXenLdUryqMZ/JGQub1Pl7KRqP0H4ceenA
hnbhfaVNMiiwKhvpJA6vo6NxJeOzV9M1y5DsZheOXYYEYnNdi9Eitr5HLzU7XoHeei3d6tAT/Bks
SNodTC8Xcg9NK2yBU/lfZPA0Vb9m3nFw0GyrhPahfPAi9uy2Vw5UDswFDpNTBcc76KOZ5y37PNgf
ziVb5zd/UwpxDSLPYYCxDqJtxr/BrXgIRM2zvGUs51+QIlo+FrYRZzrXuIKz359fwXrq1W68sGPM
+MLb6wIxnH9lMo7QnWEfkvD2Df22liJPF+Phf7hUqMRWdPEPfR7qSCRo1mYaUEz1UxB1BfiViA0g
nAKB/4tQdEbY6yEvfn1TbGvsiUoGVrTtckDMkrynvA8yrc9CDKYF5N/OKnORIF4Yu118O/IVQoqG
mynjgbImrWniJ6v92kkKil/pMnHnUmevGzzpWE3VXTSj8tigbFKc864FbtbJSYLpIbe9OE3IMVlp
k9vS5dDLrfY6CBIptbDuYwxQMhFfxp0OGV/V4Gm8gy1mraSZQ8m5IlI2xotMHJ1W355VmrCqQhSk
DsZQQFySo5jvETS9p73Sxm3hhPMEb+TXOA6w8rdLBNOnP4b/GG+w4GKjuv4q1Z2KKqOfx1ZOjL94
/p1j8SIOvfm2kBvoXEvPBkiYsgeaukEt4LryXJGqKAWTClygUnktnDVHl5CokPkQohiOyqGbJ3Vp
EYwWPmOFmyIU6RBtE1KrCJT2voDshXgzoN1LJs9jk2J//mhqtLj4pzQMdsX6Dec00bsuMc1ARxAM
iIhpnLjV9OAcQutsYlAzkDWUthqNYeiOkLSQ6AwYmxleCmkrCdruyMbX07L0q+kiOAcG+D2uU84A
WKM/0nwdw29LWgcPcfiymfMIRez1jXknDqdlDRC8pYmPnSwX2CqFQp/RFZJC/SiT5LcWU8/xZb6x
bC3bNTT5dx5GsZAuqjktFXVRiBkYU4pYRym/NciL1afzi27JusHAmrCwHwvYClb4AncyoiIPWbzm
MZ4DAqtuych7m3exqSNCFk8bbuJld5JAnyDpTl8blczfG6CJqifUJu33yEsVmNud7P5jGu2InXM1
KX4U1DGuVQBS3H7Gs5hDvWrPoev3ja77fkA9Y0xPkxljkPAOaUyNqQtHkInJlkCYMs26V5e2I+VS
MMPiYNjSFyCkF3/SP6pYfWt6P+myDDfxqRSc78/+Ww9As+FQDVnDOpKUae7GZ5l6PshdjtC7n+ak
JxS75xo2oEMnqGA7fXbRebbgZGmIcnyEUFn6H8mAqmhIhLpWYeCaz7aZ+hPeplCoXWcL6XN1cUrs
VJcUXbboSouid66A+84Dy2FuTkTqzq+kYzPPK97BndeuLps8uZ4jyGf+015xHrb5UtLWbzXg5Pde
e5ZCpL06ULFiMsetRrXXyWi6TOTQ3VMBTmSeEiZcuCQQlbw+HXghdmwP1AvSqyfy1Mw26Exao1A4
Esrs6ZqjLg3ZXXRSlQMW9fVJZsqjsbcf6zvPHYUEd8xuO7CJ7FCcyyLXXKVLoiICDDWVA1YRGp38
27c+avWy7o92EyEaH+K4cWVJ6yZpzvboNNykzl4wbMHKO6LW3M2yviaY3ncO1STlupbqtH4bQ4ni
nReEQ6A7oj1Ejxqc/7+nFQIhiD5gCmhkEccT3aNmokWt3YGa6eF4mAYD0rzkWEC/CtMP+JY5oDjE
tB5ER5YOdLNsWfzviC9gr4JCaUurEWg0w4oOEldrU7D+kuPZ4v/QpQINQgLKOnbg2XWkmXsOIubN
bZBiOvv4FXZj8qVOLgiozlgp1yBMUBdPxA8MRr92BIGRvmcdyRZTXP+9/h9o1dgLg49eAZk6sQ7O
WsAVAox7h3TudEU7IPdwxUYtUc8RTh7TxlsQU7tXnyPwfYxUeXujaOeMg07Vhf3wB5SGSfvobYIb
9DxawtXyFXRHhPUGdSVaD0c8CPzEl4Dp4puZX3ak1/RJO6GsUH0yWJtJG2cpjC3ExnyM7OE29kP6
lKOomEB+IXnLz9hsF9AB5HUoUm2KxVo8CvPUs9iWbNKg2CM3aJ6dK3vnnsWcBFoXyUuoaBkP0vC9
/gChn78DODDMCP0gSYrJORzldxehTUc1xd+hcCJcWfs/ep/HC8Ymg4/n3PXJCpT4pMNRvo+8Vf4Z
hJixU6LjktpzMFgeTvfulzviaUBFPurmCHYRpqGzO7tbfuqKT1iAJgIxFWbnh2bCPZTGMRshlJmx
uvjrMq93saMCmsHimORMHkfIL8FO2CEXrOEP4d3JLEX984AgxbcP3kj58kabUc/UAOKXxHTt5Rdo
ukljWmc9sxabloIqD1hpVMlcrtT6kCuJC4eFeQDLt+Nbl7RvmT/bjlvNpNQ3fazC8Sszx0WjLf9u
/0gDe5zNb4rv3YOK+7UmiCQemOZN4u9J7kRCjhKBqwUKSwkCBXmpcReRhM2Gdzm9wMnKEdPe2NrG
hm9EmEasaxlC4g7BhzWVwOB3NpvhZwNbpiR2UfOQfaBqiKVtDDAal43z8FFT+wTiZcXxtIJ74w7G
PIt8cNLqBhbOjX5VvYFE7Mu6/jmVqRF5RmMnuyOZJgxVWbhTqN/PZsnDABDYFTzC0JhlGmFnlldD
pOU1gd9cK7c8gB/eWvOos5YalmmUDOFNadxZE+xVkJaPYZDbC8/I0wrIbLYrWNzgiDd9TTYsfYMp
74ej2OHkoFm62RnXY7fOFgVALMaZFhdsLCifObNieBsn3Hba/RGZefqEdCS0fpqBg7mow3vsuqUa
AdrOjcd/WOKHNFGuDurlirql72uoqVDCMNV/w/Hf4nqBUTrdXc24YlnngyaFQx5V8EYUQm/+wEjS
wf+AI04+sCJ/uMOr3LY/q99Xen/X5KF84wX25ruhNmVjjDHE69eAHL3KYCdJwtIc4oJOL8/tnmMZ
lyvqIJ1sQQ8Rs/+PsPNqtKLDR5g4NaT1Fu9Nh3K0ojAd8mDVnIgBBi1+1OUtNxSjbx/YVKianHvB
d9gE1PqxOLPPvlj+t0Ogsfv9CEXZZ47SlsWBSx0G52PKu8w9lUPQx7x8tdu/bebF24tm+5Kz8q4r
zktpamf5NkCsJ2DHzK95tNmQMTfZUwFO1vPSgqbWL+FqT2p4/uhInTaYcaNRmr+pEW2A3mL7Z0gE
Poquuv6eyo8ExS3j2B+FshCd55nbjP0Rkq3WoCKBGMEmhcyzNn6UfuFEjozkYt6nSON5aktqXHVx
C1SmlqpAClL3OpldMH4LhL8sYapr6AR0C7A8jRlMjX1AhtkqIS8KJVhCG50rvmAwfmtvtvyY47Po
kudtFG+yZ8LJcdX9jPGIgtk/2SR1J46E1SVUBxlS8YkPwS5FkwD62c94gP86RxiyIqiwh+WHVaRI
/BunR9Dk8AcYUiFuUNeI+lFEtXMEFGQp4UcHEKO+zjCvgtkZLa6deTeqFoXJtnFUFfqiViXOVOSO
UHl60BcsmN0kDTCUp4TGT35ZvTJapJySMGriA//6czcjAdrUE1kaUHI5AcsIPFmB0iMyFCIGDl6F
6vy7NeZvdBlV6k2ueI0JIrucZfomNHEFOnizU0DfGjmoRqBKj+u399jWs3r2KesIo1yQKa24XsF3
o5lPx4QCoTTWbdl3Z/zI+qdWwmLHoGkxT3azEtB9C9nI6Za29y8hkK5aL4pAo30bmK6q1/9/DDqQ
kAMP6745lHwfW8i3gyPEtxgvZs6J8sNPOoVWUnUtQwIrZR8a/u4PCyzaABQSRfe28QQAYhy76wpt
r4BUO9ZQClUxufienbSuHn+tKhTZvub0bHN1O0+2PlNG4DHTS4bnlnxEPpSL5+Yydbs1FCuCtnZo
ToNtfXoJk1j2Gpf9LcPlyfyRnb9hxNtjYzg/u681oYb8XponbxbMVCviFEffeOVdlaY9naRKF/Rr
2ft0yrvRh8Sw95AE3NVMX18GBGzBYY3DxLrplPKIKaHvD29nBBDT8fvMCxe6jI0a2iMNDml43BkB
gpdMpOFr6GFBclYPkMAYa/5xkUVWXdCrtff1FUhhHbLNSiBXOKx5qtijwmCqWUpWAaAloOz+4nJP
Tm+6Dhk4ugqypZsnxJ3ZJqr9REJAT+s/7ig0EPKkBDbhiiUpJqdU5458wKgBCTtr38cT9LXHGaip
DmDpO8obtvW5qCXnz9opj8K40Grgq2yXuN/5Z9NnPs+Z2Trl/6FpcL0V6I7GV3JcK7yjfT93803e
++3gRmYIYjRdI+67tNkLmkRexUG6rkSSFQqV5YHXKurNlJR1vJ3w3A/jS88kcqIjErbxNO6c9KZX
ieH39DqOZjpEmO1sucu6cy5HtZ1/IFHRw2mY6fqbD/BX04/MscWgERYyNSNdLUIIOBF8qq50cWIK
nwKT1EJ4Xfv5T9KMLUStvze0pkpwUmmmNTa72XXA1YgjpuBCAXCRYGll6h82PINmIMK2mzJeKJSe
WtZxOOHwo12AumOx27iBpvNthgCNcdyTkbUUkddKZEvC9k3Rfd0ym+GfSNySfhvjsmbLsuUyQNFf
vGmRPKLtFASyntF/OMtG3T10GRietvtqPY4lOC2ZDhV1sb3sqmKCXisQBWdtdXrAOr1F1GfyK2fx
ZJIIP+3iElP1U3YfJOyDDkLoaAsCsXDE+GIg5XI2HiOPlUIPYoh3Yaq08UrdbN23DI+ZKvn78Q8Y
IYUWkzqd9F7GiJVOdmWTXTr4eqQoQbOpN1wLTf5lXriuvdl8qDZlGDTMCXl1stRc5ZQhLlcFq1FY
O8a2nBTjIlL3FGsSMOp+F92lPfftvpcI+H5rEuS3yh4dw/yiwP8nqYywBBVsLqNTI3+elJ3IjKdl
dbWTSQ3K2CTBcB8IBtyH7tqzfYMboxtj1DiKW/R3oKUjn8Xa0hm/r1jtGeZit3Aekx/oF7f1hxPL
lMKOgwLNP3asvZeu8KRn5c+8EiDevw1U3Shr1U5P7pj+e2HEVOfpw6hrVXM21K9B/GNBR6iawzx5
LHZQaOXfs/zpGMXIENYrEWtP9bw/l0tgLmTu3KcUP/JctZvoRfqrXQXGyt7Q0bdTWLXrC2weHLnD
SvWQbKLHY27pkDupD6vDklh+Y+ECcSoyj8P6lEcGDUmQJMKOCpRJg6fg6daBKxcy9dNfbYLvciul
FKQUHXv08J4Md9NV5Nc2rmRR6r7z7X4Ww9t1HJC09s5hPuhq6uFzKbzCtZ5/j8uLSSXrgfDQJTud
k96FpU1DzyS95oL3VtuUdKoutUhykJXWYpfJCNrH9eOy78lAS9apLbpo/9m4QKwq6avySy7m+z91
Gjws+HzA1FKHzvpjHSnJhf7vce+GEIBGstvOLhRwRmqrH+QVcPfiB9+GnOo3+C4yoQ7B7ISDw8Gz
784pPXSOhFW4NER0w9eHJPl4cduK254722jFu/xRdFYzrSPKSgMSXNnmLfsNJY4jFOuujK9MnQJ2
zhwkOsvN7bqDjdoatQTl9taaXXCBi/uGnACAWN43MYzS9uMRP3y5h+I88ULR4i3zOh2J4DS52lIu
ZxBXVjWazAl/ToX6PxYN75m2NWOTDDj5ouPk8YfdHSgYSmzS0hfj6I4WdUXW7vaWsXWXKYDPXcf5
hZWoS53BR9eZdcRSuqzANE4jsR+zdglJ0PgeCa6FChuQD4XikDCGJ4HL/VTvgn1Me4WbyYsnDPb5
eIHoYQONi2+uxjIbZvf+JdMAe6X3NPMwf9cWydeRvjN3JWEVaVeRpxw2GSCwd8ZO3pv0ieuuLwCp
ogI7TRao60gl0+qnq4ZX5u3WyDNMfaKw8PQaIhpoyw/uT8uHQ2QoA10ghfBP4E6R8gyykCZbvM+x
Cg+NTjdJm/TqTxcFECgrETUcQSpDpHppQrwJb5Pr7T1eXi1VGwbC0jZI9NefXTDe5/Nr5SFCbgyZ
qJAJQEW8SaC2JXUPx7Fcl3FMBa+bM5yasAubSjNM8I1awJtASwVAQNrlfIiAeFqjHG/gLLtRm2S1
wFxxEP+n/2cuAEwVfKc9CXvlcLDbzgUXLiPpVKiZlpVMUwp0KscXKMGzoz7OhP1v5xcmynYyWElI
q27tpj7cAuCWQpfo7isxmEi3v3B48nAtAWseMhi4x7q0xN8e73xsT92pnfqzOx+85rx+OSksCMLv
dpJa2Q0UpCXvNr3dQEYGfe3RJ3xwxeh6Lsf7MwsbuM7f+83FAIIzTjqv2m2Xrofp16Wc7vw0eS8u
TdMmZ83DcUQ4+S2PGUUImonuRT3DBcVDNQ4VXFbP+MD+T1uUNmrnIb5ZbQqBoMRl5ToaZ2pbo5H+
NkrQdzxpVkPI0IqHPG1aBMcvN5jCR5qmYjq5Zc9wNUoM5zg93Eti8TswaqghyyKh1j12Y/Jlz/AT
XLTdKOhkhqCVZWACZ8v0q3QvW04btzhHZ8m4hhZtRuzuzI8ki5/5mzE+XppOtkL+wazEgHQUwH48
PIEQqUfjV1GPyfwp7EFlRxAwNrmep54tk6/7Lz00SqRHJ7KaMdCBdVZ5caZeCIA8R85LRB4aHRY3
ioMxrB99ZEyUmGonVHoXQTGbfTxaIwdH9eML9geMtlBPy8Mv9dT+HbrX4S9qW/sAedUDHr1Ve6JM
Onn68r/80CmniCbIIZtnCoCiVqx1vT/qcAw/ZZ2BqyobMP77safDohTA5OyWdAWFfT/e03gFchZk
DSY5RcujHDZw81n6k9M5qiEleK7ZB+LicJ1xr4u3v4Tzq3DLm+chQ3ScZEIM0XPPylQ4Th7dfw7A
vhswzdlce0Po9Ean0++DJpmGApKO92Cs3hCSxzVUkbzGhkknQVPxXCAFtvAlP916c2ib9AQZiWyG
1N0gXjaSmm9cjIWnxeuYFDZqh8adbfVyrlNCVqa8srP4bvnansWmfSnJMrjRmSCQe0Jcr1DmlIHl
aIdtG5+nvePF4B/msum18UBo2uUaVOrpuYUa6KgyeNP4aegGRT5uy8lHMijNsNkc49UeQrHC4hnv
pYgbY1lubTG8e9X59gZ2mcYn+9qw6HFGNf9Eokvj+TaVqzP1KxcVoWb/Mld/QR3dFbLf4mO1i1pN
LXTMZWM/wmsdNB7iCe2cfJcCFThymR0keOgLDHn+weQtxKmKQkqDm82Afc6iPkFkpMEQKb3Oxn+a
kFyRLqsKTPlQs3uCHOXE7Yaz7Mj16KzqFUvTTj1GsvO96JJ+ZGDbSzFrSdE8Q4t5+uJ7/CnbaQSG
5UuGKLtolXO0C8O/pqXLzYY8aSTP9Du8IJ0GIKTHDocooIiU1/IslIRGKR5ymfKEiVzSSqQ36Sx+
J/vC/+7AnCVIi1kWKOzRXNNSOhx4l5JSXJ6oytTnKiTT13Gn2i64+F9YoOLN9ngLLIfBYvZy/J5w
2I2L4AZPDVrAZV1W5BMMT4aSLlMbWB/mMOOB5FHz8KMUVKt3DJ50DAPIcvTVv49X5tDqcqk5Bzsw
fiGvjXpbhCiMXfUraprrs4Ni/PThsybg7aaGLdoAotK5kiikku8Lg2akVk0KBS5sOp+bUw74qgHn
rfPDvr/TpiFJWKBp5GM35cn9phTAwPNLQnd664OC7JnipPwbqtJkm+1ftQNV4JJN9+Rhl1RQnuY0
35V4EExizp/N4bpCUzQxrpjMKjt7zzlgTfu1yNThVNQ4Dg/xaFav/FaQ9AYBLkkU+/YE/PLcAAbP
K1z3f7n0bYPdEzCZfZNjX/Ige9XiXTljc1ss98OSHYyTPBr7FTWBuJALMOK2EoE81c/B3EPAYndY
lsijrItOX9C0/IlvQGiXd7hFdOyFhigrLIqqUYWI98hMvfdpCaDxZyAoOCa7ZhwweayGDQbkFBVY
a3U3eB3HGocORx9fSrcAoekU2fOjcaLz+bI0jjzYqaWS/0TQwvSJv06tR+arzo22SADtEl2EPEcT
mRGyBVtQny719Tn+6HDERDx67yPZyP9eqGAAcqzjoC5nT5UrwQV2XaOFDKgh9Ax7fvsCQfIP04BR
nTzHCy2PYbVHbcPBg3HVOPyeWF/Ni1V2xpLUxlIsdW7MIHXFA/Q5SM5ikpTnN7wJVmlacuj481Kr
SDn80TYGOHgSGNQ0ysbIc2FxjxikdxyEHvOCODndDG+3lzQk3r9Vo+C/RZO1le0kiL/5NeBxcVKV
d8BtyX5BDY8PWHzlFfhyTJ/vn0ys5LAvrOhufsfv0xzjJ/HFNKQruD+W5eGuM9FYLU75NWqU87Wh
YK6+InX4q3Lxhhk/Fl5/9sCxwzIvJWgONyJ+8Jix4Yu8/uK70VZtAFTv83gCClFraF007vyf1beX
duJ2U8V0pKdNShnMbryLqM5Y4KFlQ03L8FM2oJ9QtBhR0QUaq6ePA3nlC4y3d0trJNRYPc7f/ZoP
nDgPf0o10oK+YVpxStSWQOm8QkyvzWizi3DWVessunmyXDPtU0tJYFSBSRVY1UyCD/E/Ra6mspcV
3nj15H5BXSuA/6IIE9YyrBqQ9MuhhKXH0OwT9rOhe0+rtS3MKi93jl0CLP7au0N2etje4ahCGSYN
A1kzrJayUWfJFoXTgpGO1QNVG2FVEF8FSDd4kQiDJrv3dLCsDrsPH3Hyx9+CzjoeZG54+BXkZbrJ
7pB66fZYz2AAmRZ09ApIckiEgWNu3I/NVp0J2QGp8ku32KWjc4qRObbMBEs6/C3nWVZobtqnBZuw
lOXPpZYglLFPkmYWHimDlJAN8knr8m+8YWM8fIrpQmn+c4ND9KPFYlbbCImmErmVcNz5dqJRjMrk
AdMnt/jPf7NDQUAMDhdqWNoDkAN8wVSTo4yAIhJSyx0S8nSwirDmfS30A3Auj04pYsGCd+8wHfvF
4h9OS+dja/t+IiatmfaE0nyDkQttWF7kwrf4mnGF+Vr827brHN2VhUlv0yyutllhg56FM1olnQau
Lj1ac9aDVBUfvLyu5yp3wqHBzT7+4r1LJy0q45VN+mB9L7oNEuxerewsCM3mApvBoz3bGzUwbIVr
ol6JtX7ccQZxJmXyqvYXOFZAAji8n2fGfguryMCFDH4THpocjFMPp9P2BFmFmJpcqs61WZkrbeNv
xslBQBUYf01vHkS3+1SxlG9hiIs8uGfiyco3g4KtRI98CuBp0k0zt8N/BKsM4RumV/81j8qzcQMa
5d7oUtfxc/UHr3Dp7CvPsr6NzwVZN19oPiYq1AdEbZaNqcMyPPThIwFUC6hdYmaNKGS2UHxW5WW+
xpI6utgqkhFif2bPWnDF7PNL8qr7792bmYBujgcRgwgowknQUCec9iR3HRY7Bl2u7PH/PyePR/dX
CuG8yG28N+nzUCDsUUeBojQWFW24KwBKlRm2v6ZKibXgFLktK9NrSs7GKPqGQImxePdB0sSvi8UT
YQRPX2QUfWjqiqpVhlosiKjwUMKdq+GfoeaMVyOqHSxi4dYLJN0DSdM7ozyfX5cBCvXyQ2FCXXyJ
cUiFrlsC7SSZ+8bZs8Y9XLo66CntQ2PYeryeG5WXQKm/TgUk6nAheftABS1MjElu5q3FDh6hTic7
Ymx2rhYNmCPt5oIJWu88bJie/Txxp57ElTgkom7SeKClKCX18FOpOTrV86WaM9yk8aruDvaSJHZA
EmAdlYZPFRMuShRlrws6TkdCrYKjKQHcIowf8QnsX8a9keqGMtSh4CeSj7ACZEhG456+YlUIWAyT
Mn63ZZLyHB601ex5RnOg71JzMw/hNf2ltDcGiLNsAyhdhOB08zBDvgM9lnAPkf1gWhJoJyPa5QS7
miGsDkEJARE13J9RsbR3rJz/mCLedMTSuNkORuAiGARM4+sp4wLikwAiluqM6msiQLu7JCHCxXCE
qJDCGaia5DSSiinU8gI1aKdwNDCOUZM0wqsuXVzhgU36WhzmmWwcT810SCuuLBQlwoXBMWxxl1AA
3zlgXOBR9wyr3LCFA9s1W2EL+YQ2CMpiD6pikHCR9OLNBEEWE/xMz8tGl2w5W+Oif+4vaBnZauTd
df2xXSzZkLk2NH0M/Sv5rrjyagNDy1xLVNtV9OmRUuMNzh5LyXRvxT1bXE9BoFxgb3kLWF8I30X4
IIbASCMYPPrg10zC9tkL1kh5OmT2v5JICCtsDsLklkt9nvoFIdl/Sdv81X9evwF2kOSaUEYliIWJ
HZ7Jzt49XR037031ndEJvd8xilGY/cuGAuHSo+1rFTepD6CGNhiiGj0QQ01e80eU2PWXl03ihx9L
E/q65M+3c1eqPh0AYaPmYG1v8GC/1xz4QTHGaFvN3ZDSxJ+dFT2tH0RXHnhNLPtwrfJgOLoXI6tA
AGOwj1+Mt4anUMjHhgMBEsEwFanRyV8/80Tb1Pxrps7atMhbF/AS5ULdDyznBMIKsRmY73Q2ALll
rtV+thq2f0VOpnkfdHfG1kiXoS8j+mYQxR8ZcpUL2JxOEg+Lt17AQJhed3E+Z953Idkb34bmFH3M
4l06zp+YXJ8URKeuP2QUgmc9zlejLUpqqVLb4Ily7NVbej2+Uhb12DkJYiK+kQIU9A4BpT+vuM3j
ducP9BVIvl+Ta2mMTM9s7kWqDlizjnEUWUkkuiFNrzwk1kZza/PMXPwXpfbjqV9YfqLY1FjDWTl/
2X0jjHU6fT+BuJuqkC3vCbGppdC770n9DPR2KC6McYsCsPNxwOj86DDLT52Hkxr/kEPmaLUv/TZV
UQrPcmybIybeZDhPS4pVH6FWEHwIPBs8/nNhXORSyjnSyI1WK/1m5e5Dkk42TWGxaIz1qZ6pjvab
n306KwPSJ/GJY5IpXV9dHIX94ZV5t89iNieqQa+vN/VurvGxwmdWs34SJ0vTq7mlCluQ+jZeXsOE
3f2+Fym6l9CtDgXMmllHzWqTCAKVL2Ux2OP1wAuL4OvqPQsk4C5Z5hodC6RzZVSgTwLtOhe+7cct
C49xV9SVeZELTJmmGbO6iIUC34cKLTxWjmUMLK3B0dt7Axg6lQISH6piE6r8SvPGqyrDxX9QxMzj
woxvXNcbOYqwlLgIXOkVh55bXwFq68WA4NgS22INrnJa4XfA0BSFWm91VrWvumdlao+hVH/V+Vpq
l7Z/ucE7anGBL5ZIwo+MFxEk3Z4XdPBZgmAF3cRh7Bqn1hSMC+cqztu8Co54cVfV8puHkVCwphbe
TfkwKrD1AWyHHMG0gcTAsx51vor65nOMt1qIqpd/cArMIcvctS01aW7GuvkDW6RcT5+s7bBJZQKV
b6Mq1DwzZou6hUij2QIukhCE+l+6ZsETvALD5eT3NN6BUsOUN3jgkQgEkr32dBvNNT+IF23RWTmR
j6T4LAuPikfed+5/vhxKdzBe9cCe7JY1HvnQZWPCUFLTeM320YsyyphTsjf1mP0m2Wghlzz5O2oa
dkrdXIHGm8dfbRf/JY8S96zV2XhUXHeG7sKeAaq568QCY9/J/wTphZP09yusf/koRPahUusBiLM9
g3MjBxwXT3y+MLiJB4agSErbq+hWjoXpSzLh0w3H3l8jxn+WZbfTF5abz1sSrShZ6sTIsDOs76jd
MJeC+Cx9ZfcV7fQ3vI8CPnjehZv5dLYABd59isYi3HiW3cacwbxBOnXnecCmQq/LzIdWqF/Xgxrn
qoq5SdFrGJbVjgKiFSN86CPAiDvpKvWvgzky3XMaHmuk1Gyb5D5kOWRtN48k/AVU+bTOLpIgNv4u
UTU8OSVVbK99loWvWQsBUkN8R18N3FsqaiUQnz3+/Y4CyliLS7/Fiwa1ZoB4MP2xFvi8/4VG9wCo
2i2rBE/ZCNyH8cFslpyvgKUE+MZM+7Jw7vv+ucqeW9Of7qZLUbSKifxuzbKQBZNhp2Vjc47pagtg
h4JSpNHlju64LjY970YUeMv40t42viZee/x+JzjcGLgszUY7GC1ktGxtPQO8J9qklcU+mDX59aRs
1XDp+1PP/u2L8B9FlUmEwDaCYDmilAQQXuwf8K8pErPbNSuvHecMdO/wjQvn7NSLQd+qgr/uzQJG
wagO4UVyLzlz8p1BjNCdLO5vW36cVwcqh9w3pAHiqg38JlYtVBPVy46orLo1JI/uDsT1kN+ZY0og
FhnnrUBPpDFqYK6HJ5KbACxu2JPndiP1nD4gRwahrBhkP0r1WzU7faed5N0+8ae9FR7z7E0O2gs7
aQE7AYtUBUSiqRJS/qMAAxGceePispufg8UESeQnrn0IzJyGoqS/eLwZost1wfYK5yW1Z4WvgIbw
H8G0XUCqbioFhiCYQkTranVt9S5a0f7qcudPJnO8UggZ0wLx+MrvaBGMlkG50BT6f9TUTPZgDaRw
aJnGmBpf7R/tVMxXDZiWxIo/IshyO3pVUvBoUIhuY5bU4g194ZWq6/WPcy/tBt16pX6AqKx9AYYq
xT5tycn21Z3PAxpBBYONuRBBj87mtJKWjkGnq89dmDFMoR8YlzMqa7gq7XgT13krnFJhq45LT2qO
lk3mvolcIVaqmtA/74lpQtiMdAJNK+9y+Gxr+NaH/9nOMDbGyW+EOEhY2BFpRgYb9RyvBAorNNdt
b6MsiM6QjwLJzwleM8QMrGn4tCal0WMVDo+fesnaekHpRfWyZUgkm4Uhuvin3xfU5ITs4RnrqhcU
KRu2tuxfH5UMIJv29MFa8mWfzzKBC57HnL63pa1VmImb9lAtBGvwfsgs7MAX2PVbKTF2jZYL855P
fRnDKoeQ5nng9pFCCqWdPDrHVDy1Augk5ZsaDVX2wkZRy6lUqFrQM0LTw7PcKfrAifbCr/x9lfr9
qidZm37PJpgad5ENrTchW7xpsK2//2RWiiNCUesFTQEcb8hcyeVPfqJlhc6dTTStfzaPC0GwJQYH
zU2JIq5l5+5Eszfr0nWb+LgeuWUsOhkSbZe6Gr5ongJ+VFDR8VmcAVSOWVfjmuxJfjN/o8CeOdds
ahD2Cwm0VuzkKzSAjQmxgRlq8T9H5q8jKQrT78VpBuugox5dsiSjbUUkCiIPvmOTZWj1HPVbdQfo
hlBjucwRg74evngRUR+h0aS8ZkqwFVia5Z+Z/I9UUcHrv1kXyGsgiqqRiuZSLx3yVDPX0sq8hHXe
cEtJ3Q+1vqKHstYZZWLqAaQzTsvByN9i6NNRHGcsn/1yCl4y6KLX+EGmzEWMw/oMe3/pu7AjSukN
4pOegFXf0I36CHnk7HFKsLlDJ3G0Tj1IoWBfHqZLxN3q1ZnEZU1cuqPWyDkMM5WT0/ukky3WN15G
lpha9nVBOFgWWsSoRWN2ex6a1PxEye2fIzVStt54j5Dl11/GxAVXm75NP8Y2Wu4AmIrs9qMwPpaG
9164pgiN55sYb5LAKWoiRPAEaFBGDIYMa6uiJd5kIDLyUoN76arDAX6cb0EpOcWwRp/SmpWBBBur
dnvkDUdMiABZZl8NHwQ0694hVVFAJ2Vi80N/WFOPXlupOqVCwoGmonsSE2IBRR4GI6YMlKMZHJ7M
YqNTdDPWmuWio/J09xNDyeA1YgGne9DupyDRq1MzuMl6A//fwZcvV+0mzj8GuMpQeZZYnHFg3KLJ
aRdkQkNxp6LW3E38u0VLYFUU1jGrWrcsI1z85ZMyIe5laMB9kda4z9r7ctQVpDa60zRTo7CH3l3K
Nl+nAhGCfh+TfZaFleryYv90ebDndF+rksKfayNsjJqq8FrSAcUmUbW4LBND9ajFgek36gHRfynl
1vhxRi2vC745yIKmeTVuE5BVaSCqx8yHANPCcrcGbPI/OcR4jnsHvS7QoBkixbp4OGlCpjnlSR9p
FtCbJrL+SPjKr1OE52PEzHTkxKxgfRpEt5KxUPEp0cn2ocmybuA4UUfV+cnzhWIPy/msH74ENpTd
DykXgM2jr6soUDVyd01wT7bwupCi/sHgrPRYjwN/FoAaLF2u70qOnHjlMOoNwWD/d/1x03s1RE/U
O7vTsbQlFAo0gtvk1giDSMLWLH6Mq8+Z0KdtVxdJ8pfN41xcyhWYU1igHHkGV0BgmX2ImsbI6gVx
qeFebcsJBcrIsxNP2/yBL2gkGMnoOZsurF0JAzW4jcEwSVLPReElx0tgCRYXzrzB6n5NzQaz0QcO
js2eZwJPB+NZaFcO3Mtcok1Ph6OApHqD41eH3QzdihFfAHAtRkETEiAjHxpTTuYMPJ/0lEwfe65X
byLMIzibnaKQIsha7Yub8Y+AVsjdl3Q0JGT9vnxUWIOtdj95h/qL0ryLi/gKc3nfHQVDHio919Mx
cGtij3O8I8H0JKiGoETKyDPtFVpLZs9IhPDQzFRLIyeaY5JFh3R1bGfiIbdVyJ0W8cGYi36mur1M
jANrBO6CKicfgZ4Hl9mzzqhlIg7ig4+4GgTa5X3NcUP6Fwf+65BqoqoidchsIjGK66mg2MxBvDEM
8lplNIe7vmyOjxIoxXXg/wu2lOGZundmuaSjXWllnXEvVH8M0+laMlQmcnWdp1NCkDIfpkDugUap
UnlXLxaQvq/Kju8sWxLzheCWm2aaOh4h+T0ubxypHpZafHw1zByt4f9XqH9IrM1x33dyBJ70JTdb
k4Sw18Lc48h+4DFqRhY2Z/Ma21TuW7SSOu2kjtXCy2lXLhZWJhvls1l4j7g3rMUebojL+YhcUje3
ougdApsQRXOkAIvR9N5fUqrqyDrR6PtQv48PVpWJdQnzPNW+BUUvWIqDEUiNaleqdl/fzkBpZHZG
7A/N73UzJTygHTVlXOXvckPAZpZc8+9gmAx4cHa0QRgLXEd9XKNvSOliOhzdy2huOcMNYU5cUXJ6
U4YVpxC9QaRRdyr9kB5qoDpm4W4SJP0I8x9OmRZ3o7ZnzLzr3XlcpH3xITdQn9terpCURFPeQU8f
cHFgZ/ebx/GlO1M8MMHGdjw4S6y6OISpCEr2PXvUJw2TqB+Zwf85eoW9Fib53ULOX28JoYLC1v5l
ZRXWE76xVSFhY75iuU4y0eEW9xNLjdMla4vgB7ZHaiY9ypHVssisWpNmKZoa+jkwdXQID5dYPyme
bopaFoDtJb/9q7rWhKprzp24k/aP/i6UaHKVY24sApALHXqJYb5WAIcOatQatQ9oYN2b6hqqGMAY
R/sxLGYjw/cjNynzNsGtO7F/oO+zd2QDd0V9o09FElA8JgMgUXSUT6lZJZWn90XV7q8QKvDmlHUY
JwtToI9vpE374cZ0jk0vVKKKYpLERg8TFt/JkPUqjxGoph4PB9QM4vQ7ewV+mbGexCGcv5emXZDZ
iaH6In9MHlZdP2OA5zxRr58+q7ybpdDM2O63guocHjyZTl6xVjFK5LBJ0Q6wW89UHIheAl0y82EY
yB3miTkDCvMHTDi4G+ggeMlGI1a/UvOscx0M5tcdtrP+OCAb9xx2beQf/rakewEmfxy8y8GeMyA0
uqKPoG+MpCztsWRRBSBEWBvp8pKCTUdC0kLD8yyHt4xhpw+z4XJQGIcVwX8V/yl8wcs82h8mH206
zN3YCGo0w8wBXFAtRAwRC4ZDBctfxl1kvk5GUwKXrL04VQTsQ3TnZwEBItHV+DddGn11PY8CFE+M
B2eRE+MI2zNhHylrp9UEyhe/JMER8DcyKchnZjMsYNGPogIjMNnC0CZ/HCFFMnPPkk0a54mdHE3D
w78jlzt2ceaa7/e7ABdznwvbBLsr/DTaXnIFIIMNrKnFXDwvNnpQ5O1VDhX1iLD5iSwzFBGdfwA/
6wU6ZWv/LlWGxgW7nuZZ4t58PeRvUKjennrkFBF/IQrpMJgvz88OPnjW/4Cww04OsWlA9KWh0RR2
yEPB7l1LMW+hHnfSeTlKm7loEtkxQY74KzX57up9QD4KiM9KkZo6Vocaz5CWLGOHy0IvcZa9pjug
u/T78Wr6EZjKVPE/Y/60vBp6n55j8EHtV8mAaD5OWEpjpxJaZxxqVv39ulpJq8CKiDzOz0Z/VcXa
c/0UwOBSpgetfJydT/IkljWyKvJvmC6q2vno6HNRLfcbTnbIRwc1ZdxZrZu6fum0zqcgKU9K8HU5
g9bovL5IgAPtcNLP/PXk/dvByZFcA2edJK/KgaNnH5aDp77Ap7LmJpDsCnUyIa71oUCDdsp3UQtf
GjW7wQye8hOAdPogRHLqD4ssRCtFcg2B8xum3SdB523AcbhlkMzEAvgWXY5BzE/E3HIe7NWyKuyl
6jd6NisOiNKOMP3fD5s0gNtP1D7SwhoqNLJpNAJM4K1wvQP4naVo2P91RK7mf4xmM1czS+uw/Ur3
eHHEEq9wJ12m+CkxFc+UU432FOCiBTQ/CESvD/gxxu8SFUoCyZR5w0DnBFCUlYLKcm2esfPAIqzC
ZJYTmvU7ZGUFMJa1Xz1C1eP6qpIBstzK1+USbmm4dcvVtV/08pwGNF9Lpmgj9uVPsXoCQKFDG8wC
P+Z0DTY/OeKvN77Ipk9amDnA5FCnonBwiryirT7cRrgGw2SE3CHpKz1lAR/+RCZaMS+Ovvv1PJU8
ih4UdFqqY8RQYeNvGclf27BcKOf/nNfSFzyHOSp6gOLA/Ooo5InS2S4KBvGfcce6TjWSQEl+GHSm
lvK7uPNJbR+mzzlOt/AYtbdt4GQ4SQVz4ENhIYxKbw9LnQtyowpe+OGwTSSudSPIBgIHT8MWxLmf
Ng0GUzWk1E/EdJerb0qb0mvkTPrT1EWH2PQkKQBbfFYeMRC5Y+v/qOrF0GwErfR7/bm1yr3acHbS
QJ3Xqb+eyrdkjPlIX7A7GxoAZYfBlOXcEStnjLgKAlfDEGSWxqsQyLHSAiXEsp+OGEV+wC3fvvTz
ny0w9Fx/UJ1W0y4RJfeWmEexZKwK74WYuXWmr2qsYhcHcAtEuZEbAP6obsSjLUoxYSMXHcdEOqgB
hbfltxyNtjSXeKhcznqqM+HI6+sWQ1e6sVwimvR5+fZ4ZFxmHlDKxeLaVPaZ8xJ0vJjLTQJ3rSiU
PY8XGClavft3UAiIicXvH4i5T2UmfdRXxy45SxEK4nPVSd3XvTzBK5t3HMfo8Dy5zGWiBN7D1eDs
235IrKbI9FhBl/gXnAUtr+xZO427nCqzvoK0USmPBj38G67J4v3uKeK4ozTz44cALB1JYfnuhI4o
YWuMtvTd7QU829T3spos++2EZ9vOHZkQbEu1NLE+0A65BJgLFnjZU3VsmQLHqg95y0LArjB8UY6T
oi5t1nSCJAqAJSBOllQleA8nubLi2pDQfP925bF7/3IOzOw0TMoLibhkKT5HL6MUW8hzNqWCnSnn
BGi9Ko8io5+eUTLC71Z7irhDmqaAhSwlA0XhVUaPv8+TqHbPtSDx8mRKvogxZG34ju+kGnZC8SzV
KQxNh0KPn278FV1rFMcXog7f/zdzt7e4J0pvfPIOND7xiXd1SswF994YlQDb6PG9HnKoke6nAzVy
appSnzW/13lfDx2iWZRA64H4KECyGZXMklGQAqBrLRwYihQArGfxfcGvGdSE6sGCWYk97WxjG68i
sP5i3HReKTnkI9wnoCJbOT6Fz2TjVOtChUIdHuUUYbbcye4vGskzY3Ov9js3ErpOY68MuYSu75rq
nGeC7jy7dbVJjTMvcarb2mEGe0OMDssrbBrVWUiABvZinTthH3e+PkrSphTRywHjBa9y235XkCJc
Kcch40KFvPmDH7VFOxZNlbyRSsAJcfJM6jqxcnZwv0zR5t5vJoRXURy6MAmH6QWJDjWAGAIF9piZ
shJ4dkpqnTQ5TIUZvpBcyWTMmub7jdxqhk3V/zCBmId8YvzVzpFO1/19NlkP7Cw4MEEIlgZzxg9q
bHQjhTuDTojSAigSpQMSHfwnWjtALMLruhlnbLcL+X1PKpeFeFbvLQpgAcEhPhy9PWJ3S1bDeNPK
pnLQQ+X2XRbvn5j5MQfTMt1itN7hm6xauS8NX4zvlVdfcci0nJe0Uz9p4TM0okbTA1Juo5eRj3Ul
nhZT+wq+ZVRnthnelpIRKoMdv950j7as3Fp1Mgd+0iGSxSxzp08WXIWObZ1BXNEtmxm5zdEhKo1l
u7QLFr842/k5BsSPlVJdjQHrzxMGrFjMJEqphT7wiZ9aw5b8FM/S763KgAgR5q3iRD08corgVwts
6y7AGw+059nWfN2h9AXuvfrDGyEW+0om3UEFUISZyHuR6ZMacT53fJJt5MbK5okHmEEck9zpKwGF
8K602bTri0jf5AS+fU6WKo1zPR7mxjBqlAdTAX60dmAn21iMCTZPGKzjQ6DHX/oUESp19nLZkP2L
1oFiYHHJ223PGSGIkYheAI4IyYrLqdVpK4cOKBlVEWMTXH5trNNpwcMY+2t7k2Es2m7PTHeUWM/I
5182/9G15dNwSId76pqCuTy+gjmccAsGsHlkDKvJzZyOgmqpRHG9wMTWRt0T174wOHn9vLBkOM84
JDJcPqQ4cmRhg4M1hdWgvYZp34F/gE+mM7R1sDnV7fTW94245Evil8O4qxChosHijgw2K2c65lva
7Pw3hLl7AoczrK+pIuVBbj3hmtQYjkCKINbm4bPqW2hnoixad2+KU3dIhBtvleKxum37Jntp6+jD
CKQ5hfBXJRRL0olqFHKpdUW3+FUyHMSqDANHFi5podKnY+nBEK+fM5Itc7izAn5UqgT1j/1yztva
XAgRPAj+nKQBOiMG/ZUwVQF/F2O7TWaFT90z211zjEXy/UUbs6bWSP5gHvTHuq6RUt/dIdQY/VlA
d2rbsJLDCPxMRvoUzrL2l23T0GO1o9dHMdh/sxrtqZwTIiuDkB/X3vBMRZTV55rplR84k4xqFIPt
Q+55lBOg1ASeR/iyrk1CuGlxmuQcMDHS0aga4nL461DukpOqFo8EiL3j26AFydLXXOCFNeX5Yo5v
kyRRTJaGEIcpD+QyThFV0dwu380HWoBM5PLIEHgvkWBH6TLzceGOZSqgOTg9wcW5Sbhcaex7Uycu
1mXffdekBBYflqJWuM8YswsoUdsY4WT1Ah0v2qlaswYvh/Qu/dXfsLR4A5cYHMd4elODlgIuuYh0
OzC8fj2VqR0iShOEtTedU6HKVu1mA1uRD4DLpqZ09QqPwcjaHPjnZchKCQKmVr6hnaKeJBVKiT6N
H+fR298Xu9zd/nIOMfqF8eGc96+Ua4ZiCT4Uvo6uvPQOPu5zBXqZzq4FlWBM1LxAi2RvU9FGUqHu
P5CFHToCepCtyALwXkw+6Rgd9Dqth24IM1wpC8fA1ZirhQaS9tMCN5FPOcr5rROxgIE8pm4VruyL
ssxCzsBTewEOsE6icod8PvoXTGkdFo45gGUKSGBQJobUPapblUz9yUaZl8JB2rdtHs8i0vjgE3C8
6qsAt8i4JVOHF5/Grg4hQg/VQiFa5q5lKQuqaBj74h6FWN2LgUB4Mq+hXmCJ3qloW9BgW6Sb4Unz
+1RaC4oY1rlu/3jBXQvF7LFZEtP1rUs4LZy6WpgfAFEDzhkiF6eSC4VY25Hpt8yYO/NTVZeHxvCp
elxE1FX2BtqjTwfr5CWHnt24vQNbv2MNS1mhFmoqWwc+fkna70PdFtGlp2Gm0VfrBG+SaqD3xaad
hzqxJKN/y3bo0MBpcrW/c5+FEF8+cJSl15d+g6ZUI1ilvUJCwqWexzOiTifHVAEN/tT/scpV3oUk
mNAarvAqUDGj/0uWIbQAQAHYfEjLweRUUHEl2TqixUuB8El35jE9WY05cxMXY+f3rt2cftZwT2YF
J6r7kZegdiu3aD/3ptGU9JkpGuft0uc0CB1iLF7eRQ/doPpiPDW9QZToNUjj50xA4A11+HXSE89l
6rHW5QH0+1bb1LdKNFKyxOO4r3WOr3W7ylzH39C6yEwkJniyotBWMKO/9T6cJ3Q7WciHZFy49y/J
XXMYE5m7L1/4UcNaywIcvRrdjOlrtJrN6jjrlUejb2AdK09hZOwY8M90ithecNINiGyP/JWwU86o
q5hB+mO4wCulU2caaGGVusLBaJxrFEFXWErjv11h9xb11w8M6w4+JB0l+DdDO5C6ZuuaoGCjvxoy
sghFRW0FUeWJNfo7qDJwLub99N1Z1dnh4sL1kwXvm5xzkxWW5ujxiCgD7XQksIMh6ojxFb8ttHES
DOD9KCeGyyoUX9a3KvF2shL0T7xgxVwnf83W9Pmtb3S1mqFaG5xycn5rK0qMl6TpJJpaIyX2+Ty3
/Ssza5Lp8U2PFO8dZRQVryTHY7YmbTaSiv8EusXmeqFoEAOgfxJxCIlT0lSlbyogvcUImISYbPLW
UG15PZOfoi/HBjtZx5zDGKYCJyKYrIAgo9p3nIQ/dZdBjZbM8x6z1ANlhdv48JYZ7zdM58XEssHx
oUxJqF1HIkYO10ILR81cyqlGan687PBYsLKn36U1tji54GnjGUHJYoOa5rt6yWFXyUtwwee6KzGQ
1UDtEE+gsP04Et2CB89gJ6KVe9SGI43AtLGvVyZP7jJvkXIzF3DNoyyJwv/Yesr//toipw1U+XO2
kG0hYe+hrPeK8s57hLDwTcFqYwoebagzoQmau3/CHwlRyBkgBVSwhI1AAMulCCMg1n7q6jMvLNZ1
AJt43BPBQwvTs0p3d+L0EyquUwQzpKeN+Dz3Ku/iAVJmIYr2IWU6C60DTWiRl7N6Kvk+qTzYkSXk
pyvhKtvr91M4g8Sjih196iUDMlSzeiUWbJOk+QNRKD/tKCw9tg1V0kBqr1Zs19WmIBkdtd4grE14
1EClWwU/Vvl2StQRrSRRAWIlmm+yyOpNvtI0jfEf7mUUE3SnF2qpxRgDgRl+mGGVaCI3zJUjE4uj
MCF7lPfitz7kSewUbC7X9HspQyqZE5dZKHte0Ojl0F1oKpjmNK1k4I2CsWZYr6ifEdiYdLXBta/p
SN5TupVv26Wwwo/YBsq9Ewj577lmHnE0pV9HBH4RZd+zgiBocto7B6111SA3xpJesdmd0tTsXPtY
pb6PgFxjHMMb1jXcd/ffMf9wCeYdXgjBeOzNKgeryPqXIF35XZdEPrGb5BOr7K6piQAizRGXDthI
kGEe0C7Oro7hNAP2Ydur9VNyBfulMQRk/KFyY5tCXcoG5KB+YfCtwFsKgMMatHaJ/4sG6iOYimT3
cFZJ2sMDoswh0pzml0dQ5k6Z6EmBBgUPyT5K7Gkqq7nHbHLKQ9sbZHkXtpAbeU9U0PzWQhYJ5arE
xjARg67qTVzbCMx5jeB4m2kIPtlt+/JSF5WZtYiI3OGdFAsyOGQqX2WEYKSuy7RhoGyJC2gSVkXJ
2i+VLPKBDuIgIoOj/NQwvJIHuf3p6uf6pPZ6930Ibhaqs6oSzN5ThdisRT/eSvYhSqlb2aSdJG6U
b0gp+gkwgKlNkxn3cM6PzWDFHIexOQuVRxfoS457lL+HBcrX8WJdSN53jY1wSbF+G7kvt/tdQzMW
+RPVpgRG6w/yl/+1JwpJJpCzxN/TxRXstEeDpBSledHUzCK7kJn8QrK7EUoDG1/ltXyGnkvHjk+f
T0CxQr/dkHfz6/9gV8v3LrQYmWeJjBidKmj35v3VrQh0u1Z64RfoLbvyJTgIFi6gQSCvF6Je5tNP
ItueaB4JC4L6qD2Mjr48kZUY8rtzWDC7AlnAAuJ5SA+hB1zhFEQIE7InXs/eYx8k8uHeNgiG8ehr
Y1GT1ZmacPBKT8/hKsRU8JTpHiitXqM3EQVo6GhBbU0XgMUr2VwPUS0o3/o8vl0PmzNwxuYMb86n
nk49+tiHs4NAqS2+fsjozbnAnoJzynXNYfVwUP5jHdIAXCD8ncU3hNUvsma63T9ku+M6G0l8oCBF
95TOw0VTPmGwm+93Q5wVIWnjI2HJNQ3ufFtk5hPjy41oRBgUQgjoSRxbNga4RVR76n7knzpsX5iF
Y0E7yBTma/VGA+mPBiQ9a6VoLHL/7xvjwNFLdtUHGYny9vwjF6vA1eLVHlWO6wUM2i1kTbfcy8Xz
me+96pUdKSuClhoe5WrF45bwDhz6kWI1uiPGTyjPnoiX8/K97fk26fWinTxB8Nu/zO5AmVYvFNZW
pi8uWp/ye50rSj423ISwGc73kXUDCer2NGX0pQRyIM+nflAqA3HH9RADCrtnm8GRyO3d4gLgK9sT
ABi99dQWuHUT13vyCNyjKS//g7zMKDcr6byG10pl1c8n26lySI7izVNaEyf41g4ri6P47gxTsYJ9
fTMyrjXXmvz3Xe31Hr0tmUTkL8LshNgCxOdvyRulO49VrdFz47CLFIWOGh6jxhmUTX46YwVtbPpd
PiChGqQbiji8SgjMpXNb4oaUPUqR4p3Z7GT+nLjhd0Ft53A5l6EZwt2YG7WjQX5M48bxTEXc9BQ2
QoZA5IktLzw4FlN5Mpo0zbySY3Y99KDpjjzwyZ4hfuAtfi0ab8vWhjvMzIYdkjgV8kWBM1NYH2eW
5Bv2QVMxpp2ZokFgnTEi/b3cXKffW00qIJPjGuj53oit7l2nBH5mHpERbblJgBOb7CKXDHS344w4
9vB3WBtjWsFvZAMmLQxPh5zNQ7H135QzC8QIwlQmIAd695ZETjVP1iW9rAzc5a7Tkak3LehbnLcx
Ud+Gqlp1Evu1Mdy4NRz35ZhTbFlbrTZLl4pMlEdDe7lOpLDpglwrQUfnceiNQNReJUj44TWvIoAn
u32lH3UDgrVNN/wC98dHwrs12c13QGevzw2SCLyrUySsKmzzfsbcH7Fj4FWIAm5EajlyXLS5eqoA
RRb9OgCkAUng9Y0pWCSzoyBT6TTb/vTi/i1Svb+RQcCm2tL2ig30EASxcD3swEdFf8ttBaIZLXDr
y6ydUocSafl+fYmb4fhfM74ZaXEbnlI2H2KMfg8qYe8QV8IhHGROnCCpJxu5MYMRef60f0Di3Cew
s9HdKSBY0J2mNHSbIAdMdpMym41f3je8Cmr5G1zzIhEokKxmd7rrMxgNjwwgxJ/QlXf8tMXPfpHf
r48EitiF11V/R10xY/KOFo7F97s37tV1ajlZFO2C1u85VZ40hJQ53fAghHSqyK3il7X6MU1ChZmn
M2IObevPlvtGyv/7gdJ0YYIc7F48s8UbhT8qCteEoYYxmhT+fpn8qbcI8QgK+X3JV6P68ptSh5FS
mZ6zE0b/56NrKRBXxBd+Fd3sd8aknLxxF6m6PQPPuaDxqT1UvuIpLPoTr/lDQbPZVv/eYNEM6kUI
wA9Ue0w0bXZR7mkzuyjAjZMQ/NKgZkfCLreo03q8zxd6Vkta2Zfi08a3ZeAK8u+k49i4ZoprgwdX
VwCa9yXjjetfoj6c17PHgwaRJO1y1osAx51GDFMsal3hDc7IzGhX/kxtsZA+sOvLXSHszUEkA3ES
rh4beyIwJ07C1GaYS2gpYnMDblj4yDC0a2o3l3l4C19+/r+xG8KSnkZLzZwkn9jYLiM9tkWNZIxp
WXMNRwH44c/c7bETfHMEN7d0FeWsiI9LLYRkejkDMPXqq4Ucgl4/6g4k7LlWKKkbBO3U5Lgn3OTJ
OPQqWemhf5A59c6sJv5LwwJzHdNsGCwAhU6CJc1mI1rf3YAjLwZYz2M5YSbcRnkHU+stm/PaJAk0
lOVKcj24bFJ6EokTMOy6I0NHoocwmuznXmDVvw+nLv5gdGM/zD+X1ysD3mvcDy4DQverQcD6gUQa
FiemDZSCDFpGOOCRTieSKTPqLC2Da9dacZXBxr0XHjx6Me/yDkgk3URHRhpAiqWvQo2YUnW2RTps
TNVPRuVEbb/TlwPEFC5KhCLFUpyxIKIqYFBUnT+e7ZXTYPTShtf6OM9MKVQx9BmDpkzC92q1RWE2
2hXIO6BflqmEJec+1fFo792YgwstpdDj6Ew/YpituulnKQQHi0M60cYf5LE8F3v0J35m+SeINjED
KI3B6u6X/F17s62bCaoHpvSmudMiaqkj3admcWjS5TdJXL4j7ruPmwF3AIGdnENa2Bw+iTr1aBqw
hDPR9GGP28X9kC58rUMebuMup5IBp64junc6DYGcf2Un3zENslWflGBWNdN9YDLI16BpGTmEy6zX
KCGIWFOciEisC1W4lUZhHYhYxAr2bTQtJ/APQnnFcqAcPv2yKdQkrJjMQZM/XrHsBNl+Mm9DKNDM
2Pn4833p5nwc+if8dZxyIwO+poemkWe029zgy3Takz6CbhC+qi6cTeARy6QuNzMWAy7KnuCTn9uM
15jze4hj70htCZmR28XJuOMKUkLxGuCziiWvhdOGDUNGZNpJg+TsXbyrjI/un7yJTyz6hhpzh65O
jh0diNWnC2Uht6GieOb3q5y8zlfsG1f/iv7LxwQTKkELuuwSJgGbYZWOhf0fMfbvnxrPhNaQhxZ2
Kqje+9nEpPP7BCNCDpt8ifsDAjG1XVjHqk00ZcOJ5GznOSZOVKxk6czwan+uRaLwszlc8BuSz4Hq
6HxEobwqLz7ZnSrjajs4qBz5RDX4yB9ZUT81fhQWiga7+XmIUXc1VMl1TtIYrMMF6B3e8hERiN8T
qrds5ly0OPqgwvFVeKnVm5Ekx26R2eHw2SykF0ZuuktOKHYWO4Ndhy6bpk1gNGCX1RBXSFEL2Jiy
JSgSV+QJLjTg2bFm/y0xDGEB8PFue/4ZAT1NbprdKW1vGAvAoULoYJ3BSN943ddkx02/0uiV4j3B
uX/FJG1RaUiya8XrLZMBAcd6c6Um4F9CxX3dZz2mzKtTrpe9zD4bpQd6HlyBInyrpdPllDRCxd0O
+wZpE4lZhDAuTfBfPuEyyjhCUPXZmIWh8/6jy6b3zLHuEm0ioFx8wp8OOTx66V1yiO49o5sAiiAQ
4Hlc7L+HKrW+uP4FQYbv5E14co03EOdLrv0eOLFwua7D7QQvRFQ8/euQtWzHgVSPHJyJsj/9H0My
DFSBsGcw+na/nPSLESxhEBCSxHllrP+PIrK7BlDPFNKo5xJqAi4oa/kSLLNFcfRDEU3T5KpeqRP3
dS3HC+JFEqUJh1b5XF1dR+GgsRE64Qf4dhlGA8HqJ+ALP8OzimsDUOHgGtMOkznn94M9WR3G8t9X
M9gXlrdixcbGOLg7i89E6r0e71f2S6nRw3fNPTRgnzyqQfja87wAibDQd8dlDyAaQIHoxTWoORpd
bOOCjZjQzcD4SOWMVcKDf1H7VL3siCYqesJZFwzz7znxqofXBWMswp4WmCHnOB1LjAuIB4qIURdZ
NbKU+2f6m2N3P+oEj/b1DIXkgshE5mlGsgvNrPXVm41ocRjYYMoxHpGPRIgmpUKRT3jrV4XuY3Xy
TtnzXwX0FNmfBUTXqSeKbVmmNxhc9h5Nt0O6XTsoleqECcc/axy7aRx6/aQ/GY7/W6a9DBfKeWIb
iNOWmtYvyBIwOhcouwGs5pbmaKkoLw33ntta86JS9/3J/BLLy58bwXPUnUKOrvqsHs5vgBFgnV8W
UE+QpaPFWS/hlLdKNdO579wVwwPDVph3UhBa03HI03WAljRx8yyxXHBo5/pNtrdBEgqnf0Z83Jov
SOPajPuIOaIImMtRGcQ+y6HBNDwjHaQj/BOCuWI3TERGAQZ4CtDIagrJ5rl4QgD4DRBxK1lFGgOR
UvWJYX+8IReluOkUq0dzsGNZAtMnopDAkmKBeMwaNTr6U+X9hVwXyj4IS9ZsWbHf+ES2taPSORAw
TDcp++8/K6mPZOHuPg6hp4qDbf9fu/OKfY6DazU9woUAXJC8kKb1h0vQfFIfUxKOyZQMwF+wmA62
uB6PriVR8Gu21fjU/QiG7JlE7CTphCke5KZENeS1ks64HpVc1MjFBNpseoExPoKg0cF3PcZXVVdy
viupYganrRTHtKXlXBIUsEmiIJ6Kqud5NtfnvQCjjb/aZZ8Niv8HBnnaT+H/zGHVQlZlXBZ1pNxs
NskIk418IGlldZEL0hjiR5AtzYwSd1TTO9XkowX7bHhzNtucqGLLG5OUDRn2r10rP+ouDmUOFVew
uoT+REZef4RTM4HET+PLIMOjCVkoV+uxZ16onUkTmzQb4g4ndx0YpazXhxSfsw0jSE3le0/+qtK0
fGKpUD04V8xkBYMpaDLAcjf3+2tJqADkUQqEEvLJrq30Zp4oGYFacrI8KX/fi98VoM3nFxOJOnI0
UKKUeY28ge6V7rhd/Xo7yO4brpLmO7Yzx0Eec364VVBRILM0G+aR/iEijVGe+NFV14/uBd+q5Rtw
LpiyPmi3UpapCs+s9EkgrJBQkptvGXgq35YDkDcEStaamL7egIkR4WWP0dOPZmUp2T01Kno3ko6I
0eZKCW+DmAwX32HQt1seXr9vGYDIXy/+YzjxoAoyie5TKETBcQi9tdbv1/YKHje82dH/UYO9mY/1
lkoO+YhmHQZ196btjOh8FS8v3ZVeRgz35mQPTubRua19K4BtTWE1+MV03Zi1S96pqawqXc4BJrLD
3c+qPnePFNiH8G+Jykv29dqpTVBA0udAW8kuW4tlwWEGCk458Yco23zlGnGUmJCkdsQnZ0AnqcfK
Hji4n2XUlo/aKD2k7DaAEHHio7P2IjSRi9wbfzc3QkmUegLMo+hht8k5hm5l6rqybRWNp+k8Fz2T
AlofKEj1P17dE+p2xS5LQRM7bDKHdpWP+xKgGTuoa9w6VD1GiR1QNQlt86Rmc2mLtbx7uH5OaCuQ
WM5gJsTZCMwvLAkLG90b+MFpfz6VyVDErQdefy3puSqi0O08rHcFL6DPoKuZFgLZaLn4czkwAwEZ
NG0/1yegL9u7aXh+C0UqIsuRaIoxD1zI3tIMJR32YXJTVW2jn5ShVyNOx/8u5rc+BqFc+eac2fUu
POCUOIED3FN9jjJbZUEU3z6t+0y4JdS/ruN8+Sg/1qfPzQ6q4hxts1m+cF/n5e4QfuKQqtl2Sc3B
bH6o/1K3cebGtGlR497TYbFGtDjBETcAmQRjNbVnnP31RAbOFHPKbs5vN5/gkfaGUQUJ8IYXaT/Z
wz6E6addQldEhr2mWxt1caYv1fJ32yBxnTAITI2laEJZcgu2lfiGen1yAZQrd6ardXytUCNq+Urx
/G6FBQPlo1LDhzp9kGoKoQR59EheArGL+Z+X6hKA/ncwZBB99mrri2B986BkYuYpZYzcmcizK4TY
57tpVr3ZAmyivgu1lyF7ydLomJCSlcqe7DO6OkcYshtgHI2lWowyilgEs0vm+fTNphCevKq0MFO7
gdRkKnWUAodmdtWSEhfuJv4GWvdazBDjcPI50c+g8olYjUkHliK7mRyToFbo2TLexn9wmLMRL5US
WIX/BxtWOdg6UO+95as6hfJoDWuz4R9zcTQtzRBZNHpMABgyxfhAxmgFmv28/pUyGA3XhorDmqjg
Kw61hzaq124AJTf/bqw7jXorCigazAimZPFppepd06pc1FUB34BpQzfmweWEbCh1Qfxc7/PSaEp1
jhBQozpjJVDJB3skUKiGaqISOs0gHVIyvDwQiQxD9Jzqk3NbLq8m4mcXxdeoVhyKa+xPd27Qm8wj
B6yXL3YloPmsMUhZrDT9b9aUzn9XI0GN8+3zaLHKsoLgwnefO26KUKYwppLlBI/4q711YiUxIlXB
1j/yUUkaMP8So7vD/HmjUsiJXf4x67ljAeCjtBI0NSEg3Wac8qB+drwiBXn0NF324GBWDSXLf0Zx
AR5WoqJLICf089UV1rnGXqNaCj89pAa7xacvHGJ8RySAvAGZBaIdQP3dxfJbjzg5YSxP1thHmvo0
spJXdYli7MX7zrYpO9xsr1tM1PB9yCx6CGRukeEXPpRJR4CI3jIYrmcJiK0b/DdkDsCHZoQI3IE9
kwwjJiOZpEikVrdqxz8WvRyjGdzqZafP97HzyfrM1f2vkHHwv64LZ6YcOtgatfWc6DnwuoYjTvSs
eRHfDvq9nr88zzHVObvI9cWBAysK608hiljT5msEOE3v2elzGOZjkjFJaB9xjVQx81+Oa/5eAFFV
w33hqAiKjZe2yqKXMzSftbVk00Rg9nEwVmuJfuWLYy4nVC1OC+++dWGm8VbR0pRotcWhVemEiJ8P
E9mziLxW1Q/j4GrqXImG1EbqS/xw+qS/V9nBhqjMxuz7B8NdIzyOdBaTNTp0fNqUgw/eSpkutunI
VCzoKiOeRGm/MkzWlMuDL8g+OYp62e54CT+VR/fN6pAnPDEXYKC69RpemTFgtQLniyc4YiCTUTOG
zzC7f/ncZ7qcveFpkoZTdR45OPwbPBygM/srWQ3+GWanhETCOkOwGIGTasjsbuhUQ+HpNwSyVhZc
eLhc0+Vm3Th3VQqjGSwrObnhzHY0CiC6JT9uXeYbOkqVba/ZntndzoiP+QfP7IXFwF7vGEDPLAAv
vLRvTjjEskBhXH7h7zgyKHJn8fS4YfL1C2WSTXv4RycWvL+mCS1A6yV1jdW8DxTpd7rT6JXE+Qcd
DmsPAAh0pqd/goNv2jD4UVEi9DRhpJik3lGlnaPo5tPzH8sRX9aQ1aiZFlVClEp7MbSBxkGe5O/M
gUw8Jk6FLUDOakM9bZYsSARXm/D04Y4jxVRGehbJh3+8psrEOFQJJLMgXrVZGOmk0w2lfSfroT6O
Twjw0zEbxN8A7u/v1eWA2kIbOMfOMc7q91zNb+ztq0k7HjYCZT4huTI5NvY2dp4sbmTaoEPtEnZ/
1QJBeMgTsrlVKosURv7CenDHDEKtZqhde5P4u4WITHLKVsMTLkBhyFck8S155WdarFDa9IyFUMci
/6Yjzu8Qsks/f5yb+5Ca6qcZbYh5n1BpxjtJHnekvQ+cLnZFK1kDFY9nQmXjS5RqbEc10hVUiHjT
+q+nWycpCNeASw8X0CMFaj/Amp4h5WLskbNGRW6AyvPvKb4XlknMNgE+rfmxGvFAGMjh44WA0b/4
irO7sEk4y2ahiEF6Cg7GJEMroqOZ5LhYevqAQSB6MpuiMrGqibDJgAtOD/EcHDicG28/L4yj3xJ9
ryZcOPYqjXS4Swd0pjvqPqDJJR4KfU8Bpkn67iOzKoeUYuTsBcZnbAsZlMx9F9GYIPD0EJdbEzg4
mtoFu15nGmpOgS1alyXfnmdz9bkusmVzCYd8l6DiUaWgLq2fm1t3y4ku9MzY6TDJAnqmMSKoA6O6
dIhBA1zpCbzli2sUw1picwfdXdlWAW/m0608qgIBk0q6BKfES7S3sX31vJ2CKxoGTiGyE5JjGqH2
aN4/7wP8+8tzaiZ9EXxS3zqtQ5UJyRfXTvwt3MPG7mZGTfYq/SF6BQfkGRxJxrgUMh/bsBuy9XVc
pM1MJr4+yFefq9MS/N2EiKxJgZhO7N9kcCNk7XJqf9LCihL2DnnjnatVys+/TLQqPKcw4380isWI
Tn7hmz245Fue/DKFgqBx4e1r9Gz4I13sQbGg+SYpAwNI8xWN+lW+J6FrTY/I29Z+FKedBb63mIC0
m8AFk4sGjX4mCXhBhWeWW1AurS1/Ui7hCtBKj5wxOV5nU+xOAEpd6s2pNJ5G1z1czw6OSRK0x0db
hZJsXg4ayDG4CrQBEs445pHFE7oW3tuiBCWhWXKFaLtHcyoqxDQz8f6GTt1fdDT+kHj8kgECTrlD
lT29Huv5jp0395NK6w2X9ipdUYXzy+b/VT3deWY9rDWa/lQy2HhTbXPxoVHvKhFtezJwaB9sNMZy
JVIWoUrajV8oNUAMvZehctF1A8lFxmc0IIGXShGxxqBBSNj8KZtJtRbBu5jhY3JDLNc2PehnGj8M
U7KPnBxRHeOobtWJ9PpWDgZfQTdNoCdNLlcq6pB4DuOhIYs1hzWG3laX/pdWN5JmxYtbn52USym/
0jhd+/o7G1aV9eTiTpT/FPR+3Jhz1Ocrq6BnI5snm33bDkZDPbdhvITzD4YNryDJhPl1+5Jn7tdI
Z5BqU8uBtIO+MzvufPNw2yPjxvAcVHggihZTphvdEUjbSZ6T6kWENa4dokEcGc0klLY7FQO0ByBK
2HkhC86e0Stnu5MvpPheWyHC49NSTrQ49MPferbjqoA7ktAzl4yGSsKszk97jw7lfhs34QqfpG3t
5R8e5NRZ0KvWzJ519OyFyzzN5u7Ogj50LXyDXvJDtxLtDaPinlP3KeRgxhblkZTGS0ej0D4p1Pob
Hl3l+QPZdHxbrOF2NS3NgCubq8iHYMZBAYCulOTyRPug4L8kGlUz+fAmLMAABxrxoBkbXiu6eZEm
226f/sZZ67rXq9DgXDDhJ+MJv5+DDmTI95f97eWMauzUdADshHONhQFpMEQsg6mQ0vrVzgbTfRR6
G8Ezi0ncDJm4MlJ4FINnckEMWRRDN8CG0+ZBtLmWp65vs+2kItTaNJkJERv1qxQq2ykwrqXHfAdj
FwLiHpta9rfMw+K77ik+pJyeuTvpwPkLDTmNZWVPRse7Ou37NQIbYeibzgdd52bFzn+CsTRLsKrE
EeJJYJTF6E+CSZleCR74lmGSd1o5dG/BAth5oNFH4beOCXYtBqWMKedGVKs6+jLTFz6NTFUpmAJF
b10r/lryb7eqqYr5j4baNWumh9GspExeCg+DK3jjURueZvpcJPXAiOksueN6qvnsqc857V/uO2C5
mcLJ13udOgmq6VNe3YsND2RyjkrmOai53hH1A4LdKiDnfUG9pEWRtBlO8vkEZaZtiSZUqWgdgh3y
LvGYWYIqrAKuVBMQsHjiXnqoam6q8Q8RruFtpishoOveLbiPsqLOF9gCublExY6iDpGCqUPI9dw1
yJLlC8CqHagXONU5JaS6pxWlH4A4IDm5N7tGS9ZxemBP7h42hCy9rqwh5ykVnx5ZMOl6JrfS0dSo
Kq05dB1aMx4GzOuPrFtQHcy7aBTrFY+sHlM/bGBU3kziPi/ca/t/4jHwWTAhRNpRJBD2ePdrwyav
AmKxsq8LLKE6PytjCIugfznDNff/cA6smktXDq5ZQH3HTeF37s0Ibr4vjOXCQ50M4ZbEBxDrG2OR
t6LYcho6Ms/iHN/EYuE7i6+hTh8TULhwJzhM3I6seLaBrGOSxGAC+syN3Hh8RaKgbkM0bDslr1f+
+dI2tho33oO6UvMFgL4eX4LhJrvHc9qggZ3MPhJ7zhw0vkceOsnxkVZcaPtDjI1mJ21lz1BfUEXB
Xa/Xf8qj/GXOTdDTlMqubOKHceOYkg116tSMv7veIqH866JO4gFuymdUDW0doVTfIeOczptfO94t
hOLdfNS2cME5dm0R8Btln5RKBXzWkq/fix2HePtW9468GLy34B+S/rCqGA6eGoR4xTjjdPS8drxu
WjFg2e94bcmxLP/kWcqKwewSiWGt+ywtotkOghgPhilYDSTuWb92UaErzsiIUxwGGplZ8oOzUdwM
u/QWC1P+bDmDGLVxschIqAk70QJx6CXHfDBlr9QOO4d96ovc8dwe+oMVSRuvvDsIz/EiEDy8OK0X
urk21SnvM6qVMGU1YJTQ7YRaBOGq4Cu1fjfKuaPV3eIVmQcIRupBNVjmtZu5r36sKHqjkV2VZ/J/
n1SPsjauMy23NEYb8PPKxIf+0s1MHLfKirWqjKfw1gTZojfr2RncBTSoLzklXkGDoCaRsu1K3V6+
Il91+8el5kLL1hqo3MOs3WKJ/lsf6KxF7+qbVm+f+cUQwYlKm49LO1hNxObVz3ndSbmfF7xgQ/Y1
yMZvjswPe4XRV/4NBAg1IIfzo4PrepazruIV5e//BAbW87ciNfFiQHxj6QgTfRXxzAu5oxYuP6A2
YOOGMwK9oMff36pJRQcrmRYlICRN+F92O7jK3zxF7PHs1fiRAzETZy98gddBT6/SdXpyHM5duzbK
967wdbwsSVs028vE5cSGIMfwpNBDYrydwzgMtsaXjsvM30MPUgY2wnDNaHFeIp6eAH6sGIN7JVR1
EaPSQHZDz87efSssrqjkV39JXGv0HRdZTu56vpHJTlbfiz5YmJYeLz0340kNT5mrc1ogTIvRuiqQ
FP4xY+QwX7R1QsCvdEdkPb4dsnKXItURF2/i8FIJp4cFSW0WDphCNOeVJYex+Y/Yb+idTkiQwMbv
MgmWT/JhgSY1Vlh241XTQ+2P76Ub7nt574He2wQIBCBqmehu3piaGoRpau9ISdvpimxRpwdSLfV7
eyk4ZTzj9EiLXdt/9HkkU8/8+6ZYWOUSAkOlYa4D7CNu70G6r9v+MG8DqXoXAFLU6QP5GETu6i/f
LDcJeRADVK8W3wEiHsXMyge2mF/awB4cTQ1sAUtrm55WpVQZfZjqZeNKbck/HwcsZSZaqRphIUdM
l2qEmYa9JkHkB95ZXof5I8yycsVbAXGu/1Y2gJrdEfKieMm3b4jSeUu2Eif4H7rUsNHYF/X+Qs5h
iQuZLzhFaVvaHN5ygMF/46jvz2ZIYh9eEl2ld2QApPI/iqmIth0iY/9ygbrUo5BLOew10anocANJ
tmq4dFpL9OMkfcdDWVdPHXnDskUmabiYYbVlytRE8qBjJ35xwTqZa79foeKX79nOeqWD//fXOXjL
e/ZeX1SZLAYYq+rmsKjLMunqnAexd2I1mKbO7dIQIRrLm0Y5+kzmo7NVI0gjsflebNol9ygt/pkq
KbNepLhX5WIA5+mRvYgkKN0lv8Xojlao6jxm11rRW0vso8bmYz4z6DpkuLTb492Fu0N2RyNzVgyM
8xWs8JfOmb+6Crroa5QFO/m7WY2EW5inq/FQO9iv9WJfqQUv12XHM4/NiuonOclgKpuS3xc8US+O
FP30rirz5bVqwyPWsK3dMOioRYH66y/TSZ9Ysesi/qa7psXJd2mZ1YLAbix/YQC0UDq7CB0c6Wc7
Ttnu/TUB5zO/7U/JSrZ5D6wK45G9MwB9UmcnboQNupQDSXXF8P4K3Rr1hgL1618YCEosKURfLQ+n
etVyutJYgiQ5s7RpG4U3uPjkbpQG97cquWUJIvgM4sm7PBaG1txBDqHW68jxWxUdcwZUErgRoae7
01CdAQr9ewKLaqZvmYYB7Whui3wdA1HMoaCO0zOJBqzVqQmP8H3138h/BmqHLUW0ZUo2UBHCfIsY
DXHUcTetuExgXuPMbFWwEdVuPley0h3MSj2htjsrbOqq2UhRZGZWo1XHHl6JRRivFhCoj3YuceEt
ymkhSOcUCXz2VzoQRj7s50whOAri0EfOBazAVq1n00cjxUdBgugxNktVevlVYlzw/XBw12wk4chX
BbVHZegKXR8AURscwIE3jxLPs0RAnRphri1uvWGVGr8njt+CVK5zILBx19jYSDuPFbA5nJwjGvIn
M7fq5daqhbTA8aLfwBB5Y9CxoJq6nVQv7NbA9PKG+nPNjntfc1QBZxocrVjQ8mPzmfXnEZgscboL
1T8r23jZTq0Dt+9zRA8wonMLjCO74mTvhxBYZIi/xEubofJAaX0+NldYLvmzV0pxB79msUM1RwxE
mZZqgk+gCOpgwAQnDS963irYM9v07H6obGRzCj0A4EddOHOCa45xUfYGBWhoxCzZugY8IY5cvl8j
3AUv1oHoxgePnQztI88jse43hjTuvBTOLBeWHDH+RLwdZHiIXTqG/5lMF6EHz5CtkEJoOSOf4mvY
GXr47dMyggRI6VfTEQfwITLt45hWHHqAEdMJqy8RhpfDeC8twxEu3FYu3Rm1eNwLivVPQSInKeC6
lMcS8DWNq3vdqp6q1fSJTgM0ni1Bou2fLA57nMIrUwKxxaNSX5QyJ8eU6N93IdU5Ppk2C9NLZ29K
PkMzBwaa/bnhHL9dqZRfVJLbCfhxkOSAMpqeH6WuiLZ+lnKc5rB3aGamyHh+DyP0v/lJBtd+eY15
8SQfSiNl9edIk7o6t4sw5BkmPFADP07yAu8/VxosiZxn/A9dFTRN1whz1dXB6AtpzzD7EkKOqbrH
hcUO/zbUze7+k43MwMt8W+ZeOdNhWLWhPkWtIuKpKAb0pfOxN/oRhfpgJtki17MwWEJtHgeTIUOi
xtFXeXX9pAbs23sI8yQIUKA5n+AkOjdOgCnaA/RS7z6yeIPi4na9beS8H2M3ngIfRE3tOZfjfVcx
4BGb2vTrXLoGqIFobDYyB9ZS+pIMsl1waGzQYcvb8xLJO6yIZcrYXdWcAipEzCZh+By8TX9zcu3U
zud4d8ME+xezCOJpXxPffoLt9S3AhtxS7lokxPnSscPTV1ekQWBrJ/Z84p/A0n5Svg1iLz6oOu89
Fncw5yhpgmXpc/kNJ2IYtiUVZHE7RjV3bcZmMVK2HGPYdWMWhWIu2S8+3MwBnQ1loUKrUdFiXRlA
6Fq63HcPubmHlVDvXqyKcsSluvNRvMJm7Z7gbdG96SOdz1mCPLfu0vWuYlR4iSWY2yY6crKojpIi
NEvHrXailfAK0V9+eF846IASJOsO308UAVwoWWqm5cYWjo2eGe896lg3sXlQt7Pt+j3uCcPPS8w8
Rea3wuCj3yQ7ZagCQl4vq4OjLyi9FWMAv/o6ZE2GD6XfSwETiQe9uhtOzjP6Q2iKV+dypxjhOLIT
77pc2rAQospjhUaqefIP0pPiGVjWm1vMioclpas7bs7YpGT16MU7Hl73EtSnsBABh1sMano+m8wR
VNsN2ktvIPWUBYXcTop58rizlPLZfD8j2vUAd6uG2Ul45vSz5PcXLqWRtc5B2YDKYVe8DM5D5K/7
aIHCMwHjE5veswmCqsTk9QTfeGzIXB8HlHcB8VZAxrmavV2M4gPPo2y1I63jGZB99AnGFPjuxW4q
9+dMIsOOagBFvNvtBNj2xNdl3yXQA9k4ceDc3ywBpzvZrRs0idTFLNHy0qYwdp9N4eFKE1NAwhKh
8qgdjoOsKdPfIYgNfAeE/yjK+ChXx3YKiWrl9a3OWUBVDRyk+gY+PEFPwkXRzL6i9oBehus5oXM6
e17Vsue2QfC8dCieWNWJJue83fVGmgYxGbbqAI0bdwaM3ZwXewEYw4AxJxBiPoEpGwrYNKgvRdcs
1/F23cZwewTfQdM20HI2bJ7NfMSZj8w/E1TekpGED8CcJOC14nLh6gdeBp8236YejShbX4eF4N+W
x8QErq48hq9Trc7u8EDf+t8efWe/6pcduIYbRl0wfDjJJ4I+ETKxUv7NFX8MUW25KvPyOcr5MKh/
o12idsQ8QgCHPz03CluETbYfQR/ytYLoed/CTJhFZwTdBYHXHEM+5DgXpOHva+jriGbWAjD6bejO
g7iGsg4h67HPYCkLhb+SIWwtWJmXA2Ww0KLmxh1amP1qSxcitSnIXYVhRzuHj9HIQIEfHWCtt8Uw
qmOeNJqBnThHFVlGnwpqg1xjJEWJQwoTkedhag7YrsH/ytK8YHBqJf2EQJeiSnx6z6wTCj9Rr3bJ
jqNSmW73Ky+9tC/N08bzEfvGGFe2kCSYH7UOUYfR6/bnVSRBLZ61tBpNGD2oYBPdjM1jOHhjnTcp
lUJnEG2L/L4jZNGUbaVtxrQ+mpXdIJZLfX+Co7wZ9Kn4voa9mgyAYUWNm3FpM5qTnJ9hl8l507Rv
uExTCDqEfvZMxtaH6t8lk2m7ErkajZaBrOl5XiHLEmpprmQR1hJuOF7qMAWOISk7uhcRQHi93sKE
V8+bVD6BUcTkTk2+9bGZxLjcKS+yZfBvXiQL/cnGBKKP0vy0RQA7svBfRhrU51yhlpIzYdB23csu
qgXQEf8eqwmyRc5R+cA4tdtc2XcAumM9+sGLLnPYindL0NvhNgrXcKt56Jw758cqe8D6uwM7F4uh
BrJonSrJBpRrz3qYXuhOvyN0+10ngfTNlBoEnu/kaHxlQqYKhP0yPTjS7T1zeO5cdj2n+kaz4PHS
N3S/XAvGZrgdzP0imeLF1nIEQT+M/X9bhtPdXs/dHo00OmOhz6TtV1AFYmuy2orSQn/U4yWkOnSO
H0zFN3rSnnFYKeRxVRsh1aK/TqoCkIMcGJMXBkqshn7fchck5p0g/E9EmaT5D5UR9sak63E+J3KZ
dGEHmMZYeNHnwSRexlM6kmqX0td+m1USQLb4fkADlqg2RE3SLbcsMi+OCljJIl36hVbsr3S2PadR
yvUe1AiTfcDEiRW5qrwodUqDk542jO6E0z2BgH0D6lHBQiF6WZ544Ix1XCVyyx6vllc9NOybzlfp
J4wQwI2NTl3mq8EEWyH/V8WehqTaG/wO0vQ0mIaaz5scXdTkZe4qgL3L63nIn9VpEeg4h2g/A61W
IQqdyFDJ0Z1cxHlfW3JVVVYX4lqwhUJVxP+wjoH33h3Zccm6ch66LIxB8HGKj8zobd1iAUuHBZnW
h59kPFBE8fzABWH/8W07hmB7vrqrI1sBg4GGHWZtPqhqjbz+7R2tIA51ubmUeZte4hXDFvc4MXrd
+4a9NsD4wC7+Vq8EjaLTe7NQEg3lZZzg88DkghW22T0nugVr+DOit2gVBBMyQB0e/LAdDkh5jQdU
S04PKNUal196EEj/2ucNpfUQY09w3yF8rKMz02Qd6zdkGUl5kmOgVp13J+xdHp/z6Ak0bNvhagA1
ZErzN5hHlUfmusKQ2DgRg9ELgpUICIb7xAvGW8Tp0luK4arsnZxDXB1VuunxlF0iz086oRKwIpbB
ohJDvnExtLpjzcEaeZEkaEkyZ/6XfAoSD1GRaMZFh/vssCksp9W7D2CKN4mD94sLkHdjHAwE2n9D
KydMG3qFUq50Bs3HlQyNZ96y9yUsgpcliSzDcr6ZZBDf0N6a6IH34bZgwqCQkeelhLwPB7AkU2My
PRisioo+KKnZoZTe7+DbgTyhXiseX5isn9McFAxw9EuNJE/nmIGa12aA7kgD7QucKf5ErFvFe7Ah
k4giNK1Nlf/hJl7g6/drHasZ4kynqq3eqoi03kVM7+POhRxnPlS4ZKIW21jJDruIEOsnqQVBYRxS
l0HMf+sIRa7WNU9evrghQpftGopNmvSLMNIUDyC9QNjuRBTLS6iltwgsmDTUobFvCpHRpULOLYcp
ZQ0ImItaQPEIL+whRXqhyggNjpkc8SOZuhzMu9RvoluEJb4p9BDYXW5VhkU6KshJWbRi9gny7mos
XSYPTDBc8uRbBlUr9wmWLAP+DBaYPKMsWFxonCj8eid7Bie5sqJspDTs5EqFnjjBuMi85s2ukihQ
EHDClrEvH8MLFdTYUi/zgj1GOGjCHUSUbe0zp8dIFm6cqtIdLCn+CJtsQSKmkQt64cy+bFohYxx2
LIVF/eyn1/chgbSYkge7wmVVFJUtavaiAWK+zbsORjVgIX3yAyvEJi6PwkA7ggjow0FhMP72pTQh
ap1LR0hr04O3xD5/riLAR9oLDArIqNymGMKeXVzn10u6eD7b9dxYOiUgiHZxcDRTJZDYiLW6b9XQ
Gv2WYjmk4i6ZlztzekJkqSGnRniHY0xBqFF1k3qWtmRylVAID74Cj/RU0iImbfRCPLSj9kbVIWV0
VROl87sg4ZekyjtWCP3OIBu3cf0gXGW74o6IzqUEGnFtY3RofGrgt772nKVrRBSSdnizxZksvWTB
5rIhcisQA2+3MEkIy94VxFZ0dKUnIfahDloGtzchBNe7eWq0XFoliAxZCvnZTYMNVzGPpkfxMpa0
TPwlFhwQe0nHZYo8sQvC7OHsmtZ+/vdgtcts8+nHRiVzU74ZTToH/5Bno1SoEJ6W488/4JlV3heK
7zkX2AxCwnlwK7w71BLXaDAYWtUCkODBZZlriDWQIGji/UCn8h2dbQcRBlM/qdoQJnbiIi+hl18c
byB0YBEywKAtPMT9aI4qsp75vFd+TqNMsF/9QRcfNIBHAHW3ziZvtMmdqV2Y8gAmg84ezfmPDNmL
ubourKYfAhcWdm0WuP5+8BeGoJCWzfEQWr7kSf/tNpDTPd5hfk3uIt3jokjNuV36mmuQTE3eqTTh
QZdnHXzTau/0k7ZkF0SkFrowpR810aaKYbX9xjA77iCllr5AdBe8nV8IZkk6jpWaILRk1OuGIoAU
rug7T+lIQKkwYJcVoMMa5j+3OG0VLOqWsGCnS01dKqR8BwISQd+UNnhGCDdRTJWRyRuVCnhOE03A
uXr01VU4CasZz8deMCdog2i5RM9XTOrSkkTvAxXLDu6kNGJIZX2+ogr374oNiSdTkcQnFtawX5r1
cDjNFMCXVcSNf4I7t71PFrKEXoUhztBkJoVEvnvH14DWClHwlvlJS90p4Y8xwaIy3R7FvLe+/sg8
CCmLJtndjIgQUUA3NmyMBH+s6s6DzDGhHzzSHUiSfxL7csMhtsscZIUqsZvFR1VkFoautEmMTpSI
qxPsALcbMbHEbyY7y6fn27H/eaDrIw7/MzReq9sdtOcdiW0P8d8cY8Huj/jqea2yNyZOLdfLEA/w
2F80FJOC/P4MJ2mTqa51b3pOrBzD3Yj03ttUKi8cUjjpAKtoM4ZyiT9pG/37Md3eYF/tzDSsO+zm
X26qvGBCKrW6eurMmMwrx2KqXPoZHRfohKj2dJk/la238c7h4+ztY2EVRMuKTEpxH4a2cbHNLroF
whzRtfycPXmFFftU8r99Tqj978bIKdJMb9QzmQPNfIsTz+7xv64nbnINrkb+Ec5nDLb8MvWOMW8w
VmrWKFoFx/e3IhEmv/Z5MaWBAS2DNZlF9p7GxyzsW5zSgPS7sILu7rRN3lKm31+XhTDTiTAQexXk
nItQZ+G/M98pjAyJl1wdKAXWnf6x19f9jlefskqlvikOWWqz/fLoKDPqln6UfE94g0S3rCtbyQwP
Y9w1dyhW82+mGkKW1pZjN41+CVwsB0RLeYYKaEdl6XHxVWu8RVXJmj+ZUWSDvN7pvE2CyZ7de+Ni
+/SfgpRoHxHJ3UTsKPsxIzybKtxf8vgeH9LWZPuVRg0H52SEyfJ2rZwCLtwXzaqxOAhuW/FN/qE6
Dfm2nhg+V6rkst69Z0ZS9XcndQ1go0qR263Ad570RUJzY8UC3fX9SJN4BxOdP2f5a6mv4GRPmQ1r
Va1zegkGiVT6WNiWF3PlFn687ORalfgNnejb0c6jLqLzcApkON1qEbs5ZMXBumaYMDpqLVMjLnfu
ki22QsDSiTdyJPEwJnIqMNlbNChV/Pet0TbjbUuzim1nPC6U+yCJmUWXT4zMY4LZ6vfrDjss3O4s
F8dEbWvbqTYeaUYbSSPZ3irvpi+HXuIHF5Y77IPZ7hBM7f6elhBkOg191ku0DXyXILIk7oK5CV8Z
tc/sbCXDU3YCogqES21GdQKWTr2zobvmQPYI6z9XXBKckO3l0Vd6ggrxRorSlqmj4hX89dEwcyiH
u091RFK1ycN4JDnUVd5KDG7jPRc+6LYGw2lP665VOM5Br5sV34Kz3+yyzMQH2SvhAxs658GGynDJ
08qw0kxFQFMIqWXIhM6JeDCG4SQeG3atfcb85tD1Q6ioFaoTzQj4UuvWNlyJfuyEwZT3hf0AHrlK
RiMVxNgtTJYn4JmvCXf4d4GCAE29XqAKwx5exh2jNc4yyLSNCUXheaD9vTAgpKsGCbnXRXRZQq5K
3CI3T4To+yimtdM1Rs2y6hHbNQeinHEO1eof0USmcQKacUUpVce0w5IlVYwjM1a7VnsfqeOM+StH
dyZaHhwD26bj3zjO7IxGiBA0VBNTd/eQG2w27CNaHP4YY/K6MJNBjZx34hbe/SSwKkdwrIXRVeEv
vr9tzmjggiKQOtlnsjbkVOEYKQlJ8GZDuJ7CllJIWhwltPBXp4cQF0o5wQ4n0NUaeYw3f/kfG+SN
RFPiU8j4qIBeEzvYtMRjD4shFTh8KkbJ/BkCPhjNhpoMGSRdPuAXVbfuWE0jzZLGB6tBoEXuzh0a
Y4neoEUDqcvu8FfcZL4bdeeH87tkXdmf0RTSjx6KTOT14W77qj3mkq11a+xl+LwLJGCM8nxrUrTp
oX8UYkb/Y0IczAJlbMVarKPVzkrlyJEEQQKFul/OiAl09dn/2XQ9bnpZ19HEceSRYewhlMTCDcmm
u3iqCve/HulDFrAB3GgHQmg4hEFk1HjGchvP2PoMyoCG2/qJdU53a22fjdhSq01Ik3dFqulwrWcU
LP0+IEWvdeGdBheDnamjv/5xEN5qz71xfoxcMUPy4gyoEHdgNhnEfEM2eQQZBytkJMK43vyGiWod
3DaV9OvN91pHet+2N8HGsMA9G/56m653s1R6Wr4sqUOzL4Bqy/l7itxrq19xs/fyPC4q2cFxEzY1
OWSZS9rvVw62SFXQhCMA7uvxEIPPi+05snRkQj9SwONDR42VABeI26nmPU1nMGLDXDT20gBFv92v
w45f9qkeWkYH+N1lZpGa3CHazFYxa2Oh4DNRoNihYHYt4x31EnX9/CXSgnxG2JHcgJi+DQ3a6nTp
YPjlicGrMXwCbpBnUMrRr2DEt1TIkfgZeLqmXSQZ9VwXtKaUdhDZfu4iqlF+wfYV4x0M+PnLLW19
YoLswwyMAqfc4uCX5LphC8IqjgZwTYl+tgctc/ioySNSWADpTn1nMqeu4cmPozgHQBtjEKwHorah
zIEkLeBWKfCEKma2olb9nCvg0o5WMmOwXGhx/rdpvfZ9yy22XkEHOfU5E3yCxcU9TK5Hvjhse7yH
5zYBdp38/3atsDXGUZwOiCY2nc8/wXIVlDHf3vJjYAIxHuH1AzGCoYwzqVWE5islc34sqHlPL5cI
Tw7RiyeTXR9OAxg5WhK+0O30j6sOYbEwrx/hoeqadeptqfQu9KVl+ZcQSClWba83UhIiuHda8B7x
pqQ6MDY7QN8MKXbqu5c+pGWqIZH0RmlANU6M/U9pkydjmg3cPAdnPjPz2tW/MsVTqNyIEKYnfEHA
zJZtLNVp7So2ureUVOFW4oYBFczMLkeIiwsmVXiGfOWygc5XLUd4jQSmeh1OK4+mx4N6iqMXRBSt
23pGfFmjT0KklwMxw4W6sxeDfdWiMmQTF6iJj+at5gwJehA1M/zHCX0afK2yO4aJDGkA07i0O4dJ
JUQA6t+ViZ/CHao8xfqmg7BFlcOtTmyXjb4WYHhIxWYLqVCKGETqohcUrpaOyQh/QhZmT3yzyccg
WURnA8M0dOUde9qLcnT7LLsW2bUQw8pLA8DGe0ksf6r3ZzcrF+7kpGHIujBfgfZL/CTAZlId2Fmb
P8N8aUcQBEdng528bn0C4foKNWkm90MoT5dZyuZyQzQ115IRJCOGa8zIby6ZoL3DRmhoVuLoMp1v
o45j8YEbQHQ7zhtI9SaaogHoLJTv811rAm0nmNTPQMy5YkljMrXKVyDHrCCbwxDZrVnI8vZgfbVh
tj80r9EX0PbWdAlubcwwhuZ5LeTHqihkyMqw6Jccfx713GrmHtFpCGs4b9H5Cv6DsO4aXdKaB/6Q
6BvLi9tUW1A8tlwYE5yn2CpWK9iG1t55kYct0hQG3VnzeCX58kEyJA30T/LPGQInCwEi/DT91zik
8UEx5sk5cIVV6Yngh+ZmmGT5lA9N8PhbFrMToJOmmN+3XINi73fxVy98hYkQzIDl4LMb2FA0wdPS
PTetdrWXsNsLaAx0iZbkreojBmnbowpekWNj00TO5X47relLBO4VrXoj2/DY8L5xl+hD5catvAOI
6rRg0F47EdwdasnO27fsI2E5PSE0zzeC77o/qjl82Ts4zXD9m88noHEMqzSGrq4VxNIRWP0ZVatk
YRL4czlqTS0t6d4wMdwYngcZvbW88jbgHrd0dbod5TgDfiJ/Iu6AXcJtBrw12nrIltaEOzxZrDZF
XmugreGRxoTO7+SZLXP5PRqd2RBGeyto54gpybwmPL6+WWPy6RoxpiNrOu7vYm36E1pDaw5iuJMb
npulOVV8sU1rZTmidK39nzQwkS34vt9jX1e/RO2h1IQqb3tq2ZcRoiNicYHGtKq8FdYRBGWasFuj
dfKipEBOnyEtMbQE2BLqCot3iDchyb5AoWZVe41dd5Fgx6yTV8RxgQyb6SfRRuWVNsBa65mGXlKo
gIXZRN5vQ37mVzGDeVwqXrujhSz1HNWWB1OZkZ8qtvMCdO5zTNqcqNTsC3Vztu9XXGOFNoo8HG8+
wlaY5A3blM0Wi2kDTz109MsfJN0yakGIQJrm6aU2DSF5PEvDSEpM3c8LmvjlbkF2wXm+HQsoGlEL
TSz5DFeko/RKOkzqvTbdyJQK+91iqpe/jnDs/tGaleTHybznXwWglQ3RJluFvFrqowBPeEnv0EDd
lwwo2hs5sa7yBaOYMMVtS6Wg3FeMJHQBTM5YSpRWkrjgWv1NAPwnBs5+pOqL47O/JnMyyY2dNsai
ubHfppn7CBEF5K7vRLfKinHGNZqOsRxQKQ07/Vx9WyDfg4N5Gl4Bppv+tMoi3UM+WtqwRIHdB3GA
RlkW0DRXDs4Rr7iq2qQ9uE13t5ef+/7M85ceRBsZ8AgEgUL4DA+hDhvvoAE4vHWJwlMIRTusr4Lj
P1/x4Ip/+CA8ue+dSp6Dwpq9U1AAZySZKvUbpClgdfcANvFkBSDHgs7hEyelda20AMpNMswfyzoA
WOAZurFj4pA+uR7UuFb7zLAow0/FamfH2cQqjURoM1NdtbmQhpRDe5rztYKxPSFJNRhAWGqVXclD
wHTQo3HE1nfMwKl3ShupLNVQZxWBYaQH7fGl/pB8lArUmi4gO+y/FlAtYosi/YgmDiX/P5dVLOYF
0nxqN70bksaIr8QaCDkU4MrDxCw32aOFT6FA4OWhv7xBBZGNPovfGCsXiSJWNbZMwiszWLupO3K8
jIdmxEXV3HrTCi/Mqg/zL5NdOug5yDNYbVYH4YcNWSoL2yGBM2Vu7hJyH13X6SNlouv74fyIaBlJ
AnO2njGMMm+AnIO1UA48FdR5fjWGXMrUHB/BOKk0YAfl5QpbPi89jb8UhTp0DHzMh1tWxywPtH36
zE3A5KEpcoWsc4nWk/phaoadrA0TWbTZR0rF4VrIeiI4L9qa80RUB6O0Y361nNultfR37p0TzoF4
nkhJrBS98lhuZs0UtXgwR940rnAoImYRhCsgGclPok34XnY+KCMs23TRozs1I+PlNHQEHpWT9g+l
Cgfo2Vnmg096rk95KD5F/HbKjbv6nKolRDoTQsbytEFLnLzGfl0fDL0mALk0cFgIzAM+VN+c/qiR
0tfhrEWyKN3hg1qxPbJ4qVdrQb/MXU1oEtrs9fzaeo1NnpsUMh7MRxIVdJKqY+KLGN79t0Jf7FpQ
S7KNNd3mbhdiTfL4vV6fGKEdH+CJEkAAWf4SDicX17ZAJHKoKwj005J56+xON9HGrDBgVSqpy//0
i0FUHYZWr296xnePkuXaTLYeKrlnvjAhO9Ar5zhtsu7RHl39uK37kzNy3cuK66rzEmpj5VnkbkSD
fhPZUvCCcRzgLZVq5gHTwd4GNeD5Fh8nBKwcfYFfb+JLgbs2sI5FmYXim1FC32Kn21W0TVv5+ecs
i5tFekvVL3jjpmclDJczu8pdblitR1c0pWTW5vbG80mohqK98xR8t7KcYe/tRzQQ5lb2yI+J9B6+
uR5lsNQSGcDnppbiiBhh2MUGXR318MP+Fgxi/CsWAyrpL4lk3gUWoIroewxv7Pqat0qIbvJBzD3w
+lSJsbVRcwI+WqLzpZsFdcIe+zjG75L2y0R+Sk/Cnmb6tXYGq42I9BKwSETgPjTymZl7Nqs60PhT
IityCZhOAvpOZe54mV2JO96DF1n7HCYo2VHuK6D1v9FTCZmObQh7hlHJhXUWURprcSH/f58NZc7z
7R9Xx+RL3eQoJuWUn0Nsi1sJ1PTL/UfB7G+a5M61j91Iwpo9Bej6hQYzZSJ7K+Nrrk1+6IgHZ7D2
cgys+54HReNNWMBs0SOkwkSBehjSAz2C5AmsNNx30LgQlbynn2NSaMDcaf3zrfTKdnafFzq30460
qNiURxjoBznd/8htlUOm1SfsDklthDmdso27nwKhpeYAP7ThmlcAopW0iA9zt3ksMezIv+2oFZ6k
QLLq8GXwrqpJ+HME4Ndt6LaAmKZt/o49/kHi7NvWAsDRNS77JD2IAdsKxkkSRIfNd9AT4OjCpe87
JR88Zgo3IqMaFbATr2Z4FoX3g7/bHWMaKYj3KG4XFmvvd6PdnoeMhISx7GiVZZcBmQ9f/syX155o
Ki0sGzHD2R/hLRVt9FPNye0B+9ylWpyfWARNeD9wvdMVUCs23E50QZGJFwZ0YMcRd4EDmFSLeaDp
EW38JIZQ55zy4B7Bst4/IY2O0gGbzm4KaQc1r4zgiAOuxR9xJWATOTCAgRnUE97+YH/IzXxpFgzD
jjwm9KQsRUt/JQPy9C94OVQHa2CLhZh2byXbmQ3nb/6UVSZimrimSuGmOD+y+/6MMUKHwAajxTTl
Vs0B2oDFfjKdbPRYgZKtgn5Kk5X/t6x1WoR32ndD65448wiRajVyMKc82UQdRmfTIxfAc36JoL8j
5Xl81gq1zsdXqlmPhaswMSgsMr57s664W5t4QyXJTb7GIoRKgNcYDTar58lkBU0UXLYxO7yEWYtM
aJlG0cmRFGTir5qIT4fkXOcF6J8bnL6VpQo0TwrBg2kRhjUs8ymvAV8jsOXLWKRmm6Zh5Kfgy/bH
dbi4oMZYWF3x8w2D8/waE5b5jKiayJ3O/TunFtO1XMc6sX8ZhyCXtOIivpJ1REiTF+Xf0FWQhGCI
VTKuSzBdnzaBbQcpEUf8Z9iniCNlH9JXkXA4d6wk8I6ju8AEbsP94Zqu3Rn4WOzre4YxNybs+hFv
KmHjV6ufjj9XLFJVqN4PvazGB0frb1O3iAQpvlYJYB+6Iq0XUL0+xm9S9jI/sR/SmzQZ5f9s4W3j
1jKw6E9T+8f/SSE2pVNF623Icm+vLjqA/ia8gOOjsxwcMfXSfMcoCzepRL1t2Zb8dWbqsGr7tAHF
JWlPYGhIzA1blkKytkbFmJTOtX/2fvdYT6mzAlODhtmBBDBpDXa9t1V5KLEyE6oqPzjMeFPMsVJe
S9wsVB33V0d4m1XjZ3HjZ42k3XNB3y5VbOi7PgkTf/xPyXSB8AydtIqds2rPxuIEBDRr9EfGpjso
DKF+rWodAQVFvx1umONg2AfXMc97jDMsztr7WvWPj40sHJF26lLJTruhcirwMToYQkBpVaceDWwT
FOYmR18kdUe0y1GoFzPf9i+73CjA+K8T1/yhsMHG+XIunPK0AISEk/S6h53aWKUMRYMnnKeOaQ5o
TAPo5du8hgI/kygEPsyzhQARSJis52gzTlVFOHqj2rkzS91MaXPqi9EwGbLL22Q2vw4aW3PdPJtR
tVc+ep+KXzQoIERwhiA0GchLeWI/2BMAEtR/9V/W0ocJ+nxKBwv7gOaQBMoq9wDGiBuDrk2n8Pj6
TtCOs40KujTPBZUvghd5lfIuwsGhNJemXg4Xut9CmwCt4ke6PEQi6CAUu4XD2djR9Anhj6plPR6M
QeTS2nlSHqiEmxfjrddz3jnFsra/c7Nkhamk3dvDrGmgk3Kcm50obSHwdQ0AjUvtQDhdUmp70Rnn
M6Ogs2BFu68eiAjhEDIYHomeyLXQfoAH1dneDnc1sSbYGBWdtQrsbmlpTM1nn1Kt71RcbWX37p7U
Elw4EJy8uEgn9WUt4/y6EUf2KviL3yYj1nxxFbvXZfIHkBWf5Hysn7HNKKGYa9hnjQ1cKekAZO+b
vjjobSOY3/GSx6/s2uuBwUGXo0Tn/gEMoPSpT+/6/bxhAGv8mOgUJ6R5tLE99L87kXlkix4tPDFB
R+LtxXgh+Tyxy4jM41j2KtP+EfwblxHp7eHVR4exlCdDwyi/YMxLw4b55P2gm2H0uP8kiSG1Kazs
UoGi/KU32iXHnn8RPwutW3sPy2ZU2sxQhG3WW3b7eUSHLdd4bOR6AKSL8d4HWlvSYZYQBATWYaWi
uPfbypJKy2fFEW1gD5LVs0m99UEEse5l+WEQvWM7d1195NNGnNRFod85163oCRgvsdvQbN39gCn0
DaCbkTbrRzM4XhrJv47uv5PRwlO2OOjXTQidlqwYkKgSF/mcxmaGnYHe9gidl9QUXCswyJojaU9z
p3m7XXkFrZ8R1lFCl3z4lnTTeMTq3ojNRfAa+Fj8A1fqlN1rZ0tjoqsuLf/7SWiKKI+GFc63z519
ZlZArhXta93GQGHjluL6GbpQ7z1+YY+PQCvbYKzToK4T7/AY198sy4Qbc/0Qa1pppxQwcznC5hWj
vAu6y8QBnStH8yYtPTJXn4Kt3fPZIAtpNzXHwsI8yzT3a6NbuzHrIr7Tn8s/hdJl4yNakEJsgder
LLy5n6BWc5r5OGHlP0QNLKIsnrDzqBbXbaacE9oSF6xRw1zojkejOha8AKY8OGEkor9feBs2bM2w
RIrUOXak1NilTg+d/NK7qT7fHSNP8hyQGNWMMJdxxngffJsn/ZoQ5/CQWkplbkc/gAXshefXXV6i
LK6Qpu8v70/z0M1uvXmCLcctLvBJj+nFp27VQ4pwwh+seNui5O+eCWU8VDzHtloDiNSWXjef1JlE
MJyzbOD34bTq1qR9wDmLFmDQgLXwGiwETFCqnAcbSpkN/DpgHNa0r4RDZTAXm9YbbLGBCiGiwzkO
ZSYsRMBTeP+c3je0HRgacI3iSfpV6LkWIZTzdWSMCCLtjl59gcKPxKeADNGQm4WUaT+qagrYWoTv
SdAdCxrswiHqVyj15V1FarONE9/+1Nl03zTQjm+f5IpfyP3jVRPR+AR4AxlLrjzZMlRiIhwLV/wr
6ay2AjVMpn97fL3fUUGaJ1myiTumZioA+6tgpL/o1KmeEY/7UBhB/xcabBN3iKik1mpPsgvey87h
g5P95wwctMXkXdYbUn/OeRZAjjNgLdjoTQg0XuBhaZkZQvcvwF+ijlYctkhQu3mD8LdWXfrRyhlZ
ltQYGRpghx1jAIUEjYa50indgVRCsTLqQSCw+4qcedxat1VL+bpxKL/k/3VYE4NRob/xM15URB1r
wdh/rpqpmLNMgzgqeYVzs5nAhG4NgIcwJlfJRZCOfnf866CPjuzadVBURvd7jkO1pITGHOC5q1Wv
gewMXPOIZkik4OxQ3DENPeJEqKfSAJGtovSd9u8zfdX3io7gzwCyWS3+23rE+bbPkoJTlOpsBU99
ICL33Oh/IkIVH0YrAaQj0W1XpixBOt2cuwnODCSgsvFuyZuB3H6IP/Fam7W07akCzwaBSsVI8uIH
NYhThVi29DQ2YCZaU2KAUaeRI6oaTux17D/RY0H14rr3yRL71OezUaobfy7Mj9p08Uz78l1GOio+
CjdxgNkIUUfbiWOMp3StQZ2tNPzAV6JDjce4UpKgv6BC91sy2P1kvfMAoGQUFNvj7djxCL4w7dpK
WnEBSoRoTpoP/xD+2D7K9M9fwoHMEC0uSnjmYZx7qCxQNXOETCrLSNt2yUYsfhFjQLj78fs2DClC
Mow8u7vhRa7jJSuzm0wqBkDiZY/KvGyl4V0bwO0UsNm/uCPr9Iml+z+V4vqPtaWgcqmOvhJ0Js8m
yQr+xgbk090H1jpX6Z/hvTkdFHgkJBthTICTsjBYnpErkwAf1+9VyLatOHVPgtnOsznhh4QiMR90
zamAXCpjfHViETukGb3cegVQ6pwwyWAFOoAJupjxy9dYN7QVpW28w1wCfsdm9hna0eQLQzb6xYOn
ncMj+Yym1omTIvV+t9g9w7NjwtbdfrQl1moeHeaGSd8E+9l1L2ygvApyZZWgWJc/EwhNVIzaCc8F
ZLc0JWwjPulzuxaYuTtPIHpfhxPCxfXRYMpBGWvzxX+3BAbPkK19lDsQvX1RCvc2Li4LsJALdZ+L
jkyQG+J4cFUyUwuzBGBF3XdkIUUoJxbwfspYr5WVQ5W3wktenp0i550nhz5+ON8l275YGj1Rzrpo
5rGnnbudQ5G7e4hU0v5ldK622THWEDCZj5uelGChZjyMSZtzK6offfUDfoeoYZ+unLzV6SawDeNg
Z5q4j6VJJQ4Oysu8NQT0LszadCNo9mgaGrjopJ6jePMYOhoLZPjpU/ne41+So6i1PC+eqyvr0Tcn
4cfSx5TyjN5caNfG0emTIDUeU/7EDWKKSWZxLNBbIlUXH3UtH1Vlh+hzH03sTvWNDHt4eKmb5/Pn
3LTywtyLRbGxsXWfxbkjlE4kKWEF4uPZt0D6DCBSI2LW0Vwd9M2b8b7MnYhjFOWJBZRZ6G9od9pU
zZghrHUETotno+NXEGsWERFE2cR4zyeVnXSXq/9UxxZTjnaTWDHlDHWMekbILX6enV00MErBAt0M
ra/QxO6xzLsnD3OYgBQYXHCgFu+0JCVOqnE3f1hWIjQkZo88St/l34P0nJAhd9PCUiwNWAk1QRW2
KpAyNCHZw1544FYMfPtNQ67iumG8w5SRiT35i4bMjED9zsfdafNuicMtTg7FztowNwAZkMaNEGq+
dHDinQ41CRylceUxHHaEV7rFjhN9R4Of1LmhQ4qVtHx3h0D3ymijFdjZvwP0/6LP6MzL1D8OQgGX
D6eQWohT2M8eQzJ1pdjMEg1QhMP/MWSEI3nq7EYYeTcO51aFByWJ1crbqTXp3wZuiDUdrXVisOwi
TA3Rs0v276H1xMrTpB2OZrcaJin9OP5II7vMuIh7HVEmy+qK0Fc8zUAlZPxDz47dGpaLKbjjoiCs
VHAhhNdnfWbqVvHcNrnFBFhgB3zlG/SRROEbImJ33Oljspcu5AHcUajk2DVQ+OjpfhcsAy4Oxx3j
CfyEkevX0fLs3/AZpnkXoLdsxvwUXtProDkD4un25YNz9X6Demi7G/1Th7TMbo5MCvQ5XmsJrjTr
3TQ0/aMkLNKZuvzmPhr+kqfuRPWm/D/GVpRRkclMyDTu3zy8Iex8bxO8tt2iNr8G3FkphZYaBT4Y
aHUUkSbsf83KV7VzcHcjOjkDOwT/s5UlQOvXGH0FffSQtsFq3+J4e24FSHIYCZ3AHfhnwxhTKLd6
2pMmMnMe2yy/XTLX/vzh3wpaOEuAZYiXsLL/wxj5zfz+DJ9//fyP5sd28zYo/nn42aqniC28KJMp
Z5CVnFRYwUIKS7gtO8xUZq/unMvo+U8Z0n015LBoftNCSDrgWwrwP7i6nmVtyJ4bYqXSftDjFHdt
+O5+O6ePtgoaRty9Du2YserAIm/MS/yvsl35P/mVjNLuS5w/AYTR8n6+g0epBE0Kk2j5NFlQeDA/
kxP677L3CJun/U3fUIY2fxMaLdCkm0tIjIsix0cWTNSD7FH9yXwsxbGDTGYeP1hJ3aEAcBolpX7k
fjwlbcYURCIFiBh1aGTLdLAhecNRKzIAy4tB8YHC8t34hmRWbcb3zkRPWWs+rsHXaWYJF8oqFX+g
7wJjggteQtJ9E/X5kkeW69lR7bN3eGl2umI3OLAzjivXLu5oKUk42tULGWTi6WhAiU5aFhP+JsN2
uC0tRtP3BSbtNj1ggh0jMoK52CmeVveVcALiJIN3cgzNWlo36BuZWdqkmWT2ZdKCO5Ct5RXumrX9
J4asJJDTQVpFHhVUYOodkRAkzo+8WTJj7ZT4MDHQsVQAMWVI3f76lkkDfWUizgRYKV308hIYMv5U
Yx4pVva1f8gWcuuI81iD/PzhVz5GsgfdMhDzua0vEkAPZsBPyaa1k0qdY8seXmUhMKZx6iFKczQ3
QKFrxk8yVUT51824Coocxo1almdCAxIgZx79rKvvsVKgq62XRxz7+GJKfU5kLjtl56gJAyFIE7Hh
6fJsTQ8WloUcA80Ta/0/lhXE5GCMP4Roxi5jLuTBE3No047bnbGkyk32WTMpBiRyZY9OrEtRvAJo
8w0wFz5n/FYNcDpPRKYzSaQ1MFsyUG3sOrS3wI2jdxV/sg9Bly+3ibymIuTc8ooqfrDw4NBYq/yK
Omok1L0AEa0eN6iVlh3hbdkepIfQ+xO7qQcJOeTwkj4T1F6QDW3lyLXYcJL+Zu4h7QcMFp0rjMQV
qSvfu+1TIpZP1na9h8BZ8LR48mxdegiwOLGe089bjBptlq+eMtkW3x4EZfwfPaZbeuIY+pna78yc
g7H2X3LJd4mRUlgg37rXoVkKyIyUWuPdTFYHVQb7B6B6x66TqOjxqlowGhUmWP3RbAt9zNaIgq95
KZUeDcxeCRlOtuJWjauzwJl4A6/1Nx9mDwQSqa0v0AUmLThxAWOcjqrkIFaPXOqrCBKKEfhFouqg
up145Q3X2hcQQJJihd6AX5n2NRRvz+XMt+Hnz4ME+H22XA1FHoDOG7J/ylPeNSafMWLOQzVxyG1I
gfQUT1IiW/1SCIiDVrR9jRjawHt1TlGGkYaHbM//g8dlY9rTvk8qWRxoX+EDaCX22nLXu0i+fFXx
AZ8nH4yxHUoiA9iqglM9YMHj0UmpdXUJbJR0eN1alXHV+4RpxwoCNsRUiYF3PO+lGHk6ca+nocKc
tulg0wFcdHZf34pelTCEYbB/VWCN1lDzwLatRoF3Ug/Ga6PqJmUatAjo6vw8/UTB/7T1QecCX5uE
/OY0VVAfRHPhZcpQsNOIDJZl0YkgBWB423LHvE2SeAn8grklMFOLRzMUw+pnL8S8sAOwWLQwIYh7
KnSVaem3NkRboiicaIc5ZDjIIqgNtd6AJlXC2TSi/2f8JQ9IBCo3kjqIgboMoC/iLkUWv0AUXg7Q
RreWZ+plT095avtSIpaY0WS+NJo0BfdE/b5OJuFgmM2uP9AQloZu0DLNP+bbutxucXLxIrKs55gF
K3yy4G4LInB6G9oJL58wZPug/sh3BAfkjDt4XwgO3rRzXgn3EblgOh9mYw5Zi9sCpaPP9AA2tGDe
MrYbhacBsykd24UbpoKdAooUT4SgaHNDxNyy3J7d4nqetpQq0BNgYdvOTDSGLvEsfRdGO5y0jsAL
uQA41ftOtMY0O5vbCWQLo6IIhml1zu8WwAePxycERT+vMmnWmiN0VV5KN7anODe4jMKpahQ9y1JH
6CNcEk8DgDxMnlbSY8SHmKxDG4bFg4lZmFR0Hxp1OB5PvXyBBzi8GYCfPCJ6JSC1vzSzD6KQm12B
7mcl/YWT5vSTs6K7gLu0ClQNcvYeOh/X4bRFBgXo3aAqk5YPSpqagQM6mOgox+1yOBrT4V1eQGtQ
eLrwdBWk7xYu/Nh0mFFuz+N/0tkgm+SAN1yvxZELmUdO4JyiGF2/MK/7eeTmyPfLNXTYx8AEEH+q
7h51UIXL3d0x18N3W40PL5A7Uv9SJlCEHIKY+T11mf8gQmaVlf3+WQymad5xD8fMdNVOwyhRUx5u
hqbEweUZmA2JBn+bqkMl8RSPacvUYuALJCN6VqIpUjTovKu+zaWAV/k/GmRz9mLHYbBOfsyQg2Pg
r7zC/JAScBg07/i5AfJWQYigXIXYJrd3t4VVP+CXoIXNyQnTHvCF9A0DWeR995r3JcP7L/68Drm3
qx1xOgqtWy56k0PoZyPJeRnpUNI0WgBXMYPLEH0tg32+7+YLM7DM4Tn5pi021Y0BZOQEVRGCeQkW
UF53ZzuR8wtNhSfQD5s/4zva9fwcjLVTi8XnGxcgefN4XmL3pbPh9EjdQ+GkwIHb2MJN/xIpXHbw
amTNxmHT91KcjraRAB/Zw2vr48KbwwSrcPuDvULm5LwS0rkbui1Olt/akaC3HuFHd2iz2w/ZUuR+
uaW+nRXqrRVCIdV8vsPwVV7ffJlkI/OjwSG4I6IQbMfxadrNOqF95Iwo0sGxzV+xaVjaRUJjVZbL
nPgH+AzCWKay/YP4e7XNNEXVPm7JjEIvNIdQhdoElhegC2b//fbXXHVu+4HQSzqXpwI5g+osF9IV
7wfmK6H1zO+Dg9/AKC8uJuRPasUzwu/SNlIt9/Xv/fihYblS7CE6jEZ4hT47Jy1/i9OVGNtfqI/r
XeLcTRH589P2sVQoXWCCTO67+l2xpmQyLxP+T4+V7UitehLtziwYaJ+An4IAqnmbkPXxaaM098vb
SSC3/3TgHvCnNkpvhBPvgo3wjpWiAwPCGNGwTcIoPZGTiNeCbv43GesVjG2SPqDST1W61Xu120ha
PiDKYhtQLcUxsOaWrPuHpIG/hGLt6P2sFz0/aEwcFcFKceL4sv4SHiFqyh1GPONckc6quB6gPgF3
NTTVNdVHB+qOcy27PoWxQGe7sP3EnNR14THMxrIGt0VA/1BfuGjQ/HuTtUPD2aSFYapf0MzuCfBB
SKYm4gQpZfHNs6UTtjxa3Abh9/ac2Nru1iO7Fu36+vIAIOyuEE8o+elQaoKfjSYrYHLnxFCHyOyY
XmcJPa89SUbv7M6H0tQ2vCQf5k8HmuaIkqfbWIimdFPw7dIXi1la1zbdgBdqQWIbvYgu/pk5y5AS
WYKBzl0S27QN6tV4GA06QJzGHfhsHDbMhpl57j9fAI8Y1F5JZF9Ay4M9f3n9XmgobHaPWPHxjdwM
Qg0EqKyK1sDvH7YppKHKNNCul7dKNIyuiNi6wNeIUDeHTCIEjp2IKwRks8sxnXLNODDXN4/5Ynak
GJzR3PHwxzzzCgKdNh6kmA7Y603QJn1TA0NKsma/Al4O9fvK6xwsQaQnqvcbzsTjsbCVACWXelit
5eiBcdAANya1Ntz98vE3L5axJaB+c68LwNZKBBvmFW+JY1iQp5t3eRKFMCgII7C+cUuFgE0yA9Hy
npFZCiLbJirYcPfC3bCQJeMNKPiX8NOjKXxG+V04uFWmISQP88lYWovMHbo7dDQ4q5bKw/vAYS73
dzbd+igWtxjDh6Nszb0MK3OnVAOKNSsFDn67a+gzkfB8BsDDtv1ICQEav5UQAgEFuVvoRHisSUtq
us6gl7zkwYDYrwLk0C0MC6cLezE+1Til+iWh/t47DFF1TxDSN04OCmxjOmkAWtVqcGTWU/fmaupE
n424HYKvaNbGDemBSN6g0NN5MsOvOH5AH4agSbENm8oT7ZcL94bjcu0J/LZttcUvPhL9n4j1sJRf
p/cEsOowoOZ47/JvgGmK8/J+MEYaJAMao/8Qp5ZGCFUOEOxX/xUJUX9xab8byKyIgFeZm+V2SFYh
dVYQoTChOGhO9ks5YKTNpiH8O44asoV7isAQhpjU/fotKVy27HGWzNIwMB6dYEBZKEgyZGlrkI+I
d9PMfHZM23XqA9/rUQp/e3iMlAU/SMcVxBz99sitjOSGXifb447Vu248uvCHEQro+Z7ycD2yVXFf
hu8Y5gyJt8NgO2OSru2paZfw9i4J2NISPctI5UuRep5GUnmeMv+3zURIbhI/xJsARCRKO3NxLypc
NyF/d388gehWxpqM5t/SXAixLLmbcYT066bdz0JEfpAyECFEpIkklhTlBCtZahplatvuitQudalr
Ny8a9oUyXTIwXUiAzZjWPie9oeWiCaWb2L497NdfNyGeVgLcethtoDZy5I1Hz3hdGPvqkdVP4dbk
Bs8v0XtT3z1L3FYg0GBnpGbBQMtURyoB4D8kzMGVvps0z6KqQcu+RRg9vjxT5zNDMsUfZ4tlT3Yg
qfD7uDR+uO/8W1f74w5oWo9zFtheab1Ab/QLwZHLXNhhHFfnsjiSed1tYwO+SGsI19dvYOAoFniV
BTUCWgWnhZHUR7vBu6A1V2hObCKBOmaK8EUGZNolr6t/uvquxVIKREtbit95D6KyMk87MIewz6of
nGOTIT3KOiw8EZlbl4xvTSq3aq+eJhCmlOUtTMun7p+gSewL6GNNCdhH3C8JMsMF/z5TU93lwu3r
8zatTz1s31AHor42AYL7uBGX0NRYqRRcn/gWS60iMws0oGO27oihJ3jSb17LLfpYG0TB2Sj6l+K2
wrBmz+FL3F+MMVCXXuARdiALOrHAircjUMN2s439pDbMsqpyzsI/zoBipa/qqVg7s6sT7WP2EDYh
Zk6ubxbSBs5bkkLHXRuf65zqS7ePPgVfc2QwUbbeX3RzeK8EWNr7zr7W82qDBYq0Ls/MoRyNNidb
G5O3mlOyppshtOQFsDDL59XGRbrYyUN4gLMAMICvskFd8aaZ28+sUN7hZBwHSV61GkPtSIILXDuy
NEJa7Eg/ZWNFopA0UthHXSBz7w70Mm9dgvhLHL5rXXZMnWKN1AbDj6RzzBfyxBev1ZFY0oUCJ3DY
2Je0M37dcN9e6YflV1XOOE7yq/geWCvybRAXAltXeWq+GIH3IMk3RgRTp6bbI3mdUoEOomHOvK/b
NEVF5rCZMpYf9iUSS+XYBqNgsNMxRs/L4llwy0Gt+IERLCq2Xd/aHaS0ASNsoOJ7KQQthnqzf+TE
+gpbTHYc+g44iomu6Zww9TkkluO/swcWEBn3/YBbqHIG1B0TENt1x89E/xRBN+agky6A28syAayL
dbPuTKACVLOpuGKz/Him5Do1hLk1wFdDccUDEzYhaMBTZS75gkwl+M1McR76JSYXFtfBqapfkzCK
A08Mpur7SZSr7mtRb5BjMoVs7uptfUgjOBtKDJeEf+2z4sIDQZSgOBS56qI33k6CzthCV8K1kzjF
hTpehP+yxTanvZ/XXNl2MGzWRGSEvaVM87nF0/fSAC7nfQMXVc69sMkMYAcL8pf4Wycm3/er4QRo
wejjuDsGurruoxHlKNAAPDgqc1dXxgRzS72UAZUdnv1J10Pvp16XQnwFWAnmhXXZMvZWFzWmhvyW
ZKLHV9aidAIQboFeMGqmGns3t/QC9gLzbQUqoUtlvAUEBHFwrkDIhTZe7PHptCWTVVRtxfQPplwi
lr+M2C8oBcO5gVLeCdxb03yit+hGtyEzF2DBIz9ssSyfJy83lJ6WGXwLg2/h7SdSVrtUz3N/oQ7C
ru25CBdWE8U5aBpN3oe1pwLOUNmKeHfcpy+AGnF5ov/qU/YW9g3/PEd65lowxGqsoJgvslNN1PbW
EvfdujkmS9b+y+KcQ+2VgIEg8/7mUXRBcuRglm850G9My397IZq2hl+mrewwk7mtB7jnN3V4jycs
2fwy/WHQ8C50uCOoGq/pt/VMy6TGadLVVaHv7O5zbGg1g95Ef7sZvfNaLEgF+ELKMy/3sbzhP5jx
WFDTPe84TT9fDSCjO039Dgn+NWe/lFdOI/Ew5PqncY9FnpX5GOZexi3k0db47vs/GjKX/OQB5Pgn
Nj7JDbJzgAWdAhRMTpv+rTTGMQJr/gkcRl/bqLlRwLHLniJ+t2n9mttWfsciO20eNTCAV6s6b+Sh
XXRkLJKlTZ2r+89aVNbkzLLpN9wWQkHGn4CD7+jNSvNPNws9ETvuJHBGvYT7UaSAzYeID0s2SSeq
UVyowywsokIqwqN6jgNgAxbABx14YhDMvHPZlsVt83nrlp703bXlN73j+n3Tw3D7h7XP0NVgpAy1
JwNuuFFfHQmr6B3osf+iWfufDVTBbJYWb7ZWtF7Ziuvp3yw3N1dpwe8UAIbMSUjcwxBLoOnpD6Jt
HGInmB3hELVXMA4Mw3GNlcIOh5oD2Slvf+rckOQzqJ/r4NQcFVVdZiRsbxLw3Mb292HKWzJPf6VR
7y6KeObH/xpb8ExpmOMD4U0Mh6WGcZOnyCrn04YP6NdeQjxLPqFaiA5Dp/d+b7S0c1OPWytmp3BL
BMB9+3jpqJTCeuCQVurc/BUhQmgh9cZW6thUohQyDfWOEhVdcJ4s2isPIZYIHYYKBxATyB+jiEf1
NQBx0EUeUC+x6ZtHgYsl4RM0viMeNJsRNOpYAZWORVXSysoobXKL7qrYHmFXJlgvC/J1d2G7l6Cv
kfmwCtQCanIGBeSReU02Yn/X7j1rMpcKkW1vNp2IH2B44k47usQZYvLt1B5g/bG5gNisu7mZyIIx
dT1SbvUu3WNwDe7rA8cdRkC7PDdjEOj7nliBBwyeqAADPZK3w15vH7JR6dX3I3HLludhQGi00xo2
MjpXsBwYzEUROWzXAnAH9dswfhhu/MGYg1vgAGVZx2gijestmoXoGs/gaFXHPktuJGWqQMtOdt4G
47VjFjMcj4saK1xQVkxbIco0madCSEx6ynzjVjFAys+IUxJPs68mkempFFdSFAURnKcjK2W8lbyY
3EA4ooBgTtklkfIqv0TvyVYxeSKWvZz3Uli4TwYVdHi2WZfjz56C+kepLT9FIX51B4FsIUEGzlrX
+R8qJQ9eKBgJaspl0pKRa1CDt0V9XRNLj1JrlbagzObhjsy8D78zS2cq8pyFgnUqGiNeoROH0DIm
Ja5N52ppzz+nZkR5a1aO4ricixBi056rQt03D4RoyhoS7Y7cknx/CLFnrFYLjk/mUaojAGZxBfWE
vQQUtDrBt8SgtyEPFRV9pnRBHTzJMIF7u8oZgB2x27BfyL3S1Sa67E1DWudYcyXzPXnJ1nFCVdXG
V4Al7vwjbcWtg8iOsyJzbzNKjo83sugtiDD4vxDVrOTfPK7HlhDgAdE195FgoZJPgWOsJ0QUBU2X
a45tVRkAV8I29ETbSm4w0sjNpY8Ss7dsiupnaYAkOZF//7oLgXvLsbVtmHtIqvLf5+LQ7S20SG0H
0J9kEkO+VYyKztUlRDJoxBc4tl1UgAmwqK9sUa5uKFhNBbU3bQw1WnIsnkCu7ZWjGkdPI+2mEXOB
smYxweHGDDApEA5zzejKcg0wNn3Cm/lWVRFCWzpULsCvYYVuGuLo17SHExgNp5z1Tist5SVGArtm
fLJiK7DdLDOL1+sYGH7rb3LyuqBNhYO6v75OssQs7DtP96pCnIdk3ER2eDmSoy8XuN+fMrtWMp0u
J2GnCWpdqXn0pDzGWZbywJ0sXzeNt2GJDb1016EeNAKYXuugMndPxdBxHPT0zSfJQM3HQmQAWbjs
VtmPe8VxbMcnw1ThDLonSTvIawaZUOl7C/IQqY3G9y7LI+4lNyblRs3SxI1cdiEpNba1JDY4XwLd
2+xhy36ppuIhUQGkEXJPp3r1iEfDs+DNdZki9Y8UpSrnFpHyPIXwmQODLY+aCBh0btEcw680ahOe
jkbSmRklVcb9wVe/vnsK14RypVm6ehEdPgTMFjESriSKv+FlneDXg40VJv9t36GkzNrr30NkDojF
xtioB/Bzst75qyhqKNXBW5Bc2NgqpUc/ggG2WJtG5/QTEAQtKFsTauIUBlY8fzp63WXQehU8l0vU
ufCGUVQdluwGhcbMS1Yv09eP99CDnBADIHB4PU/a8vz2YqSxoL9ECl1vCJm6pQTNreUQU2rs8niW
lTYzFFqR8sGQ6oAiVLx83mQ6OJnZZhIjmAHEEsUIBNLetC45E6YuHygr1diI1QzNKbZ8LZjjy2wv
zDhQgNg//WgKyUhcLqYhDI5xhUHxGwdGxkLOI/tkvbU6Lvnfp3NnIIaDZnvbh3TnjHvrkASSIblm
QE7g3JrxG9VjNhtO6+Un4NB/jQGT+NAJ/3Pf4wnbtE3FujCJBh/sBCt7CzQ7iLCLNsAPv5NNzu8J
YuyGg5O9DoJg5l6mrnambjgtRKKkuIyK73gx27ZB9gsx1HmSyMf8KA8uWtaOIptEMDjums+56skv
xRRhMmk4re7tVpAm5CNTjTVggqnryIK3uFTdJfAiSDKpd3WpzxQjhIvsXwEBVjls7Z7K5rO8SKOu
qkSePIr35Pqz0WUjujQV918z+gY3P/9Xa1sm7DwitNR+plnHdfLbALqOd6Fru3qbP5uoMovSHhM2
lpE2ODVxbA6aIWA/B0oKp5J7RU7OBjLksg+mmvmNAHYCNC0FIATtkO1WwoxLIROp9rro2kw1cFjN
rQUbSiH8Cvv48A0LSsRk5XQv45HeLGL4SaMXgvNsGKobaiAdR8KA0pkyWtABgXpQTLG8LVeVw1EJ
Wmutc38KwksEOaImFASJUjM60BFVZ2jAv4i4gwlf3qqoJvXJxVON6vkhTJoqPm4NpJ1zsIkKAk6S
8WgHGNNoN4brjUabuSPx88HLjgt7L9d0WWw6Z9rEn+Fpt4XJgM/CASWzuHbrzKfE0LRga5NOxe4q
kC2ZRgf7ae3joKjNPerThpHlkEPRaPtM3N1yppJ133XWTmVVnsrh8MZGzfyzUWWgkiNaq18w5tSy
RySAT2EzD5/ek7clSdr0ZRtwPlRJluIJtPHhZdPWEEdobKIoLuRS+jInnS0SJs/I0InzZlXg8SnZ
QVouQvH1xutDja3sUN5spQHbtHvpQi+eLwcmHHYclfUvsFjxO5NRdCJkDSwAYzGUb6I9fn+gE70Y
jv3lH9M6O9LNgZKjBbOKg6XbL446LfXcApjSi6jt+lOPWDtoXbwkfleDzm+1oCLk4bCsEZTtD70b
1K5eK1leOLsrvb1Pl50b58BHegBb2U7yk/XC7LdUsQwre2bbIMKqi+vMkOZgp610cmGcV2QgUk2r
ok5HDoGMko0gwxSWpRs1yZMoHTrI00Krza4ysOdjg08Mxl3qkRmrxkGh2h4cf6+SpIDp21aIuvdJ
A+WwcAiS5sRNSv88GZy30Ub7rjSW79qGp7UE+ITTeGhF2dgcMrLcn4pV+Egj9SlaEfBMwNKVBDv+
QtyZQyyHCeifhs0TdDPQ/Ml8ySZMKel+D6HJqOHSvDMiSKo+1apVJXtU7X0M1S3AZzHY/LNOWE0q
3R9bsDIqg/eGdH5ZgpvxkMz/c4v9+KQ/Tkne2dIfNYTvwvsRwcR+0l3m8GOfjAu61o4RfNI1ukZa
xPuleyMHY+kM1TPS/Qt16uhjsg+abVICzdvylEPQ+5bDrPQf/pZqsbbwoLvy7G0f8GjA+gvuTx3U
OABfjRaa/or9M+T3cGMFd03ffb4X6Mv9jjyXb9EPMbPcyP4OjKCJi87l60arqBEvvNpeggpL4c8p
o2AnR7BtRFaiDrnR+7iIUnVYjCgCae1uOz0IRY39ZObj6P51n42gvqr39siRB1SbsknBvrvje78X
s3REbditqLyUGYex3x68yr2ME25j0HoeQOBcTc8oJZfwwZfp9M76NQCrTt9nTNrbZy4BZvR6TQVc
zxGWxzxRfvUEhHYBhqRywe0PLDEy+l32qL/v1+t7xJ4I2s0XG7Ekpko8S+kIZqbxf5AnLUiFgfAw
J7Z2XuFSzUnJVwkdT3Bc6bDtNpIxRX/zc6Fr1Q1imgB7mdpY2/lZ1lI+VvnLJABwVWnvF/LOfJKy
pMZM0Pyt/YVchmOZ3cuTQPZ5zaITPlTYSRd2K8WTQj++Gc0ja/G2+8/3pr0NU+g+RNstOaXr2LpM
cBh6jSm+bVAuAaZFKb7aHl33sTqIcgNOpWVi/Oll3q2ZkqeMq3xFVu7XMS9RGnhjwvwxgx0tp+Z+
7zwjTUboyIMq9tYHtxCmUNBMmpDmGfl8GB1tleqQkmqF6d8okulEquAltK5AuVtoiON1ofJmxIcS
ezDHkmcNLHbbrlLZ2ctZt0KWRNCVQhZ3FfyVHVCfAeMvd1u8A5QAuqwy4j8R2/y7aeClucr4TnWj
jNagMZDHZ86RswKD5EGRH/yQ+V3/T16W06/Ynu8ui4dQmcsvJV1WWPdZFm2I11lXOupuqoOCqORm
z/B1EQErwUQQublu9UhzGtnhouhwUYvx8D/1wSnD9y25GMIgO+8dfSyneVdsqQKPLFzvuY6HDvXo
zTXphlTMD+eTt2vSrenOQ4X4mSXrbLuzrhwiI4YZLH16uZXbmFAkXTmcwST/kl/xFpBVjZklO2bF
+IHXjh/igMWfFLGOVbAFVaomnQugxsVr8YE6XMlY2JqReMq5Zfpp3WYp7sTudDdEpBXpb99wI7Qd
DTIBDUBvNBK2OCC/2n642/xy/xqSJ3LU0vQaSmNZbkgE0TEw6TIyMuB3bUV35ysRyJz3jbCfQbvL
+4SzvDh+IrXby2JO+TjYtZK8K1SgCvuzoWmFuDg+G0lVEpSYgP00DWS77F900VnWgsgM3J9dWJDM
c+q1Xv0wQTD2tWrOS5JJNzT/9SsBThFZKHNZHJQIq6js6nH/dThTNIQGn+m6tO0oQi9FxP8Nbf4p
EKmXuu+73O1uT08fubkA10Vgaqe+Jw90awKHqUM34OROilOhP71oXUX050XDGg3UzvPxKTyEORem
0cujlpFLwJKEqFuhrQDfQmdXZd+JSLmN+i46fgLpxN7Mpzog1i0F3xEG1TKD8sQrQU02wt78wLrG
u0h12Wockoj7nBtR4CAjYIPc1rvd/DRNxqdB6KlsrruXZLImJ5nIf4NM5rCzkglmPKPE12Xm1X9i
F729WgKqaHaKQad+Dqm0xx6TCvLXlCMRi81kmpnTn7/CwOa3O4Hw8DbHFrVzBExVIOpabL0ixKQg
8+fdt0ienwX5z2FBTe9gCqysip9WqvAuDyZt8UobtTfC5gGhMdsff0gqFNsyBxslZYcEXxE5qLsJ
jAYNv0s/AndbDBg6djIoY9pr8nyizhgucp6WRjbxb0RLhgm1GJmn0CyFA1UP8X5VmC5dlcf3eqBY
kwEPGeIDP6SKRJRTMq2JZ4Zytqfx0VDL1cYL3qPy/4oE/uKgcZoY7aQFCdmEvEg5aOzyM7GD1iN/
Z9S2P5oRdML+/w3/xouGiRQROlosR5wjANi30C442lZ65zg6FK7BTqZPaRJkI+1gt9VKap/DgBbE
jRnv30C5AAD2Csj4YugBqf2t/094QhoB1q9JhesDvIO8IavpxLJPpO38dVmhOJ6s7FbKeEifvdNn
zpStD5eVy/RAQddZI44xZfVWMb5WfxoQYkpOU/HV2PPVYK24kuy5vI46KEZMCtYXrdn1F0CrP7gU
nGeIkMjxfmWbtEPQHX4oTOktdcw2ieU7qnWwrvOH71psMIbTe9F1hQ2ze4/h4Bkeak3zUZROTRTP
mOOYLNcM97R2gsha7Zn+r6INyegU6E/viuSKOmBSDevaLpLBcs4KKsMhtTsw+UDOYx6vUKbtae1D
5RAz6kz1tZ4RDpn4u9gfEnXnuIEj+fCtNuC3hobYX5mpVawLvcLlD0tvabgUzKiAY3132fyaD+zH
58gTOoek/zGdloKSVpiZIBORwSDdEUrcnEy4alMjcTM+sPxY7o55fOGWft6Xk2VqJwZL+HMPrzVN
MQBhaTSC9tE6jyJHizuEJktqgJkHlDp+IStESaDcDzWBDbtyIT4KXe4wXB0vl4XdnBWFX5XaPzYA
n6K+3XvzZH4ktxkvSHXotd9yECrC/uMmCV5SxLjqonQSSQNYIS2OiGEmynn3ejNOK+7ddVc/VFh2
7Itf12x9pt48dSObrvhVCmyupROBEkkLYUGARZCu7lt/FUeu5lyJQeGpxhSt56R1O0D7Vc94dy+4
bjx7NfQ4PjDNC1BTImIK4Jry9z+INsOkrZf44nzxKeU8PeSLM9NbXgBhMkatKapoHAYvbc4O0Rfg
MrwrZFw+p4IVAsN4DpQQqb0GLGtZsfPrHr2p/TShF6Q026XTuy4KKDuUWOLsJMQLhOFqDuZk/mzK
I5WroiLDCNChkfoIarmvLcahpmWF8f19T4G1dSHYdGr4IlC+cqmA7eevum6X/SP9fzoFBjxJ+D6y
47vDRgp2jIGsReDBvxz4Q/f6m05QE8seOQNu70I+oMaQqfYNVjeTBDuKhog6z7/xTai/KUEkvAlp
JIrxSmsTYtdpEI0kdvnOQmjxl5c4CLma9C9N43+6tncGK5afM1C8DaYpycPEu+cpe0O4//FQGZSz
H45b2EXGzHaQWd/FFJQK+QHf+GGNFxm3OPySChqegHVCdVE1THI4RnHriEKuHX7UUX9xVtAfN4RZ
p335ZBGQ3NIZgQSUU22ldZI2YXrxzqMUpL/TuyaRox5yUA5l6FTxttkx15h7q49lrZXZAWjf0Pxk
RqtT1aqqBgGn3KXDGQRPM0P/iBMPN0u/8bCtff4HuMSLXwS8Yq242Sk9SvNeqZ48mGGnY3nTgq0l
N04hybkrpzEVuPyUhC+Wyd29r/iO7WIgBlPVSh78q7/NI3CEIQLYaTnKdmUXj3U+dJgbc403wkgg
v6PYmCuYzEIBUSU36W5THBfUhTOG9e5HAxBN+MA5BRGvyYX9pfg/WGg//9qBkmIGCeVUiRYctmoH
DYb6v/VofJoPZN2Rkf2z1VXxuSCS3uIGl8UoRD2V/IpKjFmnseKTaONAc5UFFwJ/cPRE+iOxl9in
DmzaV0meZr2bHWAWZUrYF2Indo/1HFbTrMrMV5/8uCVUM8oM4fHTFCucriarvVCc6kMcCpaq2HgW
wV/NkxCcaE5/qtLH8wG2vDLn3wY2jOi04KSJFm/SxcVxUy6SfuROTG8+9XU5zKUJYltFVHy0IPKQ
PaKi90vV2om7AkSykxu5ghwok8DEE0WcBX1OXcmRYQMFTCC/5R11XA7R275daHkOLy8Y1go5cXvh
5ZtVhJJx4Zw1vz71YD7D1womVL0ooXPYVc4rJccdHA2Ydgqqmzoo2FZIP4zSKIeBbtBNswRm52Xc
uSIsv9peiEXgYtXvi7BS/4SWR4kEW8qRWtEnhSH6TcoBhfChR++wBV8qKhh/5DTiwqVrNe+aQvKx
AJOvkWeSknlJi7d3SIxJeepEPON7OPZqHzO35FgN9fAcjRvuumBNu2V72tqEC6kbTTrqWnmRQP6v
kENk5/Elso7MT3KiLkCiF4BwXCxW4ak7MqBF/AIXK4ztDVV6vJg3ccHm/xxnCaRyQncmjBIrFaMf
QoITWyt0IvVrL+MzDwjivwaYuP/3F+S6TSpgyCL/Zkyj7IBSWqEA7Qq95nixPuNoERH13lZCO6ZV
nWQhgOi9pGnduQ7eMX52tyExpjXc+2Vle2Rr7wm2ahbc6Sxrb1qJsXaG+G2so/xztyHVOzmgOjd/
hlt8syA5eiOTC9aKG0cfTc7frV1SwSovyR3bl7C853N7x8/mK0n5fAjVMJODGwHzAg8TiOjJkUQw
/6eI4/U/mxr+g1OBaTAycHh9IydAjMlAOuO/81lgMeGa7Nn+cwoWFVgyXOERslAP62AlcLMGOpq2
lRmRvlMRRpYwoxnR0eTiIiMBuzXlkYxILpUmsXLZ6skMYhfSpxkM4NW16Uhh49bWHSop/ClgPmRO
lc0luwii/jO2AIboMc4HOtbzUQ45AthLJcK8tfGATHAjyrGMQhPkT/elD3k487S9sptc5wEZinZM
luF1GYG8v7CKYbCiCXI+seRIfZrOzwtZJzy8cZ1gAsMjBQRMH0fh7B24/7L1Z2uLc58FKYm4Cn6g
pJ84MU0YCZH6etr5dStXPpXHHhHlvdvEEFUjLZCNawF0Ddi7BqOmSxdJH4qU52ER2sf/WJDTEeCa
aAsGR8M1liDywD8RN9Lg7XDLgY7Uce0g25Xh/3+H6mGAz7BJKfQCxPVSu0yem1QW6Fc8vZ0QTDrd
RfHsFCJKJbVTxCkTA62rHUd1PtpH15lnkLYykqCrJlQUs7WfBDXhFd69jz1uVwS+ERDQI0tw1xCv
YMXa1l/UhZK3bp1P7qooNd8fSgMfrwga7T+l/+T3XtHV57jpRhztvX4Y1jnSFxSvEqFExU8muRPT
dG7cw0n1ueu+ttaeKkGxSZVlkwXLLja1QXMWnOcghFxUTr5n0AEQ+5VtPDfCXj3nDd1qO6N8BLG9
Lk3SeFA0HmVhXL+7BqS/6bdWiyMPYGPMKZcZcJS44F/dvkKK0wqUjEA8HA/y9qWuCOBg4OlDpNVA
vUs6TDJXIEZb2QA+LHHWCTg1ifN0bcd9qYBCdFPsEO+nnc6pFTTp2pXtJdWZg47zKaGuCGrIzBlu
GqB5yS8/7JNkXroxbhScM7DSQNF3Ea2kqURQKe4GHpikKTfOmijS14Vv9I4Zh0Dm5l7fbQcyomYo
vq8CieGKMJl9N1dzHmHkmzlrszmz+FUfVbGq7cpvGJ+2pymYP0pid0OHfChlvUItKC2lXoKlMaYx
p0/NBCCc7hwBkehujX0eLyou0B8lqwjhSN1Gc8pEFVXHmhF60SezUbsHiLzqbu0IFTy+wJGyomqw
th3vhS7FRZkpr9YKwJR0ftyqJxI5Y/eQ7+71jxE34mwyvCr/w/57XFWs7vpvwhSLeo/tRbr9ufdW
cKS/bORFiSIBYOG6wGZL3nfzQSQnyIUdfs8FRPbAIzYxJvrU0AMDav3Q4ndpn7Y2Da22FO4bF+iJ
go/WI2uyUDySeIYLR09ilkyMxp00gumaYM/Ob1DfPYyCbQp3gnHVEEOfwX9+tKNl9jNA5ofIjFkQ
OJGTWeUQvUmj9zhu7Co44cGW9UA8NlG8H2qV5YRAJ4I5wgnaU/1ViRO9eYooLE8/HhmjAaxqnU31
VoiqkmcVe2b97Xih4/1EosxvoGOb3ls/3sgdOHAbaDjRo1M+GSnnd8SaYOOX2l3zdzGKIdvFKAVC
4i5QatvHHQtgx5LrNonnok3fwdzfhNdzIbfw+RIPKkgnAGs+6dz9gb2pNqhw+QT/Avon3ktj23tB
SHtExV/zS17ycFOAFHqqsRZbal3LT1HJssDb155Drmn/jkDCoHYJEK39QvTNEfUnezPKk74hOyfq
Bpe+YTMPfBJGuiIly2uftVoVLMy7CHnTxn5BuEkxZ3GmEqOyT3W770DEcfpkoB1niZQv13IugG1Y
0mEOm8Ha5+KNQWGeyhX9SVW6qMjJ1A/y+sMiiuscmIc1mYjNrIy31qoe3zbJzgbZRl+6wrM66yqs
42g5jTsht5omvXuCGviFG2aQxMMtGnQZYbjaQ+hAi2lXhZE4Pp3oBX4CheEts3fHWrkGQja3YJoi
iyiX7gWzKJcLBSmqEpBBDSrKqgfGpLTtmQN2HQ8xQrTp1GULKZpIOuXiNE6KjB8kvhKotVhIFbAz
VCF4kJZsbTkdecWS8rrljH5n12sT39IQg2UFPr5luqNrozht9HIhHVrKuNXsqykGuSY3KmKu5T8r
coRH7COKNxPtctBMIQ7wylYtp6uDMkSQ6fzgBATLe0/h3WNbFK6iC+x+PsSrmq5/bO5mXmL0H4e9
9vV22P5AFNJfbtJrYbS+i/RbD+/3ZGiQha+EyoWqlnP+0RswwOgbifls92apOxMscR59uZrn4eIW
UbljYPwQaXRj/tLh4+i3QSf8oL+3ylwjbJZXbF4Ydj3czm1nuYosXhwkfRND98Hw9ABkwWOzxjB3
KXQxOukvkq/nev1WVUD9WbN9CHO/K/F1iby0ys3mgH3pNTVGXJyJB5TIdvByMT2hlQz/5KJ/cn1X
YyzMZ5DRDy84cLOVQLKqWhV2naoDKhelvb6jtYIEql/nwAA6UvVF4VvT4pjahOjer86Y8QQGUZhg
Hl91GI4f8yNlya3tq1ahNWUt97SvfwIFxS7IM8xY7Gsrr7dO67ROpO7xYsWioyQdnleBWCuMDiuo
A2814pTp4PmsLxZ6lqx32Wq6ID+iQvLCfj0IwxEqjzWEyETGkDok/KVXvaS5HcN6KdIy3pbDC0aa
+tR80nJy02DnSoYd9ShUmuBQ9PZOIrJUeyxRKOZmEVbNCDYNFwDxUc1r9UiDhuwHOu+5lx1azY9k
1P83Bser7qRuovrHx7zYTuUyvjdgi9h6Usuecj/DjL1xskCkNhhPhvz10+42SzlRhFwGgPExL5Zh
aRC2dx6y6F9zjaToG5A11RCP32+hz4lyE8JuhdzNUXNY26+wjU5iCDvcOJm6m1Qkl4sgRveGGBiw
VOR3LQB+gcG4o5SnaFs9IdX58uKofYHXuT/NTu8ZORwjSA8Jd4uCx/qyei+Sgpkg+UMAKXgp5qEp
JS7icnEN5Pndk815Mw/YsHqS9vsIb+m7JLd5ehVOUtl7OhNwDu8OvwrZk0NjxRVHfgcJUJvWvbmA
mb3uvG7BJXlMs6t3qHQSHzxYCQ/bCW+XvLORWEUG6oHfJtsLp9HCuvlPswaXDwZhUlW40kyYQHO6
esW30Maidriw7SS9jb4Vst9hNFwDs3mvpwkqkAPMsYZmFl+adYqXoF0XLuHk44deuMkBt7k1lamd
mGLfbwRWhv7xHhHQvEB9aLp6g5Tqe5E7bZ4rwzW2MJdC9qdovYMFXZCVDaYpAIRjLNEKi84VAbfm
OxAXM0uUdyo7VUdO7nHBL0dX6+eH2GFrlOL5VWJ/y4nTVm+ceBGDACiiPe9TAQjQ9+bgExBLKeRj
Ovie7sFnqkpa3tGKxBrlZ0EPdvEJW3lx/r9QLfKGWt733y4qSNhZrBQz+zQbFduWV9ei3lLxFZYq
vswdDmI/GViQ4Sg2U/0olmLxgD5B9vfNIcv7TkzM6QGIghydTbn8su8x+ZoKeUZvvjeGqJLjOBgR
9KvC77mzgmHkru8x59DsYuxy7eusL56oKmjHe2YsikWEJOlgdxVDmh5bTOHa+BDqz+cNutpMovOQ
Zkms6P+OoVAH6F161qSRmR7VkgeafzdPFWxsZ8fCAlFMtxCysOiBhw5TrDEd7GaScNzNdp1i0dV0
HvOC9yzG83KE8QuFcjFn4/XCSRQZXsiujqQxo/Vg7yRw9OXW7clGmHfdBUR3Oi7ZbJ+ah1Isq93h
FkM7IwuIgl2Txel0lwQRfqELrpty2vDK1dPirVOfi4Zlmgwn+1Dc/4Z4BnCqlgJg0R72xMiTpLMH
XNzp2BFHFD42gEpWe7dTI4mlWfUqTSoXc70JyD9fvcn7mCh7NxPz8nfPHbFUOFrhe94lSWMCaO6E
b0zgvwfTmRWFXlPRYurI1l80D3C9qRno/ZujsQFVW56tsxmg5d+gg3mrlrUN3kpO6202Lct8XBNw
8OxpGr5ai7M27Vwl1TmdukftTh4hfSzzpi0OCdao1DQ0i3pjgNcq4LsruQ6ROCg2UNpldh4adutv
QFQ39SQ4APohye+i3+YmbV9C3xQIJdOH+38kCkbaEKZAZQ53tBOp0KQb1/wlgzqhMeGnShVFPbwF
FhLtaI6qSaQgfu0d7VrqkUWu2d0uLtTdE4x56fQv5q9eGARAUSSWSPuGzHbd5L7jY8rZ2v6nyGIk
+p95OOj+Gj5V+Ar3EfrdG/WjiKG3E6SmJunh39/EPBHQMGwgE81L6RraDAVu7XnP6SgwrNZBf1Uw
uNRcNJl3FpH0S97M2FYc6BeSH5n38U8xc4shlPsccy+S6FQKwH9fSlpwwT5g/guObEOK6/XxHBur
2HMx7rPXMf23pQqmT3gztauTETtBUR+bu/snCOy1v8W/1CLMmFwwdsPhG97uvpqn/ATNkQXMTDvS
1+31roZKpi6Do5cJoHofsRD2rbkSAkdF4gbh9KGbI9keKomyzkqFVv7DJ69oRmN4rZgTaOFDqcjw
VvYUpqLpQEl7zqAX2ipNGDFBnb+Ffxc0mOKQmZ8VJyM8F+HtkAYUGBmm3CrFQ2scDpW+mNdKnjJm
kHZ2Nxea0uqAC2t+EYXG1h9IfmOkmi73SibYzEOlGpg9Xjc7Wt9VgGrQU4jwwpBNv/bN1izVmCyQ
KAld4XE6sRAoNAqerEXpKL2SfU0Row7+t96UAIoItXA7vd9ZAuvfZEEJlTKST45Bh4ikJYw1p/To
oNMxQUmQX3ZtiLyEMuuq/Kp0jrh9UiTbF4i5Lvx8+mAadqnlOMJ1iGKYQvhxD/y0cu1eIFfVDKnU
J99jKKq6928kSvYUCTwjzeZ6jDkgFxDBiMilXigk/r5MbbU0dTamVBymyEmaS2YqkA97i2bn5v5r
5OzSzJFabbGeg165HaLiMEQupYEw1jwuPPAKRF3JwYM6/vCTrjKTCOOUkyj1+Ce/Pcab+NH8Gq9l
h0bVirG1TTq00IXjJs1fOSw8WmnbCjQA3woZy5QbvnEW6rRhcfIUYgeTtqCwDAPc46z6FZ9dmNOE
FDGIzM8Is95BZVm41cG3JgkCMWESjfxmzQrHFO7yp5U9r8Jw+KSvHWiboUzGCSAtKQB7ewpPamGB
ztN3veej7xu1AulWQ/XBFKFHj3uoxS+/RQbFKR6he1pLuTV2aZGobizvOJV/z1Xk2nyp9ReuV49W
nw3cCKp3c6Lr4yvwJxd4BVsY8kvoVAqRy4VXnavg6NHSp1YrTsQNjfW6RZpQPN3EmULdWUzBfEbx
5+F4/vpqw8K7puPvtsojdEnuiK6dskbC/IBg5YFU8RVbwVYNFIojFBSg2kR8xZujIyQ5LPpWsMaC
4Bc+RECWy7WohYiF3zNC+AuGN7hSkrjrk3jqaUdfQEAe/JTK8C4RPLTf83PhjE/Mj+obqIAQzM2d
dkl0WbSo2r32ufCjCFL4fZdl8VgBnS3eJF8pEozCibZX+zr/4cDngSGEYrMSotI00tq75lrAmZQh
f1vuhc86Mb1ReCb3FFJdf+G77Olmn2r1vb3XFuY1BOfrS2gBFd7HONvd/oMyC2416zKQTwBDOI9U
wWa//xX77gqLLNJZsZy4LqlH7Pgk0StRT2r2sxHoN30RZoX8OofSOg0pRlj1tQ0fLP6flz2kZG+J
5JPCI30VmBmA5Tg8gI0hrusQ6BOvxWBNKWJr/ZZbTvgrMkir6bB46x5X/NnV3wYS0wWVY6XNjPWp
s37q2JgXusEmsiMBBZwQYygfZ0Dvmu/KFA6nC47d9H8fUJUJcr0/gbVx1azNaLYs/11L8K79Bg3v
kEgmA37GIWwCgdq4ibrNxIVKSJ9F6tb9Os7HyqHWRFg7NsOmua9P+38RLaGUIGSqiKIRZkBIp/yD
T5tkEFjptfa0bE/eWu3aEFil3XQmA0xUygtgMhaL8A1nwVz6HameTSE847ikMB0Ec0qrx6Wu7laN
RImuZJFIEglA8dP3uKEM/RuBmtXbY/jwa6LGIV0NTguHrpo6N4pz18yMOengLSsYB/LGepXWUvAw
FW2tRMG3dOcINn6aIo2IOjwVk75p8VdUw0czZvmg7pWwRunZjZbjZIPMzCONS6ggt/HQ1bG3e6NY
q61CydmmmX9dIhiipe25pLBya5S29ccA/Pupyw9zlX/rNJWUdfEo9RNJxXXDUyWPzhWSKWLGGMZl
8XZn5t35aL4eIniNDnP8TdHN/dlgVWrDOBpeIW5hDfNAdiGBjvMmOBy9Cntx5eciW4WxXFl7hqcY
0MuL1Z9OERytRA+fc4CwERZkLP6kDlFpqVkA8RZsdQH6did7tFxnPRq6GHzSEfhaZJbivBiTwq86
k9zZSHCbYfq/scxigx1eRqcpKMi0Dj3dbgLYZS3PylJw56a7Gz7aKIZsGJRx8pxVLjzgObVNoLTF
GRkIM3cV3nD34ZDXtuej/rFgWGz0xpGvl+zzcGaaM+KLyt8H4Z5ta2i+4q1C5zA4r4BpQOE8OxXZ
kuA3/kH62WGHbnWiv7YqLYyso2jI6Cc+kklPwDFYqfpQp2wbXoGLzAufW/5H3wHs983bpPL8Yhny
1sS3RFYCj8Tabl9+J2OGVX8B20AFOiIoboRyJfYxAbWAbmSjoyAeY4+kKQ1Uy4xosLvFMsV0ze+V
LQ2FJET/U8oipK+rXSNVEB3QxVJT+TKVjmOHRUmkGqcIh1itfwadvP7CtnRpC15VB5kZSrWuMOQE
/aqCwsrA6KQHaFaJLt68TAOSSxWRZp/BIgGRpjPqF0gbG2FCrirjfHXKKH/yvx814H/vlnuKZR2Z
OC/eM/xd85kyLdCEkmnIKDR58PrBmNH8cohpHDqtTlOXx4rtVfeOzbEwFEcmWMoL0UVV5t0doT+v
qkft9T9PMwypzN7u9W2Lt9iX9mu3He4szvhg1k6+eaSb2KPp7HqoCqXXeMWx9dmNi8IFN1TXB3rm
T5fbSc2Ft7XQlMp/t6wL5D57w3qRKwjYUZEWU4gMEa+V97uV00j8iYBImGosHr520eGhByX48j6+
zW4eeUqqCe9taEanti4F7LyEch/9DWna34yKHNNXCh5U3E/QgqC3JqVrIFLhwCSL7rHls+VZtg8x
1ICZxxaRV49wi539oIYc2UfuBOvoGwiDtp3cLeJiKERJ46EPKcqRT3m9pgoMlnMiqUesi0V5D6MQ
AIeYr5sEpEBxSrlG/h/dDYbTY60YmztL1rEfHnpu8fi8Xil7eW2i6Gt50u32vHI9p/M4sm3oRr1c
ydO0htBaY7bLi+SJIRLN5g2O6IkSUEcbDzGpYB+LEp6Jzt5mQsI3jhJPDbMtFJAnakOPPnO8ATnx
fh0fmztG3yy93POq1vQkHzTG5pz4qWbddTNrpNS5hR5WTUnN48xVH+1bwGvJ6tbR9nr35k47D/I8
1OwWkLm/wboMeD29+Na89OnBMYfO3UEziun8Azsya0YzsO77kmuS5sxgr/oIIaVYE0Mgu7LB8ONz
V++w61uPkmzK2U1X9jJsHcl24iFXyvsplzcgGfCESw8PVqtDfpX+nyIKDdsLV7ZSft5qmpmgulVD
HyzEzzl+wLsrnSMq6hnQzc+oJxh6xqNgtRMV0mUJ/DHMmCB4BWHlHjNzUOP8tEmirQDdguyxbTVv
uvMB1h8dVmx/rd9omupiKBjqyC4JfoJFR8r6Ma3rpNlBz5iHd9uhS9dDc5U36lpyd7fS0EnSVZkp
t86k3d3aYZwewh0di3BPjvuZtUz2/pswa3pZY/OcSkTYC8WBjsub8P9uqdY3spkVc0SInX3XZ0RY
oZ82L1ZN2IuX4Fk/dqQTIp4jT7h74GZHPVTIL9CO6zjaDihf0g7t9oltYFgouqpfIuCi8JUZpUgw
dLSNg2mZ7LbuyiYTtAK6KP1edDrKvXKFAdXzfblHWWAKc0RNhXvDn1mC1dQRwd4qxO8GJQgczV8G
xeg5ukkT7L89+ReyfHnTITwoo3o96QHEOk8aXE2kWQ9PlOUvxSG+GaOuVImmaXUjj2iO3pBrQAwh
sFQ+peyDY9O/46P7S9/CygNQhAj6/am4HZjSEB/QEoPQQrNuX74KNQvkCdgfpHnqbQt/1og2jak8
mcdWnyD9xAJfncY6aP8T+o5ZXOxlzZUtwqqbz2lc5JivI4pWZmnKYoTwrzPALIENxAjDf1Mz8JGH
EYH4uaVk1MPPrLJdvDIfiKDKYs9lagJb2gRBTKsr6NcrfdADJoey4EkhOtx94n2q4FxYx32mRxbd
ea8tBt7+jRXhVaj1cHu2nOFNEgn9TqfbM9AfhxSJczymTrCnzMqCGpLccSD5jR5yoAKVKTPT2WC6
gKz2rsKmeaSwDXiDNkyN051+qyeEeZ+GcEnQmqUqcjgMI2U+gT02p6z2YvV1qTdHAfvv+Rn2TJOE
hXfmbUOCvgqF4cGVpxNhLmjYDWScx44W0IHAWmmNljdCyptIj8B9B6z/ZbGH3TOZmioDKYDpTb1r
gnNTqQF87Y1WwwTfwkhrn/DdCnKFMQ6o7BzzTgeTfUzvVjNWzJnPL/WCxcefMOuHrOv+EMryWv4x
QMDU7FsiBBR4vqHjk08RAEkwIivtK06Jttw3rtkkr+gJSAr5+prNbLp5crRVhPQjhXKDnpkvD2lV
X+D34i/8yYPLOqxEXFCoCLtik+12vQe6a2b4xj9b5q1XzOmPPGoKnQYZHNO6uudf6DkFvPWHSBkj
KlSoudbImNOsBJ3CytyZC3yN+hSiijTD/sW2GlpMcKuTxupZJbZVis/aVA8qQIdRYotf7X8RS4n9
VhdOFdtGKU0MPg3GywKrgYSQjz+eC4Cb63Csqj0B+GFVQQSZUYDyc1i5WVhDXL49nnnCD9/7NJTr
eXuajFiDz/zEBnjEAXnbX3Il9/OH73r+ACbZF9DuCoDLepfrrLQlmE+A4dCs0e6igCSWIBUVxQxo
fg5X36UNmJOFVRsoc6dpqHDncfhG5rDxC59EWRU1Tcxh3vvFJqoFt8iTVFwm3pxkVNFYytNOYOM9
r6KtjaI7/xds129c8yRNSAthonj5bxPt2hjeHLzIfg/UjQxWYUGmALI6xoHPeHeC3hLttV4BI3TH
XqimL5IrboWaZQwqf4rLogegHpk7Zhj5VZv+FwAtItD1GmQtd/CCU8/c5cIgHtVeePdkEXcIlwOt
RgxqZbcsqnPhURAGUElb8bZBjm8cNnPEufgUCSf95krXwczNdHXAZzOK+EuDFEcF5vVPypcLkOEe
OLoqcK8Awqs7+oim2tW4oK0O+E82qDs8QkirhO+5pFDuToWOeUoMy63QVy+B0P4b5KZFx2H74HNk
iOeLuIpiAe4C0G1OhpHU5X9WYaHRk4Sth4Jys2Ut5sKAEmzB3BZqinXpqqr2pk+ReCcblaYqQD1X
XpWp6P4+GbUdFpM4SCA0awcS78roiitxluhvph+vjW8tHuBN6LWTAhQnGXpCKHNdN1VUsgbwHj0T
F3E3WOwQnFXLaxJY/T4qICq5i/KDPARNTAcefvvv76LSVeJD91Jhes1VF/8uhqEce0IiNhsOdz+l
l71xDwTfFDl3m/YQC0/TFJDcjRQglEvvLX82nvHJVjEg7ihE3XqbPHrEMHWLDwSmdAXhqaasRlHs
wIVW1aV3BKybJW7s73eUVYd0uLSN0C6ZcsF1qLj5yIAWyGm5u/r9ckE8unIKjryjVqSX+/KWno5r
zLccAZnk8yfkFg/JNNZIG6Z5gSpSYt6LlwZdD2UBNdy1TiKPCpB6IMArdEGAIEfXHnqe7/o77nKL
BzvEJNR9RoM5ebQGZVA1tFKNFbb+qvDS88R/q8mi1wpTE6KGI+8sJgb9Wnd9UhTNu/VekT1YcEr0
i5qNxj0QteT5u0nUZV5rlCWNXs1Fk++svdT6mCLcLckUGr0hb449EX5JucS7/4c1fGcEvi81MPtF
BT7ZJCkZavLq+xI8KrJz1cr1BpcEoecVU32JW4c2tLRE8Q3/wJyaTt+dp/V+cNq0I0f0HlndOmM5
33vUXvkg9NuAYuIAwegAbiuMAJeQ01NVugHpgC4z/po17Om1Ra3qPTzJ1eMcKO+dpNZU44Sfz+py
++J3Rl8/p/QNK82axalS33dkywi7Kcf7eOLw1nYeW+Z7aJffgxYOf0GxUmhRSH+plMj7+NrS/Xbs
5xZ0jcrP773fAA/pmkR5GjbUYNsdiqOqS0kWsB26nxZIfzoXwfPlfn+f5AGUkvP3qq5EuWwNDwUL
0RmTv3veJkfrVy0w/EwWW2g4PCLauqwovQ8Hl9QFhGYXjEhA1UfzdeocVTlCUzWIP6Bz4dOFGF3c
go/VCFznoqu7+CIS4DL1W0CKy/u0sRG0xS+UtUlCTPeCaO/dP8NeiR9al7ZvnbnUlaLbhU3a3qGm
pkUSWcHXg8IIEGtKmXqfPKWR2oobJarFc08CNfVLosGgRSormJ6J50iGh/A8NksPmgbcN1cPb4hl
QOSYsuVfQRpoXEqM1Bdmc8tBdL3C7lCD1UZrnkI/Av/SMxDFc7PJV6mDZ7iLNvs6xEYvnFgLdww6
Ao7kewYARMSZNQ1XijBbXfyN3ejcAHjt+BVuTnD31qQWlV1WTDWRwVc6n9L8qACHM2RUX3Xd3Sqb
gM1MiG+2ZmVFC9hS78zlF84WNImO1kVBFux7wo46PzPmYWlz5uUIaEnGtxCjXuh6XoOWxWzUUHvK
9Si/NjjdsuRaoicqIX7voGwr75hbG7h7Q9Ll8vdzhhh7ZpIhYIeup5ImSzTDK7GH/zJFWksiLeeg
e2EYWp185xui1iRA8yU5NmBbeUK+V0RfhP/AoGsr2LK6Ac4J/kXnpnknwWwZGdIDCcrK2WVdrFxM
46iRMcuHFxf44TbDpjOL4I1bykXlopMBQ7pRi7EOYfu22HI9+E9gmjQefrCn0w1S8c3aPKH7AJPh
o36bRKDkXwYnpUWLiGIC7POmyArky6qyorLPmgteiAT4EcEicmDtEA2j8tsKzuu/UbYkkIdvmH+L
L3oqYDl7e/2yA3uUVHEngImxYQg00XtqjPO5kqHYY0JlaJfHz1dWZ9odtLzAlZPWyCq7I5GMxOS5
1le38lfiiu6He7C5p9H8iOm15GqH0ZTHXXBLc+l6sw8nLLgBr2jVA9Nad8wV4xjoUKaeX5+H8SBe
PiMwTbmI7m2xTd0q8tVk0G5I5kpmKdhBQ5FMotHjyXhx5ii4DIk0LuMwPSE14F79Hl9zj5P5V0TC
wdD2FnjBvJFi6R5c4Wtvuib7y9+yZZoSf8KVMEd3dSPP7ri9gTtEUcbUTAiTXQLF0NnqJMstyvRW
dcPoK1R5wPKfgFPRlBEew1b24sHClTa3ZZ3xJopFnW1YDd3XVAsMVAhvOKWYZh/m17QNZuCg6t/1
t66zbe+tRXz7LKsxu+LRfR5WuOyEPwHV92/2jbL5vx8nXLbjRti068OefZhiYItp81OiS/RaeTf3
VYzoYbqAY6j5rD/AGTALDdET8WtrxrgEYCSBOavAfBkAoEoTMzTlrk5i1d+VFqXSmqD9NFNuFDK1
vvg3Vrk+TZ6RBkmsgH4gwUBFfzWRSGhxQaKL3tzES+v2mvMkDBFaodZy89gigBZ8MtArHtdcaAtt
DKlpr1ni62WjsMulSd0SGXQvwY/r5Tx4Abv+FXKwu8b4/a94wRWdVb0r4EA6y5MESsgmxZTojohU
IVYaHkiIva6/8aU18C6rZlIbo0v6YYLl0jWEpTpfn9aCE99HTuyty/qm4Jjxd+COgsV0pKjNd7oZ
YeWixhzPLya+RABa7JGIQnFXcUsNOBwsd5Mqaver1rDvGOr8zesTuDUa8ek7fi/QyoXZiwuwjuLt
mmYmB+1J8PYla3W6sa3thOjan8HW47MsJ8e+WZqy8N+kbFFfNAk3oD8StYlUiQ021kNefbjy0cU6
Js15ceFq0x0iu5SpN5onuSGb7zxfAaWpr6fAx8YWQRJiVJHoR72jATPcK4c6cfP6Ho6i6Kpk2dWF
WyVszRjGJ5xwqhuDIOSGaKyhJxDCyGv1PG+/2ObZEfjcTBUmv3AOL/6WS45Wc2xXefA6hqR/TiEY
eZ1V2LV3b2dQMBJe8fd1fZLf6cDm4A5aSvmVl7W1kJdxATAGQnmSzgFTmc6dOeIDB6Lwdz6pkYML
YYboDAYx5TiwMbwcmP+j/rEzNfcTJNO7//kEyEEdZnne6qE6uG/QhDSoOGqpkmx1WO+6rofqGKkr
7g3wVyT0akdmOJ9yqhw9tSoQ777y8uo1htcv7zpf589KKAoPVBAYa80re2+P6Vs4U/G+felcf4z8
pXQznEkxA1seUeAr/OMDlz1DPUzSgJMCduu0bgNM1MMxM6zPnanfl+zVhdhyh2isGZZklJBPYvQh
egKvoNjl3bUpeY2i/9aBnKP+9yQMgDUs2r8G9tkz8BO85XIRS8YW98k3f0Kxwkq+q0PnHoelCOI0
hu4lYKywwKFMrjqfUXG9sF6cW2gAuS0OChWIpuJPoMJo7wpwDKWUFpSdzc8m1nkEHkQ94uAwNNiT
m3UqYbxi+zgxx+tNvS+gbGKqnrf6y7Pkb65YbEbEhONM2ik8HCl21nA7t04QM/A0wPPoLLWw3sKG
vjjMiV7JHDVu5mtkJvYdYO9YCWoCno3KLOCLgqi2fBrxKMj2nmIbVRzsCI9U4yGSajrlpsOZEaxR
4cSYBn/ZrNezHCnvPiAio6u3qGrTP/gIpeLUkXkGNJ8MyXamQaEg4x7/pnRoc8JJy12jHIOu//HI
1Sp3P7xXkvQjuQlUa3wP/6TtOlkT51Vn2Cj2HewxJi1nTMBnJ4ghlViqLG3hPIz+GsDCXHd3Ishc
ZbWPP7jxuaynBK8TvSTyJeu3SwPCfG738DP7LXC/ncj7udI9qAm8NNDmA8+ktOtfhzRGX6YRuzVF
xqidKKn9DT1Elb9z6gHJOMnQahL0CS52utCpeNmY2bHAPdlxpEQIZEhDoOoNKmWivj3yVLm3b5RA
Rz3k5yfxmeo5X1ydvI2I+YYjvoZc6JstsiU8psEDYGar3a/r9QrQIpg8s/EzMaXHjVUavJNFmhH2
cntb0gT0olrnctjJDd3iGnWYMN9dTU0nr2YnG8Z7wCrBakbmofwAuSdgNy3DhGhaISk3TGBtSW7g
AdIz5i2xwjvXV/355nHSpxoXwdsBOqSkQjw4BXlQbJ1MHXViiP907JK/tTR6JX31LSwOzYBAy7uj
LObAwRK4IeyiTzWz/2aDHx/fZ83hJSbpr8x9QfpJMHPqKvJTeBsaCuof8kzJz9A5akUeY75DuEqP
qUINIH7zCqiP8/ETcAcDr6c9z0e3RF2TRPlMBq62KU5rcg0ro2mm4KIqfuoVRkwcUoDqTcsLar1Q
5WGOh3axQXGyUOQNBIQoCPp9V7JPwc+VMbJdKuNx5o6g6W7NwZTi3pZYmygo7SjungritwVT+b/I
5F3d/S3yY412QSrR/6fuk0qMt3d22/yXWlZqL9m9ZgO9hbiE0ugADgUdEA1N4t/Xu+FV1gtSZCee
y5DAUUOkJ/iSBpDehcc6uqM/2/2A5NzK1eI8kyWQEasYvIy6ZEWZ9m9LW++nhJkzj6MbzYIlady8
rvaweA3M+DTEH34Bqi7sr8lCcbaNcB3u2SOSuMsXs6e+pG2WnhPW68TAknCr0KSiuMTR+BdCNScU
GxoHxYlvH35LLdAnz7RLE6CYHQ98vZFVqcMzK1U6Jyq6zqTwrN1o/00xd7/u0u1xXZc2zz4DD3ja
axUIhTCQSxviRdLS6XlCQaULT2NhO9hrWBhXrbR1LDRB+qm772trnbowXuVUhq4+USrPg/3PRENT
7u3HPesf3TqJLoo2w1Tl+vLH2D/fMphg5BftXD+Q1t48NHZ2n5zCao+8pKjwfcz+9pniS3gNpbC7
VQacCqz0OJjpSmPct4a640iXZpptuPCxF5qM2CgJsbqXqraWDo1oPZsPO2MccEBJNfcTVEOmugS4
4vNmuc8OApHbZgbykWIMUquiS98Eg9WZGJ1rZ7yUKRHP3g4BkKL+D13cIJOe0JeohtNcw4oqYs5b
REKAEN6lNoINIR5c9Xg2ifbUA6o22xPi2MJIqmzw8YNIPq/GEM+FU1DrAPO8Y4EOzrhrA/ZXdLVk
VQ/JlhzjbK1SNEwW2LNSTfH5ydfq0I5nU1DVOSx6omC19cWigAvpiyjeQ+2oSrRDm4EdrPV9cHqT
o0gyrWLkGXJjovdFpbMSQy52a39FK4yg3fHoKWaEOVaCVw1eE8+DQGP97B0zSl811LDe07nBy76q
edrSZ4ufvxH8268mD11f6RK5AqGPCQ7jSu4iUYLJ+7Kg9v42MV8VE8TDcVhKxIbKAiRWhe+cNAyL
TufMHcIZvOr272Y12ow28H/bFFVb5kKRLU8rY59lDaE83EVcbsU+qp3KzicO3sMwPwhDBDwmg7a+
zGNt6j0DoBImye9Pq7b0uamoMdqKOqWlPtcbQ9cTxLjI/4yZhYvwBmP2rIQJMdVWjlGmdzLTHrk6
gsGXLARftUd6tNTk5ur1vg/UH1yuqy/rHQjtUAZ3RAdmxnS0MyLS58YUXNVKjTjf4A6HByGSoOag
kZNoFwWmfxtLIh0PkY+oHX2ug+V1SJK8AbwQxsvp1CH5ESw7+kUoubsetDcpp+TXF5MCpZLbNUK3
Lms87+akxV26X9c13V8RLNwdjQs5d52PoFlJWFnUbAabWDB7cMtYmTU5EBLOrL+9th9L6JeMkghf
FAJnLTwZQt5EYKJ8qNyG3bWymuzm3xhGNt9S8caFQrFxhgRy1i7cXfqLyk1s92v14eSAXUfi8t5f
p5MzxkNsGwCy57AD7wEFBVEnz4FLpToUM+WDw0TIqMuOBRlJnafuOy3GNRsi5UNiLhfwUJlqMown
Ibt5KSW4NltGk+JhboYrOV0atypWoO1eH5SYAWx+hFgkUl/5ToBEjglu8r+iv3YB8d25msrmbAt0
0tJ7glkC9AZdAzhcGZFOhkyLAydThIIUhEZsGZlG9heFDC/52kZ0aQpWrb5/RxrErkadI+zM0eo9
2qEf2j2+1C4dv1tAzNOQDcslh1tGdEWSXNiXP73AmSG112u4rCPwWANNkIyjD4asHgtFEES2oMt1
AzwkXcQh4irxOcwOOUUIs9IjJ5CvhOSfwDUDUMMok8mjkQ8+MRteCMX6TpitwMccUkY9x+wUaaNy
OqyTzRbrM6XukxMph6ByS35OcLnD4L9z0BaCaMkO9FW9FMMzUKQ6q2bhXMiGBeUL+aF4e/kKYSrZ
Kgyu821jFO6K6+mSfs5cSJAAcBRuzOTewseWNKrdNynZDPm71YL/BU1ejETLvOT9AF4CPzW8v283
xTii3oC4iRje9Oc8FXRbJQQrLLUHfw6OaEHRulq6RdH1c8lnN7F7bdl0HISxuxWYQYeft/D6M3FJ
GQZiemASlMM1Wv4hbQAO0ZB+uVLePJK+zG2YsgB1EdFddc82qpQBt3PAb6KgNDB4CXKmV+uy2M6g
TMdBgFsBbi69v33xVLgjmR/TalNgCZPhGvRcVRY+ubwWRNwNqZSvGWKN9aLUxpquTBwo9fOv919B
eAd879y9DaZlAugJu7oyd0gIN5i4XG+rJaeY+i2of2PqW1EbHwFJzkYHDiLr2gy7iaw2NhzLCWwr
YznCrKPwFx92LgYZpB/9Mir28crIjMAqa1UbqmGuKI6Uwc+r94OfVIX0AV7gV4WqX4+Tj/Imu9Ut
EK9YfTAO9WwPVJH/aOJk4hDDTGh3kfYXF3910T7sNxYuwr5vqjbjdV9y+PTrTnj2g+iPDRxenLIn
ICrWiGS0mEKO3h350Al2i/9HPDGuA5fvpQe/0oXMMGMoTKw+eYSWMTVfuj2DVAfTS8MpaYhcVyoI
L2FB13Tdv9JdSSO4YlhQF+31ps4clbJLZye/W89dORD2KtDMWJvprRg+smwMPTjXNsqWLcL8OZBz
/1ydFS1gkFb5gPfzfJ85uCkTY4WB9YzpJXurh3H/rvoFmXLkAbmvZtuQGy5sKccnIA9j76f8T9hP
OB9Zln5JD1555Ie1o/ifDed6hnPCC7EIHS+b0RrqwXu4VEOup5+WxlloOxxcTxuS/CBvCjY90asY
P/vjUIu37fKjqYtS2EAH4MQEnnQKLVA4sok+VgdU9CsP9qzmLQJVBckGUeaFod+NBJflDbkq1r0H
TuTsEnAHwylu1AAEmJ/kYW9eJntPfEXcQk48TZVDKWeeqTFeDHNAg4wssvMYf6Zg3Zf+hj8TVnJ9
X3VSX9G7kxNln26NmZR0chRZYvbWKTcwkTCBkmTc6ruHsQufaewCLvTyYoLQJBPAJUgQwFyT9fD9
10kLKCFYnyCeZdIHjijEPt7Z644Q+ns1pmBKiZ+C5Ywe7DNb1G2eyaIQii3xOD5BGXaivGAaQJfA
ps4GogJAzaJrnO4PDXEZ0qlVMHpXbWSp7x1KjQv7SJZi6QTMrSTm1mAPadM7u1jPouVEx0dOGhL2
TTqCa2Y/k372wxyJ0q9zAxaN63U+tndUl6egAd6keZ78Ew0h1R7IUkF0JOx8Jfd60nl2BOb2XR3m
j9Bc/iLLH8w1f7ei28W07TVdstKiG+2z5cGS875XDN29zKP0L/AoYYehFFu/e+2Q+RW6dI1CBnx2
96cji+vxyk1kINAyx4TSG0df+F2UtoYJFEHF3BLWCAtjGir1oRtLjINzIQ3JG9INHuuLYWJI5G0R
3ywn+agxVkwCWqY+qMNGISQfFc0LuesvsGA8fbxFfNzO4iviVEZkPox1LGsrsXn22BP6PYeXF62u
umAtJtZvGpdOmCgh/Vf9gwDVCGD2iXdONobtS0w+jOzGdi18x/U3OaP2NQrdbhA0S9EuBlWok0Rn
rQt7sqCHlDJPLMAUwjxdIMmOa9aXcK4bIxgqsGE81ebf+P3Oo9q4RrhrMWZ68d3Iwj3DThqBmtZF
0thBpqQp1Y/nOjsIaqiTiMMlA0z53C7xOdeisSNYIrLAhL++3R9FySpj9YPSyNLf/9d0Iao0SJiv
Tzu/V2Q1L0wjMn3zyk8UqZrAIIR0LIbJ4m5pAHRNAyVv6ICr4MlF+tn5Kqri//nvudpK3N0TPQlf
+6EfyxiUyR5AP/JHYKh9xF7m1AlLLPCuR2wPkRcbyM/xIWfCN4w2SGyT6OuQMpPJn8HcOSDXkSf1
3RYAX0IJfykV03SHNb2xzaUBvUrrKbWM5VmzU19TJI/AqLLJtJWWoNE/H8u5NC2wjagOTQn65L5H
a4e66uNV6vgU8MAJGCVtUYcawQMjIo0NfafLg+DZhORt4M34AkhD10KR9i1YRoI2KM+tqfMMtSBg
YDzRDU8xGymm6cVvINEGsl/4tun2vAZELbX1CpqKZigfYkekk6EW0y3mazkC+48q3kyVD3a5UpYd
aUAJlLqRXLsaDRYUpxZsN3stULSY0+3mI1H3xlReOk5/+1E4wt3NOFu1GaVhvPil2g4pJuXwANPw
FG1Mpb5cUFQhpCk5uFHfc9k/xf53wDw+OEsfQPtJpRqvGqJocJyQvVfE7gf2J8FC782V98m0mODH
vH/UIOtIG9+IXIxIY1F+FNy5sU8+xHR/3+GJG1iZoN7xp8upXrt7duNTuchu6JnDJ5IM/GUejvVn
8JN2Xv7UUAQJpmSh22N7ttPIqdL18wIZ1Lpeb8LoOSXi9DXT9x9Qkq6pQSmvQtbU3GYmDfiwBrXb
QgpO9YARKkDbm4b2heLxXo9WQz1ZtViayznnHK7sh99cdjg+Atv2tZ4mCbmp34S86iJQlFtjE4x6
mXf7yTDVcXkWJrddpvuxGAOg3gDi3gbh/D3S9aVSrBxP2jiaw/dSJR1aMw64p4vozbElDhu55r4N
vgW3fJRyK6Ft/f1Tw+onsnTcJwHrt3rAaPWMA9dXepK35GUf/0t4vgLoRFF+Ka5hb44iStVi6T2/
S/eIcpB23bku1hZc73krR7SBcVZsqpvaAJkGwWEpjMMqaf7Gs6ZB81miVKFQVT7B1e2Dtu09r7IT
gZ0xB/iTnDKQqr5LZkJx6Om98l99Oq0zgbbzLyiqmOR8BQ1xmWiv3qmYmebFRWx9wNKd+qZEpHHG
c2+2IidZ9Olk2TqjDfSzHhFkuNRU2fXhIrNsivkjcrPLQHSgUcX/7sQEfvgNXrM/pUoXiMOSW+XF
nyzW3Ub00Y0whfFVSHDR6gJo0pgnq7jPWXKnuGSWj5DEzLk8C+ezeLy5QVtdnu+zQjwZAUqjs9BJ
K91VsHitL0vuQ1SvTxxNGInFno7DmArXyivS6NRVdbIhwRQL54vM5Mt/Hk98MsLIHyZ6sID6k4uJ
e6Pp0QXkd5p0LZEuM5fJNnh8aab07+coouuHJe1xihvSqWQsuMnpOSsGr+tuSdaQrXt+No6IiBpr
Wpt9/65zYu+zY32Czgu/YiPZ3rKTVG2e715Zk7gxBb27y3x7K6C50vOkJKU9j/fiYD4wYLPHgBQ6
vh7c2UyoU5a9lMFy+csK5O6OAnQNkm3rdVXkf79XFEH9lSIlECiS17Limowr2iwFDQ0cebKa4fMJ
Q74dxADjC41+Qrdfl1MU6FTtsBROogtvHynXIbGHrWp5cvJGPUgrqHr4XsbjrGSqq9ZX65qzZ8X1
kMNVOjHBdk29E27F0jZg0485VqT24+7ETB/LSmRnxrMm02dASDY2GzRye0gcooCSw44eKpeZTkE/
2C4622Hlr39t4aTu1eEdC+RuM59H4sjeKrTH3RglhV/2XfJJwPYYHhnmtixQFm/8/gf1cSN5v//l
K4Rkz25HT3lzrMSFrRu3aSD6t72es4+3l3qP/sdhCUETeS+/lcg86ut39MP4sc4Hu/IUCIF+8w7E
3JNsZEmN+6hgs/fv03wMhjJ1ZeCrhXSrUu+KZvJL7WCwxRe9PTF8SNqu2SSlxM5JSi3EsEeQrVqj
GO3qne25x0b7OORijZk7/yf6rAsJ4QOJqizYbli8KfQorKfg4ZQNH1XuTPd9DLKKcr4aTo8kYyGF
IPwVEJefAjEcnJz8kh9jx1QGSbdcArue6C0AyGcquCpl19uEBw9aV0OrLooVgjdQEC8m+ZC6HsSJ
oGpfoq/uOMeig+vUnaSV/KylG7kizMqwFeKTl7FfhdKJHJZUZEf9009eLuvEA83b6pNSk5VPAO4O
02RVYeGn82RUrdI3sX/BY/V6t/aatz4drEfhUVv5kKpGQuzQYJau2/z5+YxJ40Ocpk2rSrTDQAn9
MthObfc549benopduxPoKdMwtOujtwpjO7V0u5lxNM48WyUFBIysu8NUQNKTNRdVctb9OsZSZpjM
+6NOhtGY0vTAImgTnadfyiV2Gkr0ukm5rtCuG8wx/phWCIKzMgsW1y+bJhL/4ij2KMJrdDG3Y8fX
bM3npFEjvULYhW1qf0qZWcSGtoxxfB35IqFFQUX60lHbX4mN3zJY2Oak54mHNmPalsOQ1n5S9rrs
AnGVEjl7VgpjnvVq0wLGnodfyTaTtbL8SfKXW5LO1HT9Pyh61zKrn87q1bAFXemDw8WjoMZ9+2f1
RmWUP4gHSrjzCBdNkTRvTpKfHde3d+N8uS8c1UFwruwB5SsinDFhwDtg4X3WSepcXEBcOLFrKca2
0QWL009RjqTYsO/F3Y+aktbVDB6TrlrUVxonImBbZ5Db4BQWV/OdQOEF+r0YyfW+q1xPi2GW089K
/nUd4bgniIi4VA1JUDJoH1dDpM7plIry4SMJxNaPZ73/HIuCGTd3KO8yAKDxkfVfxGOxtH4Snvr7
aQJXwlfuaAoK0ljLoSB+AscngdDxzWcPd2912vCp5NOj7PI2RhThPZE6bML1zA8skA9UNC7BPaGt
TNghPBc5IyxUfJp4RDsXD4w6ntI1bIcSYsFBFGnY2U1n3bccUSx40la26cJbpXXfjdJVBpqmyLmh
PrnwWmjlzHb1xRVejVsyvXpv6XASxq1YAlegivtZhfx1LbTgBlMBvdgVDc4pY5x9sDvFVIfypHA8
lwa48mK7booc+vYIFvndp7L9LJbXJ8X1JMdLzilJsmXGsbZlL8FdDyiLp2O8XuiKKnkp3ljp9w7q
JntWS6kNGtF9M+zqA3ERCoHHcN1ie5JXY9Sm6pXctumkF2skAkHZsXyErqRGMYu1U+eFFpSv0570
BQjXnkwUsN4OQVKejTuEnVFAX6HY8Gc+B0qel61pdnFK+NC+LjBciMy40T7HLVIwX7VWu4Ne6Jso
Ejh1jOAAvRQ1Amek4yFjQ9seMDr7kEJb8r1cH2Wt/Xeoar8ENIfvOzmz7NtHypeSB+8RwMJg/v6K
WQseVLjBNPEMmurDaxg2L1aUnc3u/ZEIDkLT/vqv2KqT+1M+5pbehmLAlbxBLHB0oLHqZxPPDwKV
yanRfKSeuIvgmxROBn7D6t2vVQx5Sgw8boj1W8hIjqkDvEELbCWwTktIlll9+/8gGZ0iR5EDUdhz
c75TJ1M/oj/e6L73LNZNztlR3y1FGDqLJ78+nGjMbPT3jXVNotkbW7iYc0R/LU8fVaOMPi0PLDBv
X3W4OW8gbEmHh8hDccPHIf0sV8LMhn+5RV4vWxKwDRwYX31cRWOiHJ0NWysToJu+LgQtgqLIYthH
RQWemGbtqx10Ky5UBNrvg03IBt8o0eHI6zByVgDLzS7LfoHOKroeGhsAh5q2hfxkCO0QPG7FZABC
ffrF2GAL8eElD7LzDZAdQTJiDUn5E8kB2p61SG6WU+M7McW+xovqCcqbME1VaoJq6iDiK9/brKME
16FKXxhZrQHW5YLo5eeGJzyIN14jeiQOEoU8wG14grfj/tnjZEksnJgk6PuWsKsgFzy5qcgUFcdT
Uf/X1IlYVYpMgaUSvLN1SXV1bg2DvADHbsz9MDrjCBWdpldfxiMhOEi6klR46zHtWUVH/qyCIxq+
MHqThSLXxjRV4uhNXeYn1IVAGDgtpBoXEYRzgTn+x76sZ9rnby7oU5rNx8Lvc9gXcYEznhzeeelk
ntC+klad4r9GyGM6Kz5+4nWwwV/9wqbX90IWE7CVOpP0d3+bvh9+md3ZcfOWYki6WB3Bix2mku0O
w5+8yxq3znT7XYb9wkOWjIRoF5b54rF2Zry8ACoHh5q9aXxI/CwyEzBrqJs4dKYk+Bb6IXeSNOdK
DY0NlitbrKJf6LisdtSVD51X0CGrRO9e2sq+6Q65FCqPqFvH3CNB8i9gaL65JjZmlvP1b03x8yZs
4eb0lIZSUnHHhBz+xpc8XI2ajh2hDR3Wc8KFuaoH9jv211NKralLX1vBdTI6eHwz7mgdGlQj8eXA
xfrlmlsw95IIRsdhn2r3GBP5SrCYm7LJeyy5481chjI9J8/+f5gYYY3xeGA29R+XvGRxIJTX3NMV
545zd+urOT2lOPCyOQ0at3Zkwzs0usc/pFkBs3ecg89ihK39t4Sx22JSlnU3aBTE46OtoW1FDITK
7lXoehwiKwhw+aemd79VN/gFd0yfByZLpcCPu7oURwVlTBLKtAhzEqrNrb6UQR1Cd5J/lsEJ684a
Mhdqwu5A3/f1BN76l4Eyb+7X7tsdUwOk3/SBtPvaMUTEZZx4Fje0nnTzN/UbEKX6vp74+zVEeSno
w52N20IXD/2bbsKbhmtbrufz6T5rkQ1OHjRTFS6b40Hb5gpZ935ZF24CNWMsf/5AJJDIhpVTqOR8
xyDqPUlq/sPCpyAc9zrJSd5D0cnelckn+isHSL35BhFv+HcoGGF8/oXZ/LScPcmW+PRUEFxNACy0
3oh4lSuzsgknykhtM8JdV1yuqcXkxnc4eSmYg1+hAuLLwptfIazgMV8qtJcAA1eRQg9AT8zj2pAl
HRSJM7xXkzOBbl83g5hyx8YIQcpVq0PVeOFO4yKcaHylZnU6x9/AzKnTycTV8fRgafOJD5gTZudS
h9rFCu3GcjVu79BkSoZ4kemQaMqynCg/Y+qBfBEYd52Gl287kbfMgqyKNm/vwSKQCIH/iyWtzepG
7SYGOAFeRzaZbeaMSjq3T4CLPs9ViZN+Gm/juzjzfv2kYS7rFl+S0OtuyvGgD2Tr8jwesffxze+v
UkaN8hVbMJLafd9vNtq9KBUKxsxjG1m9bTlGY1Pqi5Jl7XuyuO+3OzWxT6JGMlkaA8Pii962jim2
cDKEjX+Cp5VfmKlRxaDxvrEil86zfn7wGmnbYniuggCY2+VZTcSqPLPsV3r6yzo4Zj6nTa88Djwm
Oz1uP1TyJ1sCmfaYi5nGgFT+jb1uMZZWvUDH71/aw0kIF2zKJinpMe8iXI1FXGXb//IKwFg5fDcS
SDVdzD9YL36tMXv6xXa90IodsftoPeR5h5z6FnPY2UbIL5bT+PTB7i4Uik0SPtN5tvPLxojs8NKP
1TCvXXEVaCksdZbDI0xmu8FhwYkbAbVlXnoIIluFjeaS9J3vu4brI0gVmpvJyRn1Dggfk6PR88ju
s2vjp7cegwOatsa6WPuILBzNUiEhVlLZ/5X75EII4uxudAVfGXWxAqR0PJkXv4GyNTeSVD9AKXWL
VHGgPvx2cOHPhRaJL0R+pTBoxKFfLZLMayGYw3MBOfI0hOAWcjJV55v36/qdtWcIou31ZvufZi3V
2ebfNjev8J5N31ddzefyGd7/uWGrbbCnkVGERkVye9dr/Poj+UIX4bbEBJI1B6Ky9MLWqoyhK6FU
MosuyjkfeBmxSc2UVWx25H7osK2dMSG2YiyXFYp0UIIOq50RG07vXoxwKzXaxGYTwndjTEHDs9q3
ajUUetW5Di5zjIxRv7KWJP1EQWKGVvX5sP0IuLU/IVxQG3SLohVKXEk9t3JznWv7CKeC/XIPyolr
73RaAbVezCGzzRHHj3m3Tskz+a+B1lPFYCJZXtTc+L6CqtudExeEuV6Lm58eARc5RWiFniI/TBxy
Ln3v0cYqJ0tgoYKGI3vW0WgBX5kRgAC/VedOidhvyOWpUTs4sQwRZl1rSzR+3eJynLEIah1zlMlF
93BioMmYhSCn9tTkJpNYCD9m8f9s/+u+4VgdQF7MMotprXlz4j5mG/onztKXMwtY/6M8nqmDMAsP
utMAKzKmSmZ5qZ/753/qjCZmVzz34Si+xM8f65ui/wbusIvowTU1DIQdnZ3YvzuDnMj0PG0IAyUe
peDk6eMNG2S5JjX/zzYZsnFarMHErkBYir2G2e5b02cGeOcrO/NRLZMcXwzSndbTeGpulKa2omBm
zqsjMcvUEDRirhvTQXje/NnkK6Vp3catxJi4FxwIKN+OoWdkHDzBkMl9SWAN9aMAvhNcHdy7PUGk
1VRwsrwjUHAEWb8HX/KFGAIQIWC/hHQtLeBd5gd0irSyaFybR6DlIXbLQ7RMpRL3niROsNbBC3ab
KWGPJ2rqIPXg/TClNJz5Ozh+gDZGIwBtBE7Ukd1noGxarbBx3abVE4Pi8nBxpwlyDZwoxCVVI+Xk
miCIBEVHsI9kwsdK1qghtwhdJlsNQdwo5Qb3GJesqWUJ9q3z5MKPe3aOCG32kiTtAlXR/Oxq+4w8
ak9fWrRvPRWevGd1ymlgNBWw60aYOkzDBFEhA6Sa4rhU6tgRyVc0lnhic3s7+e/fLhqZg+T4isqw
V1inpHPUFMqyg+5bM9RJ5oY52kLn01U/oDGIuceptztLttid1Qe4u+g1skX4eM8G3nPkko4QInkp
DtOOcFTCIaiytTS836QUzS+aaouMOoRiumSl8TZd45BJd9xczw1shSWaI+EJ/ppcG4kfG8vMXEXO
TOc6HvYFpLbByLs+pio1Hcj6EVnhx+SQLptRRL4J7xRhZ/NbN95Xem7lN0Z073hU9JOfQ721AX09
fjfGjTSf1RIcNqCDmfPM9Aq7JOaPM1YvENdaKBKVhoAmWMY/PtHmqSVeM3AzmgI7e5fhYjgLXuAz
YJghQL9ax5sc7Vv+ZcQUHQS3lMve3ItcRHkVkNMXrFTrir7V/BPbMtUxc1c73bYXHeDbuH7Ha4lk
U+3qYng0wnPG9Nv3Nb7D0UkTL8RaGJIDD2XThjgMTakiaHz/wgvkhpJMKCsTLcNNgXbbjiJQdrpE
Ww1Quccp/X/ZdjozirIttV0D+hpVZRDT4+xEvst8e15eEhbJvhLbgxgeOIrRyfuIhwONlDaw8nMl
soLMD1pnQVp4u9KBulWnWQv2TIQeG/+sJnKg53ANnqLO6TvCGkSmQGX3U6q9taPb3xPZuTNyQXhV
kMvLxWZ/Irda/MjR6WmuDprOZbPgCg5iUqTulj1Zrvr/e5VlcJNsoUMBLL+drgl02Lp0AFROYpH0
lZf+z0cX6WSMa0uaRF8wHLBjg3huSW8seTVjLHSrKv4qLa1HPwwjVukzUCU9dEJvGeiIHYPC0qr2
mPlfpaMWxIIzNgzFlGnmYU9w983YEzUcDlxLt+CA/ANLKuyeiX2jlxvIMWLAIeDmfq+5XCHKmD3S
gJaGAASDf9nBKshaL3KCswANYam+YTgCGVfumtaAyBpmtl5Luk3kUgB2xPcUVGy5yu+Ap/SGls9d
jCv9Pt7wwOi43i48DUKuZ0vUpTAni5Q/RlmyG0mxVcwkaR9ouywSkFZ6J1S+g/qvjrPQNyV+3atE
MxfoiUVMADDrn1aBe5HWX0IsdfDvNcQpv4gaT67o0GrU2AF++DdxaJhHVWaii/tVQWo/5zHv4jkP
3CLtVT3ZntpgnwXxf2XYAgjLm4SkXLtgs3Z21sBegUE2iruo2Yi4PNQFP91OynGEPDe90N2Oj4AK
1kl61HCrOXtcDg92iMpkL7nJzjEN6R5N4jqhR2NIhPOGQrtkkJJkUJmUKt3Oufa+MkAcBR8zJxEj
dGBEJ8O8ThHXmi+9TlZ0bz8r3tYgnlMO87rzS3y2bXJjFHSYFaOEm5SrvKKrZ1jF98N3EQXoFTy5
uzXl6+StF9AzeNSm9rlKqkT3fWePdWOJ8n+zBXolFOREwqSeDnkFx+gJG5ryDEmTgpuj1eLNWdNZ
1Ps5BFDUsNmy1GEEyG9vvy2UkfyJi0whoKcxSayOdCGVksEe3uqL6WxO0ijPvyR+SWDQ2kzHw8lg
Qs+Mrcxe6DVYootKfq7OdC9f5V5a2dQoexcEUB3ADDWxfq3rVpMU+DdJCJIadSdk6i5UaoR8IQ4q
YiiPg6W1YrIjKYatj4ezmbFO4w5CBMYemikTu8t9xdQcmI0g8KW4TrXolY+3QNJMyYRUN0pPmzef
S6P/p+4xXjIAqxqoru1asl9u0ktb8tOYSzgLImoSHj4HDvEvAc9M4Fq/k3SSErccUpQdLzj33kEF
BN+OVkgg+kkHaonTwWowkrgFGBIQnFRJXEZpIBUSJqRqmTAPqLXRvg0fx8StDGzwvjHYX/yJ0OZ5
xDfGBOheeaCgMQY0wJS2CbscAfDTU1zofyyOEWTfBiKmQ0ins5sqEa//SLl3v8m2SYdbc4e7q+zA
dXkKJR9SoKAbk4cUhshNDq5kL1KDj547+VjjvZKG996jMKnv1FDqXk6KWDo2OHlIpNILu36P1FQp
dHmM43Fvb2tOvruztJFr+ra2hIRZ/bG6qmBhrdP7RmzBAfA+MhDqDMNDyBBVObrYv6I3Lh2Zv5x7
3cMYwXQ8jGQE2NbD3x+cCnNR+z99RSKzuOEFWfZTPimKUDoYnaNQJdUJuguZVOXFxyr7Tg03gcOR
mHkjW6ae08Gjj5PpJhiukIDX7/KGkQocmer/jfW7K79y8xsPFJQoIRTn80HBQ6kb9P4NhaCRkjKL
Z0ivtrnO/BovWOc9+hvYZHX0TaPEDDmAAGdf4wQTKEaqGSjojPDrOitIsSV7Tq/0xhWlD7hHt92W
VJGQ7ib1JKL1+SM1Oced1rYVXGX3KGTBs03mJjsxtKuJNYMVur+U+PruW/L5eihpRtWJCENanKB2
MhYnGTbqYoXdr6LV+W4UG0XmMRRwdW3BhVXRSDaJxgh5kE7JDg5Bcw0qkkGRv2sySqxMF/5fShvA
IbyhDMKctxD0pf7vsAPOC+mAIoRjQPdHEAIJr4uK68Wd5ks2IzTZTF0Bn07DKvgEuJcy2aNfoH0i
MS0wOWCKa+8hRLQxD3RlLE9o563N9fwVlzrae+3ug7jLCBI2ersluM6t9R9+rQIPgJadGJGrlANx
AClI3NZUkDiq+co6ei1ZlMggvQiaEN3Uuz1M1cULwMauq4sI0bU8Pv6rvoD8IcIG4370ZhsQzFby
Z7p2sE/BAP6NU/e4Y9n+NIp1UKbumvMSAabZMJfKrP+a1sZ8faDKeHfPulR6AdJliPZYqlaJSFqc
edDYurcAHK8FinOE4o3uNvzzYWue+hz1zhjkZdX5fzB3pawu7m9aZswtMXBKgXGg4FBmtsW28pPD
8gyROk1QZSzX1Y8I9RAtgQu7RRQj9MboFnJKmUB9g+n4VXH3q6fZdW1hGfI5ozdUTyD82xGY8DKr
ktBwup8b0jJK3JbWVDCqAwoYVjlH933k+knAcnSAD67j7mQaOVZO7H9xU6pTeNEYjZRmP82koSAn
EFHkbpTSQcoqokB3tDGFSI1utD/L2TBCImYmdyha+LYbWDRKCCh70ogDdN5pT1ajy95nSapjqRc7
69uDg5aLxg7/gLWPL7+ItizIwUGgxXFczc3HA83wdNKwRmX6wz89GoY2PqLjQaS25mGZOT+w0aGW
ySKNVAdo/J4B8723mZOSj3jVVSZP9rDcrBcP2yP73wwPXDFkQ9uZfkwzOkTdzV70d9AcKefeqJ8v
pBlEIxppyGRNvj8BMuLHysaZFMxmMwa7CzanlbA+atlKu5/cqDoIEXuArHsBe0AWGCEp9msaHJ/E
LJ+MqAFhQvlFK8wqE2Xw/H6QJ+onChrKlvtfhAG/qDA9pQjb4rBzO4nkMAaO5i6+EjBLXS0oKvV1
Yn0RPq/CTdbpQj8xJY9Nn2LkrvgZEukW6KxCck4uRKfXCuEH4c5qVk0iot5CKlTKfuPmsuC3rnT3
SnZZx6yRBVBTcyHyZaqWc2qoyVUYokS2I6tmDmrBCYVLgyVDGr5ntj76dNoYGcARPNzIUVjQ8PjY
uDldsmeKnksMJKvbAW8iWvn+96RuRZ32Xxe/Tgz4gc6CJs96ujQs8dd2jd5/GgLJMCBCbSCkoooM
yaIv+x1YFybyQa5amRL5L5TFMfHUVwVwNwIyTZhJh7FYtmh2ylW8f0RUlgeeWNTMZNUypjTxjh3U
IAy1lZ6V2iZ8C9oNdpEHfdoLCI6hTqRHzR9ck9gl5ThrNTwOy0OttW1a8LdghdvgeS+/zDg+OWsW
GJ8dBWMACONwU9WX3maOkRjoJr0hoqlyOKkwygtoydhmnjZk0fGuy+dJW5FwWjFUhj0V80fwCug9
Un1Etm2PK+rUifkGd9uk50VIUUXxC5SGG1k+FOUqOo7SdpCNfh9RuNuZsh8+xMySC/q1DLt90lWp
fpTXZYrJKHh9piyg/TW54Nkqgqc1XdEDW/C3vi/EgQrz6S30bKqxlp0xz4MCnbAQFC0wllZliFbP
GtagUJ7Z6RI5QPPBwYmfKUOJ5ZWy3zAp32kw2bgZJ5Wd4HViEHrFPM1+1L5SVRpZc+SjscQEWTQ2
XvBYbyG3bRR4sTkr2ijwaIYmXhGWorVb1SJlFydNQC8Lmyy3s+jLNSmtaD/VDgqfAm2+0fSpUvN6
SJ3AxjlUcbsohYYNjUYCAKMNAfuZbHHnQuIpAerZjkzZWk6gELqss7HNnT6eRpzTe0RFFyD5qS0v
QEGPTaO7A1Bv0MFFsB4a5xukqC/QyR5kKOxHEum9J16HzdNoZOK42SGG39JMbXQIGYSKTkc5iXPo
4mk63mACASIVrxTzeRElx8rjCRrC8KyGB/Wl5v26WRbV7r0ZvBiL6AeVxjfJ9qFsGgHnapvWDRi7
4+nJY3zhDsK9TmDWtRKJi67raJd5XHCkP2G6aUwWvmh2HlGLY5tazxBqMhk/zN/ZwqNPcLVddOdZ
9nBPiQf/i3Ev1WVcdGA/2I7LPvlxPLdcYk5egcq4GakNAbU4IVKI5MxFFdobnWrE92dfcFlSY1me
Hye5WaiKj7X907b0wog6k9+2jvUizjfJdFJkMUPUNpTIut6mrhXobvuAgjo+rKswQHDX1FBDYSVG
VRIANFuW33CnbCO0W6e3U7JCsxQFzraOLke9n+yj4+9v8Cg4GdbxSDWInvgN151BYsbtCXOVj2T3
eb6N7ZTvfOMkXuFq7oLwrqFzV/CgiQaG0JlqUjLShqElFP3FNwYOh7soX6rbeYOlVgXUskce2Upe
0dqo6MSLP7oF6ub1h5+NnBgLEYL3tO8N0GmsJ8/o7VXCr2la/629WB0256WLJQ/B/xlGCy34FwOS
II6mHvJayj6vUwfX/nFN7NW7HvLg4J9rZNCXeJQlRZGEsZCdh9593SSJ2B14UffIRhr/B8QNskQH
w3boN4pfNDL6szHWzj0ORAeBati1lxQcUkh4uLxM3hV8fGC2ZsNwvO25AMLkN+bCXhxuGVHJCtdG
G67CRws2jK3J2XLyNmo+a80bRSZaAttuL+XiPwdj3N49E2r1FLXqWCfaTKIShZdpO7f3y8Buw4jt
c/ATmQAyK+CVjrijAeOjWwgpgniTjBjo7JkR5JMdy0eo+3gepKY2UhXaMxPwv4it7cSpOIBuHXsX
SL8mhwgvFKvglVbz5nfNY42QC9XoAcTtphO8yg9xyn7ojBcJan138rwQ4HHgP/xY6OqVLok4rKvD
F4p+bFPmJrmQQgW9CJSK9QkHH9cnwFZm8GjNEAXklDwBIFwfv2zgECzzYXe6ekTxQENW/fQ5F/8L
XTURLgnxrR6IHZSwuVDKj4vCX4hUg7Dv0J5v7WZMHPRPmo0A42PdcdOYaeS3BoSua+JxMRFTGJUi
ZIaMbCrt69PnNB1tihRQL/krTSCznpoimhbgbMwOyMlpo5/icCKKLon+fgFr88RmlWFdM3av6LUN
Das4x58CMPIElmqL28QydqipKt9mQ7MByNeiuU2X6IE9F3l839fbKuEMlD/CrFxUxh86LCWekH2B
orXzirfVXtv2NJRNVj121QnBOeaK0KOpqowzHrsYLEVY73IQWWLACiGqWs4eTs8WqPEAwQ5NE+6N
HQm1GDGLOyahbnkyJAEyVIKLzQ+ZfRJLZZR77iot4tTEA78pDHrF5dvYunI/hfReOjaFQYd7Hh7+
DVDhEMuR9WDmx1Sxst7/eZaKwCRKQFQr9+IcqGM9YJeBcZQCMxVr1RXl/DF0ewZfRWJqhtf3+Rms
AaY9UBBV9jinxALzC9HP7v+4cY7GeFdAYeuEXexk/cWVmNerV5mLf5CNbqC6ngrgiGZDg7T83xyx
5jwzeWUNRoktV+z2N3q4ngz7cXbwCiAQNlfGTP2yusfKoAf5SE+a0qHnEIMloaunL4Akuz+vEbZr
+lhDqdd0x+YA63oDnQF2QtMNmoQ6Y29YivhmbzJA5Fq0EeUq//ceIzlqdeUZQJgQ3LLfvgr8vxUH
WnQfAZuwcB3ztlWuT4Ep6UBQtTnicO0dfbcxkisnBtThKH8aLg7f3oHrtMSeZayrXA4qbfzNdHcm
z/dVPWex/1gNuwscMKwctERr+sfX8t6ETDZfSZwDS4mVm3fMpDbEk5AQPpGwrZKgHDP5uMMOPRK1
kt2yXHdZIaAr+dY9yjdFGQebYjLPTlqMlRPXuNQMw4ye0dAxx3jJMzVntaPMMWKlDPEE676b3NSi
yjkzlXmh7Fq73f5U07SJTCRQnJafqSwtZab9Tv6k294ZurFXWxPtGE5Q6A6Cn12h/2KUWD9FMbGM
sdj7AgO/Mef0u8jz2THBtLpjUl8E+Su9LeUUBIY844MsrHCskqnKXMxxopTul8pz4hDDjUo6f8LH
QHugv/beOwRDiX55x2ytcM1sX5nNs8URto0nvtG1p37suDur7pahs+Yeo47GpfgX9aIWtbuxuPzf
V/B9PvC72JFh7V3AiaLQ0K/V5bxqMIYCobW5KwcSNR+a7xkl1oWqn5QhJqJsZxLWWciRl5buNJAn
og1h7O5q8lVct4f8CfcNzm/XaVvOIIX+gt9ihjGHuNV8NZQDOfE1Q5zV9HL0CFinPzVQ/uh016Mc
9C7bl2c4F0RmcEV2OTOeu5Cl4DrEH0LU7z2zANCcU+qNJ+ZccObEFan7xalM+glN2t3Quq99wYel
kWNV9zXTlXWHcef4gZV8irKCPLtPPu3GLuQcwKmN7ViPCAcPbWxAb0ebxUjqZBe65UsrvNRiGH6m
z5YYF06N8lfD8JqgbOC7qvNrH9wwm1Yu3aRkUEXSe/DwIptBTf+SgPOEOBkBbomxV04RNq3GrEJ1
CvHHjX5BPXe5l+gzwc+OlIOClSDaOYdhP1SSQ9Q93GULvu77CFXiRJLIMcxZMn0s4yzxuEg6fS3a
WE/RJc5h/Lj9sVSgU6DOzkIGL6AP6Ra6MdYjY7otlTUulr9jQrZ64tZl8z0Ce01uFWLC9upqZwXL
bI6GPdKOE8d6X0u95xvwwCxctV7QNKJjWAnAMG+o3jfmp2gnwUVK72vRg7X603mdeoOuMWOlucqa
Orm86bZD6rowAz0obPvvm1/VTouJYI+NlkuzorBTV4eIu245MHZVQMIaoazLAP6vougQfgMc3UIg
lVtgVUvaRBDEgCfRKIXJZ65/iDIB/YkwiZSgORumI+HoIHlpNDVEfT1jV0Hxn+NS0juF99mIHkhr
1n6IExv3/d2oBoo+HDY2wTRPdpCwLsWyZGszBq4fZpHvFqm7tagjbuINfBLDo/ZhJ2FWKno88cBo
zIwhy13yUjAtff8n/hQfV+00RC1C6uCcRt9qmTMSomVa/AX5O6f5GJ7Kf7hWZ9OeSXX5HUpjDh90
4fiCpilyKEQp46sTEeCIaYNJLpCGvoJz5kxHiiC/g2DAELFBhR9Zj4OAl6No8YkI+pYOvmS/an7J
+GQOo4UEE3nJ/jtgniBqtourcQ4M0O935zBH3Hcxd3LI08nfgk1qT3gyLhYFt1n0E6YKtkPfXt4F
RfZZFfaalzSGVsWXn0MQJoWLUHSmkPZN7D77GXGan6rVm7c57lk8V61xTkjctYNDvbXPFM+/gsRU
tw5w33RLDTH5b9KyzpC5Tkszbi8ZYWz7vNA4bvb8RvYUgZZCWPjSjyuOrSo0tDfDDSAnx57P+lf7
ZGiBwA8dpyscbo1wASZb5xfReCP0AtGc/ZsRKXgpI4YdtpB9yNnDZxO2X3M1HERvWcemErKI3eps
DsxJUzHZFlOBdde4qUF+YciqTVyfKJFKv3FSYrrKq6dLzmrh22h7ssIh9RTWoGI9p16bPWiFAlNZ
IyhUsf5b4H07XzvmigesMCWhfTwRz03wCgq2xU3UQOZJMgnqa7kRcXt8m2Z+y3PFsgRKbUbtUAU7
GR648jAVcDui9U0pJcMhYlxrFf7AD59OnqX5jFOhhFNMmSGfAtFAXxMju7bmyD14wXpv6o7I3Hor
mCRXqiOR7hZpx9BtlXoc4mEoy9yeWKBJaEjPT+MAquciwU6XUcIgh9HvoTzZrerDUFiUvgyQzmD6
/1NepE3FWhSqE5ULQND3H8CBQRkS7IWMECK7asXZvJoLip/7Zh1Opg1GETBvQqNr1CIRWCBUdJZX
OyrD0uInwx2g1b2iC3BGzcbqe7lsufGJ3SQ1o9MYc6Me92HpLRdf87th1DDciGnbr/YXbyOd5Giq
D4gf72PlxyTGR8mc9Fg02Ob9bqFuUrjnH5qQ2mWxgKovuM522m6njmwu9D3CKhcQuKc2l4Mwa6RP
ujnxBP9rSA8zUwLhoit2OU8gMYjprhzqJXsDAFQDzLwrYXz9XaF3lLDEpYoe3kN34zjpUm71zDRY
3UCFv3e9sWVZgTYD7Ho5xtjHiHeizg0BL+TNmoi7PkVm4Xz/8U9sOzmK8ftegSI0KoVswc77t/4S
n74x2EDRuaTxOMjlfgWCdvBIY0G+ANCrTZ91ddjD/VAGBc/CfCrgiWhnJP0KE9Ubk7ER1d8X0d1t
4uIPRXM6gVNAQ4xJ36UTQxa6lkhPNgCRFAjz1UPuMCoKs5zSF7x7Dn5uLryOtJDy5krAw9d/Cwj6
hxzgWZgbkoPXb7Pqpu9T1ObeOD65dwS2G24scniQHjsGazie0XPxzo3Ar0Zsjgg4SGvK9n1Lgknb
W+/f+TQayj/RPw3yCC7+BU2+a7iMH0Od/34SPucjiwJQA87oFNaUegMdRNdbslnrU8GXU1JGUufv
Fx7tXMkyccU6yVV8n28/v0EUb5bWvw8d0K1WiJ+iVRox7ZyWu3BRL6lEoTC90d242kKw0dkMgfKf
MZQmASWUIe4PtYc1MWCcPg+QxAf77pv+RVfNW/mWEyIhi4Hz0o2WBI/qCuGR+0e+4LOpIZwDsMUI
BaGLYi1x1311ciDD9F5uQWRMY2GTs8GmPoDF3QqZCRgQy7Eo/U/aqhKwKXxJkXirpYzH8hpgv57+
oxteUYlYpXSM8CCeEp2fKtjzLF1aGAdoVN53LgU3xD/pNYI3mfjpBJk4AWictBwbv6yQJj7fHfXn
s38LKFSb1GAm+TSIILQH3sJs9crutVngzT78UaNhy5jVdrVxcAO/QZ332oxtzUXtLBGBUqfbSbRg
VT2sNttYlqayk2X/6d4qHcHp6DHXmGTin1cKECWbv9DIsmw9MW2LSr3getlkLhEZcOMK/NohrPfe
5eAHSlfSbCNFQ3adDefXOZqKDVD7oiPyEaiIjKlaK4+K3ALR76y8Tb/mTLn0sZbsXoy20gZ69jmJ
BDbYG/0r2RH1XvbyVsHJma4CMEQ3KFw8UWh33hSYfBD4vJuEMKu+H041O7b5kVaZkIt/kuw2M2te
kP0BvxYprhqOshqlEfnZwCvoD7JZVURk3CTi6Ropt2ddQQf8Vv5Wz+D6XC1/VEZm3CSkFMe4A98p
x4sGhzI6UuKM2/gpF/NBeDbGwqEPIzazxnYEgjs05E4mXyHcwBPYsT8yWzSA/B1ZFdWxSWvOqP8U
+Y2j6Xdt1QLOfrCTNcxhi9PgCMe+g/A3s6PH6LZfP+IgvQ8i2AZHaf+UUNroC804ko/Cda5JEVrK
VyXXHnOFfGPV8o28v3ohlvkPS85yWKV9wEUhghcyX3NBPJBOis+pICdvBq/7K5dzu/3lRRCqhja1
iA2i/pjauFH9SOqCtwfXqAbETnIxc+UiAyaTAu0+0WFWYRn/JcwpYMeEZpESaUyEhO2zcYAciH7M
MzPerHaUNJ2uGHlLCp3S+wVtxK+C+gzxBf2hOK2Ma3T17XsTBRatKjx11fMeyUr7qIINgmpjf9DU
R6VQl+fScdVsGdplSJzqfvo6dGeGY1dwRCaZI5Fwdl48y3NmmzRQIrWF9g3ZDEvkOVmfUVNY38zc
TLD0bf9COuWIyD7lSV+lyrVuV4gfnPPGymxijyvvhWOOVf5VBhd5LjkGh7ZyJ9ELhvUZS+vdeIss
ZpnEhG6ga1tLXgcnRs1anofW/jxyK5NPAq5weytELU+kd4gCasASVT6Mi9l8FBCa3oegBwdkkBJM
JCivooEhfsD+cMhI33UfKQHU7x85i/vWFk/HD3+SG+fUsWZaWWCvbBYyjI+McDXA/RX2SV+CWYt2
hY3yAldeLzbBQw4q9DyCNRbF6URefyQ3qB38WgVVUFktDV3JM9spbnYeESdRBglgYRg+UpWtPPIw
jNBtrCn/qn0c1HeSZdV97sbhRG6SEa8nXkGnPhjDubnGSbnF0+VGmXpietU+ZEpGGKfD872S7JvQ
fMIuwia/tPTy7wixsmha+gdTzUbP0RPJ4FBeKsGwIwcedvJdLRaTXQjd1P7Ka40OKNxsUd/iQhes
c5CI/VzWrfmml90ZX3iUZoAOk83nDEl9+LTtIdQpZ3j/BAcZ9+wCA+KhmBjP9QKuDTZUzEIEKSts
Aaqa/UI+PsoULU9ftNe+jC7WgSsJ9ZDv5ZuHYNQtkhjO4B5eghCkJ9gd9g6y+7XTx713fwK6Yao3
Fed9+avB2RdHDdtkn2GtRwnic18Goq72AG1SbNxERVx5Ot+qM5bS4Nk0Ou/+ST9+scm7Vw3cFV2B
C8AG6ovrWGiR/Ud6j7d1py7eWb3Ke8CO7aEBw+FZbXhKTAJVbPL7mtd1zXOJDw7I15zMwkCp02GS
wvm25DehM64iEUbTmeLun+mcMMq9xJ0OHrtpQhPtHK32RyOvhUtgrKvqoy+ryjJLc/e8LfbDTY4K
Xwc/qGjbcaXnRP+shopPiskET9LNrGCZDcbqQQhKJAtVyEsePOuS2aP1Ti9p6pC+26sQCfbU3YZN
91teQc61/XKu9JccQsz1ta/KwI71RWAoAPVPqrDiUXMzeI29uqzLh+dUIorz0ndJKW8llQSITQlf
7WVwNxrVTyA07/MxMje0zC0IO+ONoTWOFIlAFxoYIgQHFAcKW8pWzAvh7sDNnIZV73SEweLdiC8p
Pm5srEr2rBLC5IeJWhAoXiA2PG7jnrnksrGLNTbBZ705ye9ketyWKegaamG4fKRsX1IgMXrhJMem
LopYXw3AMGiMjUxnFkifL1oCIqWZVn4UihYCrMevKP2qQTeKIepulaaevlVz90FTnQNo3fhdtAs0
XzAgjxjkqfLfLNgOXGbVTCZNpNJZIGQ339loaBBvAY+Z2cZbI/SJhe5q0YItlLqEeA7y4n9JvrFN
XPGe0CAjCgcOiVO/WgdvbQaUS3KeP68fzDvPDusgxupHq9tDKYlLwrOzef49ecBtgrwZcGIIhCjj
2f1q/VOtat+gUvSfHckqGQ4oYSOj/2ieCWZokYvLJ039QUEaUdLWfy7GVS50LmgRfi2ZSf8dknMd
9ty2tWeBTp5j6EI0+S/YCUDqD2bHxsg8zf9/PlDIpEsQqgTrqoc6uxgncl1o1twsWEd7tuP0QzTI
TjG2+uOqihg1bMkPx9F8YWe+J6/1FkgVLqn4LrHrPk3Z96ZG+YpsuTYZBSY4ELjB02mR3V2ghtT4
8B55Q2CVy/PCRpeuRbk9dhDr4Ta5pGN6Pcep4WIP+LWAfxYqnSqpjV1esadM7xB6lY8aYopAydh8
Rg+sWYUBfXpMNvhh4LRoaxmHZm8Xm004bmePSHw2MdK/KrgfJNuozrcvuHUJnSpsgOldivJ5bdDz
w0QutjRtRYlg8u+gt3FqoZ0uBagdxH4Ff+mY7iKzhHd5jrBu0Gv6Sz+fhMwgzuGv0zBsOKltcdDk
P6jll2/gfK9bddMbf1oNc16MD8JbEPnd3bbMfKXqq1axFxXIemCbEajzN9FO2hbGH+y6HnNBgXg8
rZzoV3DZmt5stmQoF9H7H3b8/S/kRvbHQaXwkS7pZ+6/0zCfXgT8laPDuShLj6yAYyVDRMKKWukp
H5dMn+LH7U66Kh2FIp/GrwV+hwaKMytvrywcN8QhDO/Br+kqVlfJvdqVyePdezKQJfm2/dnde5n/
OrYqyIcyzW+Hs8eH9k64qjIbJNMN5pCBTcZkVAdS9/CYYyNTTm9Kul0M+qE5iQ+5SV9MxNZ8Nb3w
WxqU4ly+dToNFPwaMAh1GjJC2ylnVH0jc7VuMH4pHDFjJ3liNUXM7srOTllCx1ETiTFhZxK08Lc2
105qWL5mCkoBwQe0qZWp64rGHu3roSmqufRx0DACF2G+fIkeFTEO3rPumIprmlg4yLkRZRAuCS3A
DCXkSlrvr8MgcWLjS5WVbv52UMlnZYqRab45nx8ijwkZPxLJbdcoHq7nRauy59xJupMWelpqqoWc
VEY+xnby6TCLdd4/cxhMvC1Tnsk9+PvjYU3FHv6CKYNB+cY8y8S4EZtHCwHkQ937IAiIJmk2SFQZ
jQGqDpuKxC3Qo3l17Ng9FJpVNk4gpjf7eCXfxFOyhEsHbAqVuna3KDnqwH6uNDLBgxId3AkT7XRv
Bsp/byNs9P9H5Kagjqh9UsqzdYxUXQyOYkOxiLaZCp7kuXXKRB0PdzbtvX6LkFn+IVhveIWuD0nT
LOdDmpggM6q1SdgMkmRfbQamGX22RP1eouIo9nGZrh08sD6lMfjav6aquOpjlwuZ7pIpNAAL+Zfr
IaV8jvBj5B4PhAtGmr3uTfUqCQdPiUjIIjbBPTms7a8K7hmcUGfCFQ881lAKuKOp4aUy00fXf5X5
mmCvtQ2QeOq5cnoBLOliiSFY3W6RHX60b4jNBm1GXpm7LttjiXbDx/5NqGA/ZaxQllNoA0LWhcKI
ub3h8+A+qKYRUgZzSTb4BXPPdkqtjdcMtE2SB3tqrdKOMmz3q7cHol74JlXrHaFLjMIPMbukF5wv
Id5ryuEfQhDuv3cIDSpWvu4yaNSSisM8e7sAGNT5IZJ+UTkuGQkOI6kAuDNGOdIa3Zgx5RA/p9sO
vWg2uhdGx0bqPI2h1Bss2yfoTbdP9LzEyNAy1MU2qsc0zKmiBfGexnS3AAxLtWW+BlBv3UWFDn+O
Z/a1YGOTJcBqLYTv+oNFYdtlYRVCk9nv6YWkwYGKj7+PaJgrTt12Mxub/lQL6m2nGSNOma5ymMcL
I1GmYRFxyotc5PhEQk9gBvqORijn3tWBQj5iIw+W+nsKxK1vzFKX2G5AiwAdPGW7sfrwZ9rx93q2
uDvPsO/vZKKDsVVpH6ELUeyFz4SNMDp/XSa8UDb2C/PqILccfYZ3ZghDBJkDmP3D8MujRF9ryb7K
1PWS/1b+RX7QuNr3VdCgB6c+mIcjmRwOmN99eLytC/3whMtjKshRPDX7fU9/bHiXiKT5z61U4J4e
4EiMFSR1iI6AYeR8Leep+WRXbt+RA5ix68jy3telFxyKwTQl9aB/v43+yveYgXVSt+TJV/dIp0fb
1QDjlKkd4B57UlK12t+XSlKbkfJcNlWpqSakrtNVpNkteAhZEoHngCAmfGxXdtbau9sCOyegw3Pc
WnSmk7DCAw8Nb+CzVDR/8YUeEtMBwtnSk9TzjYz7hZT82/TijMGNeM4/YsTIOVvl0usu9Ya9jFMw
XLlTlteA/vkRKvtu4Jtxvb+Pk0JssDzu8SVt+6hsTSiWTtUKjxXlr6huJFqaDIcyvAeRWbcCI9OF
hpqSrMdr5AMigV0MES9TB29dsc4aBFR/K7h//lBohrObD/vZaLoIWaI1BdnXpa60z744A43CM+MZ
KH89QUbRf4mnw0DVXPbc6tEkUPAxhujs7xQT1LTuQaxlrVERB1wZ0qQX8DVC2N79X1rDVjFuW/w5
7KAB0bLNR5vIcGo9K8e7KSnMoJSqIYHMBbmYwTRHOxnMPp4MlRlXaSzlBO8Cj9H9nbt1xSBX4Uhz
CZJcYloMHivubnb8EKZtQOhjdhXqCrEJvpdN6ehbeuz4+MRyYCa/z21vHRAfyW0eHzHoFy0h7vhZ
6LdHBf/4zN7RUj4qT1g0/4S3JoRlJ/xLGmGHKd2k2nmVbhENF8loJAFLiwXTcfYDy22MSxyA/3Pi
5h5u2wzfHcqt+8+FFgt9L5A92QpA1qd1lJdzGVSy3QAlFa3PJKRmqiXTYt0vD/1i8a20uIvCPB9p
sLKKgw3CipC8U+PtwKDQcARMrAewuoTtmLuJ6hP3ncANCTroOT9kVZ1HNduW7I2hCREXxUwqovru
lYhl1zfOPJ8/KjcELoV7902T6fFvNG4NRR5E1WFCUUYMnVzQQD1GqdBHeNTMkpQAL2ctFzsZcZKx
Z5yTtlDU+8V8u5153GoPTTdWrYsmMLhv6OU0G8ywyC6Hafw8tJ6aGTLEVUm9a+jImo9NKrgY/TQe
qxwoRQi2/A1t8ZekDGjwo5LohFRhMjBuzLG6/0Qms7Gx5KTyhrqHVIOOKXwB2FEiKN0njd9QlBsN
bc/cAV86TDRDR/MMlofpCvU8yA+piDIlmV8cmvHWyyoSV0vzC8K9DzdFEFWoVLgJ29Nu+jMsZubs
1HR2Sf5dKiwg78yabwwvTOggdHNyctbMxr3zKwRmkjCGyzeX2FrA7O2hGyo3e8EcIiyf903zTUgE
FSRp1TGIfd5D80kcb586VipHkBWCKqGzxtKyQQ/J0mRrrSjepQWeiARMPOKJ2x0dqWAZueINYiGC
KCEejMPNv4rxbkvB6JQ3ykH9z/AkmQjPEq2fHNM8y98plQGyBKFa30EobNr2HGUFUQ0J8MVgDjHO
FYJJfFMvxeYIEldoy2u/c8+g0O0x1YvE4McM2ljo0EB71dX9Ymd5t5VaqjB8dHF7IL+EBHgEyiPJ
pRh3AxwnCPdVYjZCnpAE0SCpRQR6MYMO8mGJ4F9hCxCEnAVvdgVffTjZRw5lMa/4QaK5Gc28lrc8
SklPp4OrvoAL4nX4xDUl5+tX+LpDSnWahiK6wJv3iRnSSsj9zE0Q7l6cEHGasPHQedy1Wk/VhO01
YGBVNQaWwXDeMFY0m0cw/uTAsM7wd4/mLAwypKjl++L/EhmVfGcEIXZkyrVMZAGzyPrC0La5HxLj
j3GgTznZ5liCrNbN1esDsI51FbzOyg+b6uRWGFq6wt52gbPB6UmF7UKeHcTis/f90gJ+68dx3me6
RzVVVmt0EjIEuvpUsBi37TKuR8h38ishZGZFYOzAz16M/BO6LYqvizPZ/DkaqTfqKhC7giWxx709
SVDwKVOEwcG4mvj6yupjUuIv0o0wkGqhRzxYCuAMe0npTaOWnO1L4wKMAo2e7Tfkp57etzSbZX+Y
7bAbGJ0E18w+meWsF4Wv7Ywnw1j4CSg4xQRgGYabpl0c3YNQ3J51w03+ufaXEjIZkjHvta/amKeu
UlicFIRLgDxqKBTjBlkHFk1Y30IJxuQrFVWZYN4P43rU+dRgqcJV8XGR3WdK6xEc2v1XXbCwGrh5
SK69bWM/pIY1Bl0szH64CGQMnhH0Lxvacry9yFEBGAU4D1BOik3Fru6doGVBdogzLGDr/7DuffOD
kclWTbDyNjxH6dKFfCDS5ctzRpBFMY7Hrb6Z7B733NF5+xbh+hiDvEZ63OwfZdSvjFfTqxzYykD0
DIDSkkOFxi6CRcYMwtqSKVq62opoZOkHLPumB6fi8V9biDTZBqt/+v7Zdpk6XanVo/8srvT2CHDn
lAEvJUvBpxjtPf3F6YZRbYiXF9ZhFufyGvlR6ylEBHwNNLLx4fK68IF0SUNglABpcP60M12mNvwU
wCfptoyPRw4F5GfUIgLrPmxXePbBy2wIQ1oO05xc8/kWJlXVOHGiHGoNbDTSbNYI/FwFfg6bn5TJ
TiOju6CnUxixDM5MUfX3FH+MIvQYpUKRMXMxt3Mx2U6YymY3V4QZr5KMFHLnIOSwkZXn/C3TdJJR
pKB86qtKxO2oquU4zeEwLXtQwpE9uXgd0rTUUOvKI13CLz902EtA0Gl2a1ELNmdMZLSmgVhPAWP1
lPywqorOd6XT2F/iH9nGRlPou9UA3TdgkvMxTlHHTjKKbKVzuNExMeCK5xdRwsoSXz/zepgLZIu0
c1ypfYKIMcplG5ON/Aqjbix3nHO7pEPOk0EQ0Mw96aPeTHfi0X06bMAlX9Lcr7wDhs209dwoHNE+
djqEBFwDqxPgKC2Mwo7QWAv5qCHQp9HRh+PmhSp98Lvsdhg+3IMOlKK65T5jmb9+a6Ny3yy6vHQW
qU0s0IMw3Cil1743DPOuHaKDkzZSjQG48XTsqrt2DJa5/3Yb673Ov17rzr1+57PPyBAsru0Sv168
ZLPimzZ3aLuaSZq/RPU1/Wtih3owLJETKmYYgVukQvdu1/JdYS9N47vwXe14Dfhtf8Taslh3nTiB
5h7pktidBv5ZR5WzhUDvEDt4TCQFLKSBvqJX4Fs11FqJbPguEQ2P5qzlI+a/W+ngVevi4RMA3CPk
95QHRbBSsqPkKEl1M7rypHtX18+mV26OCy7Z5gO3wqRxXvh3XS14lwKZGPA8QBsqpvE2W8legYKa
/K4xAiLUDt2y1TV6fCxY+69TAZBGAKdyOaIyzI1LWDN3aPAQFEaIqBZ+0x2dupCbyPMrXORu/rbR
UqFCKxQIpAXzfFHzAnFCCkrrEn6hGjAjfaSeaAvfaOqeaGTw68mCMeQIlGLf2gH5e2YUtVgncGwE
K4xO9Cs1jUNR5u+Xr3IPLCPEgQV1pTIpSRLHuBUafLhkuCnUxB4Dr2d/uF1azSFlpdXQtlDNQZG5
Oj4UOpA0p0LurkOK8efj4YjPZHyrCP2e2gIj6gFju/IoIG+YKGwHiTZmTR77/qgtsYvM/ylbeB2z
yPswpcrAK1gN1nqt9kGytGROGOrQrDP60HPIQqILrCmfgmujQe23xo/w4Mvj29/9PM3K7RBV2Yh9
TZUyvlcVoSpQq12nC6Vv/K6D/SGwYuzGBjjvcCcy5oNUFE7jz5f0auokrq5B1yMRPN+1abAK7CW8
YuVS4obzERW7M1Kkr0lDT+g4AVFeCcQnbMXikLtred1CR4Lq7YJ69LSPxeIEsOCbrHAbowL6L52N
DMr269fiJJhvhmFN/NuEiwh82pyogK5VwYjQJ4OwemJ1KjpJG7Gewlu8QbyAv5WYhNbOf6Fkats0
Uj9KrpL34lt4yIAHeuSrlPy32nM6pjuvLvj/8scXpIsFagPpn4QpJpae4R6EtrvEnIfzVliw21aj
h/lxOPbv5EyHvrNCWlriNZXv0DotCGYUFiQnpWPl0ILz0XQxngnACoQvw28wjwMyI/JQSsVOpSVi
j+4Bg7vHy2rfH/PmpJfMgPtNKmYlFSz8K0Dp+XSZVHlM/QwL2cXcft4xEKomJPL6aP22Le5t818j
IiNFt2mhzy+SWo0Rh1KcijA0to20VTO5rcDgxyR6eGzy7InMqrMKf33Zy8CNUm9wkEpmqbba++q7
V8KeVAHOyOKHbwSH9UOBNIwsYdIV2OhvDU/3IovKWoV/8++rBuJYEl2OIIQKLlbZwOposKP88yzS
FkHuHa73LTZgTPSDqMssttlxsIHn90vBcp5FEIzCS1T7RoxlrCfVutjSFl/JE8mKMomrE2u9XjP2
ivfQUwKEK0KBhbnvFDU2mAnn06UGUwlSKbc3rKANnJFUtT0fjKhCCd1H8FmX0ZC5vU5kcoynbs36
YV5nFblrDi+IwFOcL6iWA/BwB08kXBQpTFWd5vMQM83/oGAFPh482LRamnjoUqMLX4XtX5piprFg
uEjyXDqAf9yHXfzppYKPfaM3YMzz5ALFGHTJ4/KGOFefK2yMDJxc4DFCwgj8uYAQkfHJiHjWUDLY
xV/zRtSuIgOODJd+BPz7RvivbuorQazeqM6/8K8mw6l5Fcmw4CLLVmxsUHED+eOO/TGQlCcsguPO
ifii3yIu8YnT8p4ejQaj0LEkdJkOJCET5wmje2T020UBgdUunzMkbnsfv8V7B1jGkNnKjorsYLw7
/vTYVfuJsqMExtiyRNr7W1ZIGS8WteX4V+Q9zukmYFNuK41Gr5RRJiz1gAmK9+YHGckhQ94bzyNg
zRirvrXljwb3kxUmWmff+/hWOeq1MLikooHyFUbPsS08hgZ7EwBWO1xM69jXXHRqTiwZIPaTnps6
RkL4lLPdy6fHsn2bXvPEIEuCMoxAWiol/NGvUJ4fZI2LvZe4yPr1mf61SHDGbvNk8f/x5SqpxTL4
IkIIoz/IRwFZc7p2hOnF8Cm6kvy/jxzSaq/CEw5Lmw/M78pveUsy0hSXqI8u1vItQGFyjHatq05b
YtsT+QcgNEgBsjTNCQ7YD9zQQxHMAYdQ4Z1EfSMJ/aIONzP24H604MAyvoIafef716hDuTw990Ul
8fwizILyyOCE/oAvrxfkPvO2qA+7RIRJqHigUeWb2bsIlGdb6QLLTlxQTHg2iZ0KZr4fjiOXQB+z
of5UsBgewHzEZimu0Mrj1WSYjWymCL8nZLE0pQK4dVOKWJHhm052kQmaePlE7u/3YWSqqy5y6IM0
IAjfy1Nb1ifhEK1LTpw6V0Y36lrQ0HYdQ4xMptFm4/7eAXEGX5TSJ00lToAh7OdZU0UE7cw0MaxY
HT4SaVUbhRjd14r4EruhODV89awCTRi2qJLndWlyv7xebvr8/+55fDTDSzZAbiLi9JNYwIa93csA
kuPsRlnPNpGyudYODR91K9VjlL2iBmhh8THni6V0C4iqavgto9k3p3QYSUHxhybrLSIJ68uumOrV
xKpa0TaRH/6GlS+S5btxZ+GCvcmAvbIuj9IN+QYsHKWGf4Zg+AAm2XlKp3mUV5ZnIyQXlHus7l93
hLRz/QXeRnL+JhPM66x/EnJhB7N/cIwzOp4OARKMW9IxJyiXgCoObdhz8t/P6uKdlDzOW6TUMgpp
ag5FBvSGv5BeXyO4QomzzmMzpcVJPJbbFf52nB1laMobeskr2IQakaODeOjZnLyjeeom0OuG6n4w
HtfufdpqDhfJ1J/pxArCn4jo9Zr7+6paKWICa4dVXe4ES95bDgcvjknTNLdOri9FjMO2ao/YhxuC
tCD5DKkyiIBZo+h0goNSg8QG8x7LXxejUs2NPZa9PNFjoD+J+IEJ6NbpuXLTc0J6fWQpLnmQhIHj
CnRiaSFNUkFnppVNUFOKz0l55Q2VRt+vTqQAA5rt/skJiZNPWFNa/yXRWGAjDHGPxxZzI9gG+BHs
TDaBI4JEKCzRL/PsZcnBepA9kQSa+tZN4OA2LyfNHvHfO4b7CwW8Sk/5KC/yuJhsQGSxIjB1Ia8B
RzX7HAoft0IQ6TS1tpTr1UfBzLPVhbEeHO2x2tZvMPiIuF4YqPt8xLhPlHn0azQubeSa+r8btBYa
4zyWSS0RjdvPWFRwp/kcFsKihp/lCVHJ0+0jUdH7nV22Y7uwbJLAig/Z6symbxfqAk0vJrtNE0me
t1c7k0jD+kqCgTsz7ToZC4NErMsjjrJRLCrRTtOonK5o703vEZkhxvOVVLp1c+rEXymbZH/+lXRz
1KPCorJTRSc7ykhy0A8phRb4YLQzjyZDr6ATW1w77YuQhfCunc7caIxYK5BMprr1CHW6xniK0u/j
MiFQfCEw30MTL4o4TeXnqH0fS1g7LK/FoyKLxRYrzrwVyGVeFzL6xD/u5lgeZzq2oxBhLonft39a
xcQWK8V0wn5p11S+sBv7iEsVE7nSVnu5vIwS4ogRWLyQESqFDrNTNpQCkI7jbNy3awKOLucZ6/uB
s+vEQZy7lhUqHDqn/m7un9eqF+Je4fSPaN+TIduQJr9CrlM+qPZrvVyVc9gM+8r6RdiyK9AqftOs
4xdJDu4UhElVDex1cVB9MpdKJM/afZ/eAPkX1o7sli26M9+v7lnKi5hquMhWzPng8mEyQlqq+4Wi
TdA6+HlQCOyBfRrxiaajRDjbI07Cxprbu9HvEI6aWdXB4U+ygW+mmWzCz65jT+9GqaRT/HFhIcE5
nUBfcvj9ZyVOTG4f2LEnBlq5nRuO4SwWdp9JWBEM8N2pPiY9jhsFA/UdTxAUgNnJVrRxuW+xcssX
oGLkZl3238G7UHHYcyeXe1BwcR5Doo7tVjTVNl6iWgkmC0YSdUI1TpiPSmMQN3pVU9He6pcD6U+Q
AkllQnv3Nuj1ZffhXNJHJeuCzyB4KJNmHIFwuoAV0N0ZEqSqlQzYNxhwcx2W8JlogIPb4PEK97zA
oehg733niIy7UNjywHklw7Hsq5n9g4nU7t3OfeaULYFD3/NfGUP07R9unRT9AbGafe1Heq/F8F7z
8wPOLv6ihlq4vT5dUqp9i8GuLJb39lFSNgcCpy5vz7eshpuqTxq5sefX7VtD3XsALhmtTcCNZUmU
u/qqXWSj1tI6pUKMkdyQiSIrK0A2Al3sIJCg4RezGSkJ0CNwFB/aNclM3zUi4Hecx1zvlLSUsgUA
rIp8ZbgT7yscLQOl8CsxQpn6DiD5LVPHF8s39fiPVA51JLbTsTBDQ3k8WvRxvI9rZALBVvMX7pC0
r7Ng6xdSRUZnVwoy/qRNW2HDfpP0yIhdvJKoUDF7nlbBfDMNzWDGE97J1bErCUa7QhS63vkZxzBn
Peo3pf7sswF6lLhSROWMWqTqAqYs3MhcU8mf85SnzkPl2mjjU+7h8+0VGGQU++Je4pts43T5xH6x
EWSXjfMdiSQRiJIl8CUZ7OeI7BnvgQ6wEgSCDMExY2jzCoxAy+Ydkp5WrkEUJmXe5etmSXJKLfCl
+uJgVG4DC/B6ZzZkwJ+fK2/YThEVHAqOtzTo3BAozbEEeOti4aXiptWNpmVJ+dsaKtRVGoqcsR8m
UiUwoniNV7YN4CF72glL7KnbWRyh2YngEIii0yhoh1qxFi8oABUcSMkfYX1YtFGJFnB+iPXMyhkw
aZtraDolZbRPvPrIlO4GndevvX6mxOzBloqt1060+fPXrOm92lxJHonghTZHG40hwPWYUL0xHvRb
FSSni69P11Fdi1YLstx8tWzQ1QAl/0RQZg72uhrSJgrCgZw14hBtzronc4XiiDz0KG7UngN0EcFN
grO87Q+eZ2M9rl+kbcEEbBn/B8SGyr62jcurqh3xkeeq58/PFewzmpMUwI8GS2krKP1fbY+Jft33
aJiu51gbkaN+E3A+cyXRl7GTxWCzxTne1kv0GSZJhcBkFEZEyiaWDsR5v6APXmuljo1DaGiqdUMu
/jVGVrQ6nnvA5tUXuMdm7gh3vWWjotSJjqMLLtiaS1otcbKkJ8YfUuwIzC4cwqK8yFmDlqww36g+
dKOLTJOpWiP2KtO5qlw8op5BkfQirliS6Ah1kW3Ftej+ZpzNUMADYWwbwCWQAt9FzaL06ak8UPVn
Qs6qTX1LKlMdLOHLry/Fhnf4AFVqAzktHOoNAFGr9eyMSRqcRXcUuXlkYYvSEJFYJUKlBHf1CeX4
UnXgeF4Po/59b5c9IzhL0dRpn/5QADOFvi6d18yPAbeKHrGfdNgu6qO5Ofckm4ou/RCn/73jq7P4
oO75A0Ebs964IjAWdW3V8Uoi+d23wPhiR0cFDs6Iov+YTKlPPq6wph2eFc2tS/Ubo/vC5ikJqCbv
9Zqru+OOAp5qJ2d6EC/cq9Lnyc3knra1OevMS5aw2DzYZOyyuSzGfRLyj+w+a2sqFvwMDCq0UrF9
08IR9tjYgIhj6C+hzRx1MLMUuJmZ1VwQ2EfA4bWbjhl6KXLcrzhxwzK7aJG9LDjrQGzqyudSpJDC
rERWkBcDPzzDAmqB3ee4W4VoeoOob0vhD/rD8Rw/yg3+RywqOrYObRbN2H3JUSzFoq5SF5wIraro
m+lgQWUV2cNhqS10vrXNx7v3ZPuRfD53FbpByAF/hIl5rMtPVwhCU9/PlTLnphru1nrsQmYDd42N
/mngw2FXS4HRZxfyS6PiHWM48DuSsaFjF9mPPb+RTQv9was8ce18b/bUbAbYZer2zdniEOPZmP5L
y6SV8wJui51827/XVqfIwp1YC6V9IYs/SIk7/nfehNKC/fRXq6gFE5fLcjhpPVIrQ0Uc4iyvFe61
jqCz67+zkmuS8k6qsVOc8fgRInW8QbcfinMwAtz/4Q4mTdfzKw1DEiPpUl3tfKU/CwUdTYrnJQ7l
I0pD0Uq+4gwUS3viFhXzCvdZufWrlLlJjfjc8KpCxef37cbBzYR72l9bYvo+2141Pb7wbpa+jwgg
LIw3d0JKkbYTpuJIG51TLe/awRgaBNCEVl28X3b9D77tEPTM44CFTaXg0sNKkxBTDzwOojG+ya3w
KTKmOX/48CBKz5kw3BoUKJHyyCc/m1gNPz+Pm/AYpciBIhMFGxb8tWQRsIHoK+ac3EN+oCZdsLQk
leOeuSxXEfqHgeG/X0OKPumksz2Ab/7j5A/KE60cwvQuMidnLHRyNHnaO2fHihLR4nuKIKwuenIv
NnXyZWaUwn99R0gJUuLk6Qc/sk38me+eIjmdbhBXiae5YL2UnwmpGmMZkKo0oHrFSaXyDP2KI3Hi
Pq8uukFrwT0pLdmzBzk67aWziIl2mYCkrZZxttX3+WNJgZ7J2tzq0jDWy4N+RlcXYloe500wn5jk
myyqfj9cMY+zRvadA7lehBmFtFQ6Xh0/KmmzNdm9zvSauaHoquPB0jN7Eh/VUQYnnHnhpWY0qW/B
PHquwNqOEI6QU4gApaPiLX/zX80u/4+M2eVWF19RbTlp9/qK4JqRC7Tx7jAa/8KIeAQALkWisgm9
Yi65gogZEHF0KVmIFk7QKeVdwdXcLTCkCVBdXocoDEQ9GU2qHpzsNf3JCUbWZIsb1FxARZlwi6hY
CML1haigj9mRqj1K1fvXzhhujgvxjXtrQxSrMfc1rwwR7mbzdhS/dLnx/TIeP1OQldAkoi6mNiWJ
xsD30S8iFvrY5S898f7cK7TzZmlEtkvBvzgnoOt4XRXYFe+WY6Jw1vNer3nwe/mT7aJ/vPldQl0w
9zoFxRVJnzgaBMPQKTuevyUZXr/tQrxvZxL4GoOJJ0cFFzF4qn9aIQuO/ClnO0yCoUm3fYn/Fuz1
P2Hfr2beTKPsUazzTgMbn8cylGJmZWVMOHLR6SeqvWB5E7gK7GyDXZfESV9Wd2Vmunk+Z04yv2ZU
MhfsiAIUhwgsz4tBHk29vi0Vqa8xwpcy2EJLQYVKkNGZM+3kJRgihotV6KWtRxHzS6FL5UvTOkXk
Wx3IIgNijxxGfs0lC/6vlpl4hEePA2GUT4I0QAp8iycbSwDq7XcDHD3vWkTJ1FWBFIGIt2eU05xk
nJlPbh3IHqmh5lQ1B/quZDr1uHUfQKe0bKF6k1wGprN4uZBJdCganu6fyR+iHCY9Y+Zn+3riozP5
PqneMBQXvuHTPnt0RT1aVimo53PCDcJ3nHEbsFLXSUV5w36TMicotcnty2RgiZwjMNIULLPYfEWT
4NDmJHpQRJrrXVtT4TfE+yHrCiEy3kvruL9C1oUWZ+VSGw3yeiFsf6ZtJ8mnDhhgHJuLHFwFytRZ
RYbmHrT/vRhVbs3Li7Tmu34LGBww+1atarLMGmgI55cYt08nS8QRfi+wStc8Ceik4J1BuVVYKtQO
a9+LPQy/vMAD3cuAhR2cKHOEWRP3MkZtth1GschSdA6qWOdWmcWQOoSvHUhhXJDRL50zi+uHRWb6
F4/KK1mzQMf+oTd0nF7wIkU6MJrJ2LAc/uypJhPlFRFFM1HMLPtw9C4+fGnQ3cHAHNhSXznwSawb
uqIIl+4OTPl+Nofr5hbRwPslH8UWeqnvsq966KFarmv+N9cTTVgF+26o1jtsQ467tX797Eb1Wt32
vNaMFAvTboSMuMT7KO3JRHF/gzuhjdP/M38mnskylij5eMEYi1gq24Hj5P0xFvIx7vbe+Ixgua1i
Pl9vvekP37XCrvaebbD3uKMavK6lAX6lLfH0fKosLHHdXoPZ0yWV0krN425iQxlwds3r3CyWwo3H
CiE1ai8cU5DfN3fSv/eKiuPiD6HTV/6NBvrJzlqg1c9foF9nqx+p+e9Q/GBfhBxRBmz0ZN5PmF54
3C3Q2J+xXZag7loamUxWQW1nhos84llguAG49XftvrsxMfVzgg7QSYZkEg8oSFLVl1iCPxSvYJDz
oiVgMcNDFb1uv8gUEd4rB8G0Z8JL9dbeQ26Fqv+OsPXIqbQSh4GnEST0J7CrqfGlUB1xPlc5LldG
yqrkhJfLmnuN2F0KQ5mPZYp2JEWLI1oKe9LXDhpqAfLoQmVxvUjY2irA89oKL52uUJ6Vrot83cCq
uljU1vzZ+cMQTKT+kr3VMkDB1QT9shefEdwqghDL3ejqbkoLbk1aDDueh5B8+Xd68lqcMQeq59fP
DVNSvOaI/5DMWfTt+JLBRwTSYDgE7DhR7ma0+A7RE8AN1elymKE+XwGBgbOXRnoxxCRKARXmnk5/
Bb/hylEeZfbOIFWysSHi+Mvt80iZsTvXzdsLqevbHTUnF6gXAHO78ZZQ/xPrPU3aajLMa+AgiQ8U
DShutnHMYGIH/EafNJ7C2A37GSsFD3HzJGfVHepo21/HcKIO2zcViydLLcV9IlslVx0gepQkNU5a
4fEfpZANZt78aqR9IfFWY8rENUvlK1pmLTAnX2gWACENAEWxAxLAhuVM5JfVT+mpMTGL3ToZ+KzB
XH2wpFxD0qyDgJCmaF+JNsvO4i5lC1n5BpGKEURgeGj/V69ITXKDTAXNiw6++E0pzeejSb65ApXa
RyBfbSpt2p4MGXH123w6PHuWq5gCgtJstE3YhUbynPbAWJApz94Y3CUHJdmfIDhxvPP5U41SRYd5
puXPDQNM2jlwKJR/UPo70X/eBIcjNmvN/jsBgiXK21fmu4bPQosOj7Vqpd1BQKeV7deUS9Q56TKW
h15tB4msYhPmvgKCxoAF3GL5Ebq3lcX+U8wBwlNcmMBoZ2Cz5oj+yVm56/24IqvEdqnmSjLmoI9Z
qE2WUN4EyDLWpZRgbMRjomt4tdfZcg+gy1a4ba4Cb7bv6XKFZs41y0Yy4pRMHQt+FRLspt6Vivk8
THnyyWHO7okKhl3F5FnbAv0+UDg67ubGWDllB1QqkO5z4MgUJXhMdpIVgRvFlGWR/x6du2f3w2rX
9Gpi+MyniR3Wop55y/+j7cLWSa3mTUtPRiDRcB4Iw186SXePREbLi5VQaGwfrmg0Aw5ii2hyEiId
HBs6Ax05Tq0q8NBexb0C+/X0ICo0d/8ECoMW/1/3N3Ovzq9nNRdRZKMyVSZR2OsovL/GgxOGmBiQ
cF1MLpu2yVL0Wc5bIfJYgnQ9aZ/zr7OWm1eU0e9nGOEARl6OUwg94J69A5a956BYI+fO5Mf7ZSSR
6uUCMTRHd13r+wAOYn9itDhE+p4ftCFXkSnpwSIfah47yRZtG+ij1d+kSZyRGOGTMICsuUyIA8f4
Mi7rsJvc0/cmo3vh7FW727eMbANZh9vINW7wgyZaG1LAQeeVob7r0nsI4I/6xReq7qwGFtVAyTXp
VYv9uc538uenMtCriIkxRJ3c9N6LgoUa8G9eLKrSxgtF9v1K+o8b142TTVdCl2iKC/0vdsBJm1Yf
+Dzl5cbDIqdw8eCmeoSd3CjJEEfQJZ8/gF//2Kqv3ZZg+5yfMAeG2GeP2enAF4i17BA9wDt2iOfF
sAxhXbCF5+9U1fFsa5wv3jYk7yxqYzNL/dqykUPJbjnUd7YSHCJGqVRF7HrdFOo1qqqRD2YRFGsK
quUlSA1AmX7wLrKCMmKTnSmeEmI1mshZknoWhFrpvDrbbnebOH/QUA0ycikGIRKbYCKaVRGA49jC
aSogoQXDyxaQhf8dYTkpdjsnuwoOu3xsmNP0J9EEN1lh0Pt+OfQuYEB0w46yqzHU2xNd4bpSuTdh
Gg3gSL+CjoVZB2UB+l5rcePE78/v9NkW1WkNI1Yu/lTjfjmw+sp17QeYNnQIkOpGm8E9p3AmJIA7
drTiMN/MP9sL30uBSJLjWiENMUTb8KJf33I4Wb7NecExtt40K82dnhGGjNxmKzLnOAzxLIGvAzL1
Xnj2XoZbwKOMQJEfC69CqyoEO2We60Od9W0qrtGS107BcaFNXr2Ql3dZTXpZCpuYVcZou4RaNHnH
aGGIxv4l7cTaThoOPlWU5aF3MuAy9nvQqFi4m0TdisyOKAn4RDNrlKt/VzznvrSOTLNbhLi8mCG+
dhn6xeeQYHmZyLwaBBVCrknNPqERu1rTH8BFkOf8qBXF5zAnANGkXS7mtjmmVtZn1I88TJ8lwnNe
rbz+N9Axb22qYRJf34eZmFNZZp5Duy8cMzXAp869VknLVuy76Uoy0jF7k6ut5xyDNtjT5R3YGyr0
BeDu+4yWk+q0vkcRBVtMMLIERJZJXj5hkHEQ7qqtWdXhxMgXlGlPY71OPLTrIkfUTmNa8DHS46oh
gGcE+5RbZtvacu6/ZVgWEp5w7lCbiEUyGS05N+z+36MdGiErE6KqUgPjs5bShLSAoCWaIMV3LxHx
4Ii8J5SA+SpYKV5oMetW8txRssrVZHQJzOhJffKkNLqB+r2n8/jgwJjAp6q+7hrMZDGbW9Bod2LV
ZVZPzW82XIopuNSOVbY/fahkWFxjEMdDpfppJkn6vjLrIVdRlfHyMVzJXihZZFa/qJPckc5D6TQb
kI/oAAGir8GxcMYeEjGiGqDNNJBWtHd7lJHM0iqN/tCfxQHZQDjBScT+vzmLS1nd4QzgXC8Lfhuj
e35Wpii9aOUejrKSMcUhwKwrpH2cYku24UmtX5SWBiXYGzQ6U6An/sBy0H+7oSax5cFPs306Fg4f
Rb0V9Op8ekZ2tP1zlxoGzlHG/+u7hHF+Sy4h2e11FxIY51BbgplsnDoBMDs08VA7UFgJxSlqq5Mo
NC7oDrKevb6XL90eZWOt0AMsRkQkrHvUvig2V2R1+DNpGvEyCfbB9DLt8czL6eV5fDWrC2ElDHGN
Xvc5sEvFqYFs6o8iMOk7aiZRyqwSjyoDPUmQBEQw10A/DnAvyUmb3wDkchOJv1Ry+y9+LvqqkUzg
0x1VumzxlV+XKtN5oX4GpJUlp4hXsbYwFZP5SQTaPFP871Jsrr1pwFYxPagix/poGMbzkxAwCJM4
VQ+QJ5mDCi9PHb71HyHDNqCqMQf0lX7Qc5xDU6u35xsmjXAn2FdXJZYikR+xEqISjchvC8rxN56b
9cQyf+Qs1RE7iXDWNqX+Y4yhZvDEjDE1Zhzmfs2ORBgzwgU3eHyxEuRdFAq0ZgIxXENG8LeFiGY4
0u/UuTeruiPVLG71IZcvTGUvv8AvMxPBP7pADxVZMfiRtwQxJ6Znrw8a1tFVWFjfO4z0frGfMsui
SvbBpfx71L0EKJpd4zKHgz/vHR9pOibH+ZceUdc9P51n04jYujQeIgLPulD9PntLiHvPOhTjizea
Eiy/OUp0mnitAPLkLwbQTecLY0f16bqM/B3yyOYzb6/Xx7u1EvTlVIqqH9P//MoB0I1EbD/nD/gr
cJfPyPiu0F/vG48E5grbixDK+fmhspXIa1rea9SgwOP9svvdk8yZ/5YRx46zwKQ54fSzgpm78PDh
mYZRTguQNn92g0UJ6NvGbhZmkmOfib5dA5Cj7HlakzopMDyE0aOgzBhCqduWUJhEfizV9q6iS+sc
yV9ceXz148FPk4W13dBPcIEOsBC6fthTxpoAx7jLdkUvVIb+AELjq/jP4If+/NvBqVPcM3ZT1tjL
JuXwG9Ko+LrPiGvNzR2nFK5gwN3wNqXmH/Lz552vWbRF+AzLRzyk5iFQbpcwjIZJ5aY81afKjIHM
0q1aapG0gVQ+gJINj4VXsKEwGxl9LzwUD0ofEVcEy5roZH0BRF/bFoFZzgYbzd3M5SZ/H8cb/kbT
3XdOyjGixU4wfArHZf0ULIGiiz7exII1Gjhs5FAtY16YZWKNj7aVf9PJ6tP5R5XS6ex2QjGRuJmA
SdlvaO/JJk/45a4j/rZV/5lmrSmprKEUjZ87tBRiC5gvwmwrkNzETTmQ1xBJWKFdxE4SGiRy4nBk
j8lHoVaP415wIn6GPCYZQktozpFx7GtRkx0Jyx48+BWdpU9MwnhmOLyyXQUXKEZdHF3q8dA+pWqW
f68dd8KLBELcRHL7eEYllFgv5XEK74YT0UptRaH5tLGnKhGI6j3A8EsfkwuEwRBlAGOAbsjKNSrL
j/oPT7sFpRLwMQtECK58FYCNCPo23I4l4Dekb209vxFq408jQK8FfxNIHxWJV9QcbL96bkPEnPXB
j2rGSkt7JJoQ9amDb1ZXD2e4uoFLLX6mRj/SuqA/uEys8Td4r8VCivVGnQx+9QmwWGMkgP0u06RH
EXH0Yw+NZJAaLu3jJs6IJqleVWvQOaImaZGeIweYoiumiPgj7fE7AjsZDVRSOaYp29jrvp3Bsg5/
0JJUFWT6A4ElcwzyQfrVOFKPNhsHyTgwRcWRTUmcZtuwSBtYcLJyJ3M2hDe/ksTtwDNvvK73gGL2
0uy97D243lrcZmAk0irmEtWI+yPfYzWLNd8P5XO+WD/U5XCZxB12EqOjYOT4VmVgFUvJiqXq7yl4
JkReNO3vobJWBCQKdSHdXsnLuNVR48S/Hehy/V03DQAcJr7mTCnKV7MxTNao8pbSQHZtHc4Sag/g
rydkURpUbqM5vxPoGHl2NTHdWmBZFhuH6XBi4ZLUiGtZcQ+j937DBx8V7a9y0PeBkuzlu9pbuYOS
nhByfKlDI7ulyOUitZqMQtn2kDWUd1k7ytXXBZ2gfrs4NbkjNN7jeT3tSrfoOshhGEfIWnAio0OG
1ChKDYjf1j0NO6zRE3QCzcIMdxi3ysgDVeaCA8nW48nj/vxRl4FgxBJ/CQF+5caQswv6oOZX6lbL
HyEZKKMDeAzJkT9B+xVqWfAXPQtBapIBFVTaukjxicD6Cc1yol3ThW2qbRP7tgDp+1VOVQuMzB+j
pN92Wj2+41GNUBXT1fC2aAOxltnxSLWd6ot9wX+dhO/vZKScs0Gysx/brSMRR1N8YaEBqLC8pc0W
6CK7+y+1XUCXR9vK3j8V506anz+aocH1S7JXQ2OmkX/Gxcttki/VfVtjkDs+iFNiwYHD3mVeKbri
4NGS4YGJI/kHKl/rlsIOHIG3KfIc/+F5xFgdgc7/Im7LyE6HDKQeWslWpXh/kjDvPZ23SII7/OFe
/OUylx4qW3fHGeMWlWqSPM3ejjd4Cea3HH8ath/+mcCGwMy/LWXrq7G1TkcTMSAzFqUhzFMYJOiy
LGFE9OfpH7BXHhpwOIbfJvnsWojgCoqBAThypJJKBjs5aRoH8gkc+Vw97es7xMEBY0aJOP3fsuVM
iIW1ALgwkUVrvNIQqfJJg+c0Wqp8V17j+Lko6tPeBw47Yk3j5xyHyWYeNXjhjj37Oatx4B8b5ZNd
WLWhMWVyJCdGUvar9FtSfg7/PkjwCAEE2d1nPhMWc28Z/1NOhjouBLxWDMfQtlIkxd3Ppvs+/hDp
ttSnjkoRYnaBiUhgjJRxndzkJHjAESMcVpkyOd5Pvhp3PwyErxWM3MlNZNowoxh/ZrDMK7pltI0U
K10Xdq/W9E5TNFr9JG62yE6249n8sdx76wOvZPUFuYhd4OZOZvUl2AJj1Ifk+JP9xCYkLTa5QwRv
i1AoEExm63WZsMAnXBwKVnbi/H7Yj1yY2xrIV7SNzuAtzBz2sbv+hLOs2crTpf+boLaOj2eeNItk
5mdTZaLlQc1V7a7xCG/8tI0bIPMpcPWoDcD8TXR8dUDWlJ/RuO5jrf8o7KAEal1qLjJu2MCIBj2G
i3kAB6zXK/L5QvQ82dZ/Oruc0+pplpRdPYpwDiM1Lxovp4Hy+wRLLv2iE+VXMpLnKyF7yAXNT49v
rYJrdC2ivM0RxfY2cKCbYOWMEkp8cpFdQmZQqLIwWTsMC8Ek69V5z8OL2zSdj+8NnRlcbZCChy2E
dJ5GRTq7Pu6aOnUlyaeomkR4HzBUcYnEgVVXT+/1Tbzb9LkhBo1sKywHBmbUnj/dVCTf6RIR3KCI
7ar3pbj3QOJYYUf+EKlP4DD2ipZPAXEOYwMlQaMcCVgqb9NhcttKPO48oPk63IONG1egj6xVV8U8
0hMy0l+ZAOvxPuvTqbsRMa0Wrcdu4ibwfDKHRbkz87DKFfhY+9CJmScqH6u8zr6+SvinZnaYgtxA
ctgb0A+qHjp0D3f0H4g8FJzv6Cqp+7EbOvqK3oxQbq5J9cjhWihll1gh3FsNarcfrvcjy0bzL6C7
g9Gr1MapcRs/asyVAPBnPZz06njdcFJ26ngcLnhQyVYWEOa4+vdWjpSmZ9kCA63O2TgrmYFKZc5C
4X2XJqTU29/C4oqRdmpctIQZ+GC9nryGsR+vqJ9ouB/OJhP7VXRxmgflCxS4F3xaFdISBN6gyiCw
kK9pfgQe0ywo9fuBdr3KrifM9/bCvzWNdYucH+hw8qRBBFB1PTWJV0YFD+Uc8Yd5nw+wZ/RDkzpU
A1bn+0yMrkl5jjN1xhgdKFmxoEIL2SJS9MaJyJQea3+vib1psWl+dKXD8+PA1HpG+Wxjj2qWbuOo
zFEbiZcDa8p6aeHgVemx6C1yA63jP/Fo14GMVa2kKjBIbis9zvTJcXc/dag8ZzU114ZfcV2sMP9+
hHwTvJmoSbwQFIKOexV2g7ok2vewFQeCW/vZ0hi78BEx2mZ0bhK0A8nFihKTvbbKKSR4QdgmXYoX
16gIhSwDE5yP53zhzZ1Di+exOpVwWHBwptI6SF48u6TL7Iii0cyFSiOIJmTeNsKaYfyPmhjdqXcE
q9+jvOWCR4ejZdbaEU63bdhbjZcmAuRfpTpcxFX/SJsxz/GrRTx2nYnxfafnYhc5/mRW/8TQTzgA
LevbdhGuZhLpYaJ8p0Ljj05TC1nEh6jKlN+eBhBJz0VOxec0cWoOYQy2EBZJJwx0UKjTB/JQUvxj
agnyESQn8WRN/Oqx7VigqzSymjK6DXtMoF3QoqdPUmHaiuwWCtTUgFGG/izemwjSRXPOESFP/la/
gcs4UqAJN3/5k4HnYLUkF5MSlY+ezvxCnFbPze4gknYqOO+T29aHBEdWZJp30p4p+qI7hCGHOlUo
zx4Os+TB9AGCEP+DWE5TbaOZfeuVMLOBSq1HBRKqK9MYizm3ZpeBbm0o8yiXOE/CFAYjvpoAXESe
3YzX8igq5WvO3JRLw0X6jacs7Tm+9Wbl8pJu82eID/HSLvDduHesOKcr+5IOb+0KpozZwMNoPOf6
6LD649NuaR8t973maHX7IPi73/OHmPX0h2fj/tzUm0A6SfVNPKmW91cpqH6C3OMGOQ9qoXJUOkE3
Wq/vs9nueL7LiItBsSkVD+hfmPoorO0ojlHOEdd2aH8LoL8dwh9WmGXDhO5/Vau6WylwAQmwnZWw
clzsgGnrM+quHYT8ng8cSssx0OfqxnXLjHUwEccy+Y8oV5tiZmIoqRPOY8VsGvW4cAAPGDcwLGND
S7h/Ho/JpEGuaIrBRGk4x/ovjDo/ICAbYNLWqChvIZQgxCjgLXzGqOBYCHPVTGt55MnFT/Dir7zz
w7lkwjwn0EJtkIhWUj2KO5crp05cTbfhDzmtD7D2z8uW6fqOjRTVAqYaVXcvEHHIBb7lOY0lj5kM
TIKEOQcX6+PAFvK399lQU5sazzXDcmfa/4zD3qCfK5dJLE2y32akiWQpR3TZCm7hFu7BhgGdUmWp
fgyBFnVYJaUsBv6OyBWB11rShsdJx38EQkIvqU0CCcvyBvO6bJEqnDZjjxn62KAGOmPyEM6k7E+b
Tyo90rgiYODgUKcvUgT6dLv5mF826OycNYREx4LirMeiL020UWa0h5XINwQJRzR9yJ7uPULs78Xi
voVXmKdnXvosIM85JfZu/QX0EpguZaMgSNmB5ttaUTjada7WGVXMB2ILcNdkSO69D/u+hdu52Z41
29biDulopsGql9UorwP0EE6f1NgMOwyoWXVyherh77xY2GPauuNYlg+GNKgOBmDgWMdKOCnQqmt2
eOG7UeHRghKnmQuzCWvWWl/Ma4CyMrbfacTpa5eHGRV1znbinY5PfelfRnqfYFgLUe3Sf4UkWaUZ
/K47ZvKpy7GuxlszWtgtaMp2OU5RJsYUc6jH2eanbCzuDF1Ymy6NQwp2wZ4L7P+hJwSvVRWZU9Ru
2tGLeRjgTixOWmGOsqiOA8WV+isW/1WyqvN5Rl6WPQ9LzLGIDPLiinuZ/n7UCKcZjHEBALqm3qzf
Z/lRKMCLpjhWFrHUmhE11EAzVo/W5KDk0siKQyPXFqMGI8HWVB9ZpEL66tGu6kWzRo5+uUJEgdeB
COkKWqr/Jm5XdXtqGPg33eCFyoJOo+IdCHB/7Ets9jcqjKpNHpaJ8vsk7tz9ofvUQMTmO6Bf6AvH
CIuEadNDR3xmeUp32fZxdnfSO1at3kNERfqsDsAlz+AALSkNVGno2+2XpVoHSeW04VJ03LXDsEpB
VS9qN+QfhSM7zrFjibt8V0Aj0r6GHGANWnKblvRU3labvdN0wwN3Wyaa/cWRfSdgMe/s9rzNIOU1
txwNrEShQXGz879Xg7Q50/raab5XTgSLbOwz5tYqxa4b1yXWuOeE2evvbDhRbljKeIMevMDvBWVu
7w0yo9mUopQazPFcOXzCIeKpywSFVVHZ94SxRu+uZdeq1lQ4Y7sZ9PIeC3Pn5hpsG98FuiLBSlA+
DvY/woX9phd1bgm9Wj34/aqjGU+duBa6oLuMecP0tcHKOGwcK2FCC7bdwndfdLY1Sn+vxk4Yc2Yv
Qyby+HJiFePhXokNb8Vv0XjyyLnEQ/CkvFTDiHgthrKpOf5XNb1DaH1lz8n00VKvkNK9rGKt6Kmi
CZXphSY5GpA8aTeVrf1CR7m7drWbRHclXzoqZ5+hVYioQ7vVcev/4bj/5yju8QIakN+sDxRYOrVv
etNsKr/6eBxLw1eIQyA+XNrkRAf4zgmNf6mPQNbxeDv/Kyy3sq3+KSdRQWsSXFVlKdsREw+0ALl2
CJHFy4wdnQLlXU9nhxGY9MCk7ylzJ3z7UjiyKC0veiOPzHAviIJTJrlSOfZUxxxUZ95fQzqUV8VL
/OMqBmKOEFuPpjVNL15gIb7zOH5v25BGW6bK3xzuxYt149oE2JVRwmuuzkblkLAILqK/3skX/8xY
bII7+n8jxnN+wSeac0p1XtqeEOWcn6AWpoutz3GkTuRaf/G+GrN2nySwQ8umyvqV3MnXUO+RePZN
Y9ifD5c6wduHCglUHGCcvmdU7SoaF7lkq5VBA7rGP7tkpAAcnt7wDLvugJLV9ZHfxpb2nLlphD6u
ID2Ov/x5lKHSdQYISwD2dTDu43rL6Aoc1sv10W3khvmIUZzgO/21LCruvrjDYN+v40ZfXNmSxVWs
aPbZndA1XMM3yzjGAtpBSmlxHTyDt9TYyhJlvC66FgzRmxg9Oj4D1bX/Wjr6tCqRmaDgObGFh3cD
tAio2yBuKuk78nVQkWyRTxe2cjuv6BsXam1Aq7m4/perC/qfDlPERUrN8dGF4kuP2xOj/K0f7j6I
mime2K3sAFClwlU9sJmKbtzGAKPHecseS27guy5GiseWW38I9CwBd5TB0hh+8FRpNFlje4KIbuio
gCoVh+/zrDf8lYPpmqxQILTC8xjXt+vMpuZ0avJBpZAUFeFzYfbP6DzSpFL7TqaywQdZXvi3mvnG
IIJE3lm4dMuT0fd0FBEMWUqLfOC21U5eaCs9tOXfsATMAmReZR5Xjo7QPt9t2VJuv1nbFBvpzgv5
5yVzsWUwZMknLdjQsYAtk3i5v9ugFWgL6IZ6DPyJ26+lllDmglGYypGD8PpPdnQKH+a0QW31ubE/
AXqJS4baScYXeq4nfcvWkxMKbFzjClldCp+BuZpA87BFuIguOFbjmeAGB+AgBgEWvIgZcI+aT3Mi
kE8FCgeK1HywiP+YBzZDQogyanTb8VLNMLVy6imzHcQzLxdSmXBhokf5lRGsygALQctcX3cv6R1n
0VbPTk8WiPnKGFYlhWmXp5BLkAWrnv9gDA5iB1Ye7An933JGsC3s8QgfAW9OQnFiyfc2WrHT5NDh
rdrTCMqU8RnRygIIJ5QIE+YXW6Ico5YQOAdl8SqkRKXUQYm2LN99ez0yON0Uq0HV5krAay71138J
5txcmEw5FQ48UHygcKnBKrF3qA8jl8VCqYxvbmm9zC7cwDshG5YEDIfHBlXYFcjU2/SqUn1w4G8T
pZ5lbe6P8WShdndXiGSud8m/ZOFpK68AV7CP6QcBa4SunwcHOVb0m+gT1IcHrXB4YNRhTAyjzEJq
06FtOjEO8BxyVCq+OW7+6pb1tznuHt25ztZ3bzvjAW5B7qZ8H31OtV3/sRXiQ17n+TLXtRhXixBg
eLYxfptWAlWJ2nZPr+WrGUt+U8Xwl+wfRCZESnZ4wWqFa2RLNcTM+ItwWxKoxi2rYXrYpWtBqnS4
kVxj7EoKbsR8bjdpDZcJ393ks+tlD/1rqG8vUMScsWFLX9dBc4HR70ui7YwI0HVLwTWFoz0ytL54
J9dNvKJwh5tlfOOzPQWMyZ87pLc1xHfOCLaoHKueXs4hDaoEW35A9JAMSaoEzZ+WPZMNdreGJuCf
irCKRVXrzx1gsTkM+v16afBDDBy0aYV8uJNfDD1ZbIJ4PY7LoU4CGNuc1UIZBL5E1XDJ+bE8U1gg
NiDx3JUoSqTj/xuH5Ees9DP6tEa+J7SzuvHpyVznmNWqHlW238+SSrgXPznMjrzDXbigIQxhllzq
4LmDLjS/dpICr61wb5psbHKCaxvAKOcO32MrVRvH4mWXOVHw32DyZv1QRQu0q8mSpqrHqPF3I1/M
Rirt2opTO72vFFszigARSCEiFiOijNMBmdsL55mGLQjRAf0JVT74Fay34G4Ef76LWOo1IOMCQZll
M48WVfpDFMKnIbZosoPbDGzUfCbRyflRyf0YQYC/5CR6eksxaAjaM0URVQUcIubNyQ+rfhFfC8tQ
LQWS3nfqD8AWqepAQCoQJGlhDxrUnJveDlxuXArgXCb3Dxw7mMKzdvMcmE5gNIY3s2kMK7QR88Ld
0kEIuzXoEuOJopIommA+UwUaBZNHkve+CpOOc9rHcwaVbqRiLr+J03KMyb//GshPwMTbTEcaDRY4
aDVdEHLhBJAXwaizdqn5MvTegSgYJjuYOG5rUeO9CXpVuMvvTSDD0dxSYZbff13IK6QgiiqcmP3d
enq2m4r9A+rQVTlm0URnZ8HZbOh1QjydzG6EfDlkjlOuB95F8ISFsbBPNR3saHZKXjpWOrV7+n64
SL/+Tpj82Vz9CxuK4rn1erLEHPDSAo2DXytGNyR6ue1r8jAsyzm83pKaDETgvbgfI9pgXS3JlDim
Z9IJE6C816kK6itZ/U9IjxjXiZvmvlgHzozbSvvjRxwG7QwlggUa0HDPOL0m5dQTJtNGVg+Bo/Ub
aAZzOqH+1gN1g7eSaAfH5oFu4itoa/NPHqeLY/LvceDEeEwh5hRLKk3AH8lF7qjwR2/b9/ig2kEv
78fV7i2UfbivfFwODkopPMdOs0VRw8bfRznz9lfBkOb63Y+DZPwskRGk9t85Q3XeeSGmlpQO8BWj
eShmnRhRMMQSp2XJZKsrZCi/7A1+ddtJzxcCtMDHZMpWz6FgIUkfJCQ/fIefw0VH+qihun+PC8X5
RmEYYGh74d3OJJRo/zAe+wd7ZYxSRybo4X/4OfKd+Iq3m0s5xhwDvnjQOHvfZL2ssIRBYuuJ3V2m
08JDUN1aB/dseMckpkrj0f6KWeY0PDIvrGgSEajvk2G8srnIW8F+zoknkfhwanrC8ZmCp24bIahV
C02JpVCUwjBgw+s8wDC/pREIs0veBXNj9cm1SDLPHPAjC3/Soe39QvwMSB5TpMMHuYxzf4KdFE41
/x4vtBvqvhIumZJxxvYGX28EbwvnD5B1/4lofbqjaEqZ50a02wN9yJTsZ4wqUddC6G7i8c8HHDxm
EM3N3K3HZMIhsquYgsL3zxbiDY6tLVexDm3e+xmIzWnZhB/DqJ8vY2KeHztrjp/9FwDlb8B7xULY
cvb2ZsvOg/EZEs+gmPbmEWZSRL9qLn+k7IhDzgO9PFGAgErozLhtuVomO0qL8M2tUmG6XXV7+fjR
szbb13J00/4bYdnxuBMFaizw3n6hqM8zrcczX3RIHdl/DT5wglr6q48vehp4PvFKvIkn9GNZIz1v
tgPTnwRzbCuKq4+BS9vLF+DgCdJWXi5Qyfg621oTgH+M57JDgm8i/4oHe7nrbgYdBo3KA4+qe0nn
36cZOf8WyN9Lr2KhLm5CTbU0Udh3LRK0GSbnXBmGX5E23UkMZuztwPBBLmHkdJfZLudaYMxdSVGj
EloU1ohWzb6r3IDZ0tZ+TB5shMtdqzEBMAaBuSwZdJ155dWnn8LLj4lG3c5ovOBY9Y5zcq3qiFE8
qG0nPNiC47my8bczI3nbJKtJvnGm8ak7tsvr+ej022kmJSCAkItMmPKTHoZOUYAt61SHpuqQsMMF
+juo4MATKkfVIL0HpIrICR3qWE4DrEsZFeTIhcl2l6OgCQ2lBIPS4EUlK5rzLW/hdcaba6/j4MB2
2s7qNeadmuU0uL6PO5PVsd2ZBRvIFwulj1r/B8OlCujsHgBdrpk18G/oip/yX5hB84507FtgVaUQ
6dixPb1U1gd9C5OEpnj3/YC1OIZdranWz2SpnSDgnXMdqh6xnGhficPQPrKkSY+6C7jRja1BjGc4
WFSaqjPEZsX4ho9ETX+aP8wj2/MJZxMVUBdLxZARVJ+VU3g4tWfWAK+Q80SyJ//NeBB3SxEpz7HX
GdOBwjPcZefkXQEaBSuPOIH4Y1qw/qn6MfAJ/R5khlsGC6GIq8pf9gFgvpZ0aiPrq6qQd0yPU+J/
9E6nsNQOkfFTCCh899vTJWayxmlIBGz0wTOYZ8YmA5ceps87VA1ywCqJ0XO03AN/YqEBLWwJNCiB
Fz1P7VbllNNhq/XvZUPEQXOABw43v1js/d+Ey+AzbJCPw4OqqBLvoPl+7pBmiM1Njkcg/BRFh2Cg
EQS/uDP17V0BXDI/rgh7JLqu19UFMHEbyyEqjutkNafGxFUzfHzB4tyAX7s01po1JldOUcqZ9cOd
f7vTExH2VzzjKiLsTpC2H2un+U0lEnUdF4X2+G5PkLrkOZ/x4ogxrR7t0qkjxUcsfM3WcRTLph/L
BYgILbut/99KoMrvXJgr5J1iwWbQEq6qi/yH12ycTdancSYUdrEr0uQ245AO8H3Sjsv1nEDvPW4M
d5cYKDFUYnzZh7YSIunp9RTdo1zjdoYJ+rbSt8KKh9Fwd2q+h4iAktZ0oPRfplj66aGxhg0Jnd7e
w8SmhMVEJ73wfqvdJvPJ7bgI1Ix46OeThLeZFxZ7RbRv8LI1bg+m+QCvyYf8rJrTsAp4QIJfb6lO
DVaBYmoMP06jRPcHB4l6ey1zNDHo00UgvlvQ2ATuoXMhduZDVQUwHADdgCTaub+pxDwwOlEAD4dX
+tLA62HZPFuRJBGqySHID6SweJ+1Hd0sFo1bwuXqlYD3ly5T+tkV3PCcKCqFifaLqz0JBmhv8YXt
1kQqdnmz6WrXiuuFbQkiKev0KT70RIzschFQvXwqKD7yO3oSGJz9Q2vbg/FMPkDAHFWFMF02FR2I
VwhnqCF0zlF2esqUHWXgeOUYJeKUm08odnCpEJDT5FdqYTvjJ6d9seAhO9mNd8Zh547hUh3a2zan
EDh6vGjz0lKrFtW4pR4ldHLMwzxSKvc4kYvPFiuyK+e87M+g2axnsV0LtKEx/SvA8z3NWoAfzlGy
djOK8IUsCxN9lotCuujbDmYzOTF5KBeLmSF6QY+aoFAgA1LoHaL0JkLQiBjpa3n2xeZFSu+/PyAJ
MD9s3FilsPPeU+lYEAsVoPGeectfJh6aYudjzs96DuJ+uzEzGcE3B2CMZ1/Ql7p0aTNN1F71Z8Xm
D9j7hT08fDOdDrC9HR0eS0YIBPCyWSB+ZuhCfXvo3cD+DywVJL8buR55EDbsJ8W4Ufb5L3ng4Y80
8euZEsyTeiQdEBDxYgXv++Rm2ctZ/+FtA1PxZ0xO5aaSn+jpuFhTWRxu545GO+DoY0momMOVRtvh
NEJFGxEIRHwhNc6r3gmKtBhfMTEUsebQN84lx3I9a7jOvJyBX13ncAjq1qbeMasO/TAZXlzVR3Ow
qQE0FofVJg1ANeeqdso+0pCTvYwOzSvz5GJepARUjcJeJ4ztpyhOcNg7HTD5n0M4z0ke4Akz1A7H
uq24J8ER+v7+YMIXNXnoSGLfwb+Ks9WRaceSWrXUSjU88tG/pKlDvVkaBz+PGfU3YUnQPDIGIvxv
pLj3GGox6FHuqSVmkXyYdfiWgVNCw46Xk2VK+0lEZ3As5NF1cu4O0EFHINxLK+9+XY3GjCz+baXT
PSrN3I0GaO1HpW6cXS1W8qKZK8inhGBT9D+Ge7M/d8S3klPfGAzNG0PI9UblxQH8bgEAcbG9Bo1k
IF3Y0d/B7iFC+6bR33gcQdeSx5e3doOuNZ62xrkgxhK//642v7YT5tpCPabX916v5m651o3JLIL8
8DImououI68pXYyuUKJyGNLg3ESVeqTRRSzyRkAHsMiTnjv0fp+y21mUupvv2aD0Vd+1Kyo56aJf
ekxPNPo0bjIu/Oq2wQoE5Xk+B2lTEmZm9b3o4LzE7HbDN5KlFJsK+hCE94qgV4VpX84Iq7TFeBE3
s3dNXQWEB0Giu22jCLdRpu9up4vYnRSes8y26Wdm3kEVIJ13hGX5A8ojlqLZJxCEORP/m7PnE6xg
kz7wT8z55Pr5yjC3vpunfvbj7szpLvbG317C9m5VdxGb/wF+yM6ExGqGDuTcNurIuXjQXGU2/6wT
v/GcWGlrm9p34EZlmVhn24Hx1lJTFWwkzmQzSiQMrCCikeLMG42iH9Iqm2Xn3Wmw+0TjroWtwGQw
tFfRVi5MmECQmyBBLjpF8ggZmoGcG0ER87M4gBWQ6tL6Cu6artgcuNCd+4LszRjTq1oFjYfpVTsB
Msa+fRtfYhUcyXFiB0jKYZVOR56kdHoaZbk/TaaUwTf1ahr8M8y6ZfCdIzD2gAaHPq//PivITHhV
rsMuJzxwiWhDR2/M0qa/fs/yydqqYo7lNDdwE/np0zmSZsTF+K8G66KiG2mlnRmD2G/qcepz41oZ
916HgVFf+ffymNSgg5exMKVBYbO86t2qDWX+NQAoD0Xr90jdsW54OLFW3swCDZwjklmoRUDXWBna
4npnmamyUJBooUrVTg6FECPsCc1zBKuVipqzQ+xrN2kLlbj0j2wpEJNOyIXzmp6ktWLpvceH9nll
kGvPzd1BtaUzBK/m5So5Cvik0m3qMRGQU2khIOcgaCfMf3GezyWKvRsES0hWJRZbaJbxoHd/oiR+
d3rdJL/zdtSjY1wjHKfhKEvEz8e1jfFmR/sp90v/CSJ5hwxd0Ah4Sj6lGX/pdWYBdZq+nMVvma6h
ZT0kWhVP7JYrVgcu+5oqAVnWawwsXWO1RDPwlmm3LWvPjr+tZaD0MoeCHUZapLqLAmL/4uj+IWVv
xqFshhg3shepqJlSTToBtIH/6DzeAwguIRvQIIq9xKU04iyelhKr6krOyW8v7FyY6JcDuWCc4MP5
CWpQnbc5r7scFebKXf0/Gd0iYBuiyizEMaWazs5dQINNKmeqyto6Na/DGxF371/BvuY8jHllAOZ2
iUzUyLjhuxUESPRH0edn6RsEXgZCKdX5j8MuLmJFgeJSCQHmgB3KQ47M1UgdnhO51iqDgipmzn/y
pLgzT3XlDUwY2OAgQIy2QzB5qjRwY5xsyH8ObjM2EspE4dQRDLpJJlNFB417La0qvca/ipEVrOMV
I30+ongRHU+VYo7oi9XGCUMDpETMMW7AUn532c3iT/o+Otitx4rlUihIoFiLQBHdX9zXdGGK+dFc
gGeWB8gCe7gcwhUPkCBoDVjlUXiQNJsH/jh0rnpSY1WklEVFR5h+pZUb1AQtgHZAUtc8TD3Njt/2
8QuwpRqtp9iJBGUUz1YcHdqPN6AUT7BiukoEFZNns+vYow0yZQJzg3lqMg2kdWNKPmrKP5vm5FcX
5tQ4lfH7MiDxlOBH0J62p8QezL1cvpChtOWFcGdLZJh6Q7Q6qXM/DUrQ9GEhWuloV4SrdD4nBuvs
5uI6s0pY2ICAPcQYv220J03xzUW2CqGkybP4eGFqbb7OzhztS7hhVdHbs/s4c4XSy9Wjea7QoZbG
zWMy+4pS7Cl6VX60Pr30TzkTN/5yRL2j4okaveAaJ4jxydYAphjeuMbNjtmt42R6yFJx2Sh18z10
dL/bqOPdZTUrCQsWviXmsXGT8BYmvAmgcBkghnuQmWxNn4Y+DleFQ5LCDfr/11WuaMLXSJPIhYza
2Y17wYW1U1KAFRqnKG99nVHRowtrF0vEp92UCnUVu846XYUNMlCFfeptizfhYJV4cU/51XGJ2R/H
/ulHJ4+gdTSaX/k3+KgQTZWMuJYziBLKwGApNLwhRQW/Ix4LXfuuMJWcdedw2SPQCJeucCE+FRYb
Cs+IvjYAtqWHyKd+26HKbQ+BtZQRtWWCSoR1KKSPqt85mAmFvB3ticzLoyFHLYr3cixzKvKm95WI
q34gtaIYmOk+XnCusWH2bc6S5BNj1//HqK3MRmJ0039g58vXOb6g52whxZcukpXIX+MqQFsqJnX+
ZId2rGUkGP7hSCTQPxtERQxhl3KhlI/2sHQ0a/8w+q213e6wUC6JEYxLX+ibDpZufXAsUqHZnfNX
GwoxrXsJraNaJTPZ/CZRydJnfS43dtpmaQiYde9vSGkaRr+i3HW6bJ8FJigliooQAaUz9vunFSpb
iHO3rzTFuDntrWPD/qYu8zVCfaBHu8iJvIliQEPzbal8w7gSMAujK4AO31f5xeCeGCYfo6PyVK7I
u8PTAA4KQCecapv8pKic3SNnevpP0gcnlCrOSJsm7KElxFpx3u9NP9kpOlLXV3LlaakzVuM1EX0u
dsMmeDNicW7+nDzUWEmqG5163IPNo2nlbRck0l++mDuiHnLxY+i++penoBA8eD7hzfXkIcxw/dCl
bri9G743huoY82lnaEHwQTEvuHkNBpzGwzlWVsTiB6+wseU2fVqabgyXj/Q/NFaaLBgVO/iC+jO/
UxzXSZHKQZEH1j4gxHbHYk10Rw3W6F32jzZsJVaRsAUGEMkW9R1nAi1DHQw+biqLcUdiz0andEwK
LY3Sycv3yktgjKK14TSsr8Dafgdtx2Zstx+zFOxmNmfSto3ATDFpwVbjoYGk32ynN4RlMsJTpr8e
Ds2CGLFKdoNqyqSpelBQ/FcL45ceSPQjXHwIWLGA5vslZKbg0oyEY8jquEg4AM3nL+LLdi0YMmfP
Vj0994Dvg6grLdGQkbLguSEYpO+2mh/cda5/jO2jj9dkbigr1g2JdO2tH2K0fPl0gPjhRU7grmLr
wUQGVnR/8llMwMtoZKIHyLrtCfGrHFEJ+Q4d1sn+LPFI+y2DooFOyS7She6XUNC/GnkbMggy73Ia
/xjlcPqbUJ+hNQcKUqTtR6FMxb8NaXWMyClXSkJ8Ybf/vKj78pJnrM7qX+WisRRXUMbR6CaJjTmd
0XtPX/R4i4ZSEWmm6XE+I3w9wGowjAd3ryHQldyD/16/s+zqzBsASczPGz+It4nU2Xa0seAjhGp3
mixL/nz9LQwoOj17nW/48K8rqaryidl6NdbgWVAu87+1s3VHswBpXoJBkGIe4gLpIZLL67nipvWk
afeZhw5VhL2iGD/vN0prSBi7PoUSlX2egQpSYWtQ2+LvrrobpgOUt5XuBdkuZvK6tf94CrCcMLNd
HaeqWYKj9QyQS5ZJuQ0fWB80pz+7oW3sI32j5qRhIXjW/6Wima929EdPc+aiM3orAWfquaW4fZpt
lVf7OsnSnisenuusRv96rb7VSXiAd4ZOWhYCVUZMQ+n2adZMsDqsBD3vB0ib2EaYtBPtfFbgEyhJ
QHHPtkSbqesRQ6vOjnqlswRkeGFINGCCkKdcFrOEJOT+S+HXH0TCKfzSV7aTiK9gRRcOUPaHYCT+
R2cNBCjAD2Vxc0Tinq6slBuIVhmDaceZd0VegBWBTDbfXQonRO9Qp4lbCmn1sQnRarg6Vcdxd5ON
bPTGmn3qZkeF5O/EoMWwAz/GOVhT05/4GvxHKN0uAvLelZ1n6ct7VTJwVtDVIlmwft3oP1g3g0mN
lIZQDBrQmePpP3q7Uk0udgmRlAKcYLQTDFopOT3u30M9l0BHElW1DJBz5FOIzbJsPgdoQCSd9o4P
zZStZ58Fg2vNZNL+km5VBmZ/c5w5KSahb//w4k0Cd/+Unb5kow6Lq++XxN2KkJyoLP7+CiHVJoNR
ReFuqT0g816cNBTECP6xpQf3NmZNRV2OTTknmpaHK18kUdvzVmXebUhtQrrEWSfvXABTSxhoJDaj
bCzmqmzIQgR7ImMhQe04s5/EnqqesVMl0wjbS5tRKOmFZgCVXz0g/eoJkqFdePeuf5ItGfBUnw+C
A8UmckMwTNqtrECrH1o6tIF9XdtrAAL7qs+P9mGOkvXW789eHaXb6T/iQtDkLan9wJO1Mh49UnqL
vw7dei8EGtOuLwEkrI/yFC2krBT8Y4+mWaYJgWkVZD4CdYP/WUDe9WrlQWmVs1wYxHPQ+yKxVC+F
rurYxlYIwLa9EOpRlatcjBt5HMp7WaPF3Vn6/NqOv5y5qKb33NIHpHLNZjFAfr8Bk3Avzj4dR0nB
FNSdf5A18ByxsCWEummsJzIFzJ7DJiYYKoZyFTgbFCQzYXA0ZLvkbgdZOUXu7ZejLG0gEqL6Ae9f
HIaDCzQQ1CLbX4SU3WYmC+G8aHVb3JRmvSCrEqTMsPyunPmuQjVHkNfRULyXiSkMoy6QeEp9qMxB
4zoMIr+V9qetKpsXGDJaK+EI7VSKdSs2Y2mCG8dTowvC/Dx6Ft0lpJ3zfwjfSzdMmrBtBkWKWcNM
mjxMyRvL0FxlHaLRUN8ZBckTLLmkROUrR3SQSGlXLx14HjLeiyxy9WaxoNy3zEfQoPU7Viix2UXn
Udbx+ApaBp3C65aEByKuuUVeJqeE69acNVwWnMW7Yx6eFi0ih2PtkpvnXO7UT8A5eJckp7N1ZBp2
nHUcBXfc1XfC0xEt8PW9Si07UgBDtoVW5X9F9i5k6txkxBjw1DTHDMQIkKszj6UR2ngzNibATMP8
YBmhXrUKSd/iG1TG0i6pDPlzn4JBiz+uXQtTn/sX5ua0e7QY+a5LIcpNTi/2xcf28FYCDDXXCeNw
xo7JYvj3lqzt3HCJhQ+FAf3RxU+aV+8MaHKS0mYg/0RF0xdFWZWs9jacuvgkDfJhtvt3oz616V/6
s0lpAjoNWvBkw52XqnTwjvvW3vpQmH1EULl1dB9UkAqEZSLwV0IMf1lFRFnctV22Gfv8gLKjOMOj
BkOEjUrrOeN1hYPBMiF9zFwcngbc30NShHuP74ERqbCfGPiDAs8kOMgURBeXDbiCPrRIhn5j3RwH
pa3uLpDsneffVU6w+r3Y6Ax6MNjWaPJao+Z9HNJ8HvZkWSvocIdiG9segFktboSN/HxPas/ho629
qHj1kn8hxj04q7HZyR+k/7sdSVFphOJzEDpLSYSOn/CuZ+I0yNEb82nOLgRHSbZbFWkKoOZPJlp4
3+b/5SLCqFIXkBz9Df2TV3q1wLuolLsgig/6rWhoQLtPDqZkF/YrO/XLLf8/lHkBbh5kH1HcHra4
44h8wgyUaJrKAzo/CKdjRJtWqBpzHf23PAW3yTL1eSCGKMmpoZ6mcErkzCbLYALMibas6eN/zGTD
ohbU0i+shkFiulPCpUljcQwJJMZ4eMKbhag0m90PXVh4Jt0ydrEYH8W3fJQI6PnqCtA5br/QRBlb
pEid9vqo4OZpntiNoX55c4nGSSZTzPHBbjmJ2z53y9Rr9pRZH3NfT6dpM8ej7j8hhSB6kcfJeV3k
GIAu+6y1T8t0WnPYW9A4BUCjdt8dHdymUSE6Diw3IaFEUfZsV9YWDoyhXI2QSl+ypyRJlSKlYZni
mAwSi22x52iiRYYLj3rkOG9F/H1MH2rF8xt5zuFeYWJdFEJhVZNklDXfOq16oqfFzw1wJJFGFaZp
dg2FgElY70HQU+PTH9Eys4rdToz91P8Hu0N8UoZ73ghO99Pmy4zmZC4qflbduxoKy1r57C5ByuSR
NCtiap8sj9ifj3/nb3kZX9l4FQAFh25lACWdlFPx5Hx4tLet9wJPiqT3hkoKDlU9H8MGf3svXgNr
GY7Aut6siCTm54SWFoJ2saCfbSYkQaAxvKR6qZNOZKV8hmVCT//mHugPd+NlpTEEasXK9Yd7wOu+
UFA10IqhK2wTGtRmGvmg5y+XJFnJfmmU2xNW4H+NnVjNmTHLXSFpp0sDRLhWcIQiMkwGT8NYRVdX
nOzGz/q4aLXPpNwOrlDRSFOsY8zYvyWzKShsI7QMgLfbJESkakVVubLJ94ohpLqoDxDK8l9y+LAW
+AbQVn8h/oLPzmoMuyeO+6SBd1Lzjraja2jsVN5a/i5p+1lCy1uwDECVdcq0qdG3Q72eezeWd4lP
6wmNy1cPUy3gDW0tZ9g71tqTSqOhYNiIdICmXtXIMw1scTmJnumJd4PL1XKwl2zln+p+QvQeZn7r
IEjeCIy0TB3/NITo2QlIGGxCYWvNoRCo0oqJNGnjMH9NL1OmiXwBJusDTkrL89o2+3REkwgL+RzT
Pdo+bvgqSom0WtgWqbJsgVF3w8NRaUDTXAMovVskO06ML1nWMyxm8C30gV6Pj1kUxqwpbiypV9wH
utJNiXrprHJN0tz1u/ZWSCBKUQd3kUWerXlfsCCH55hCrOPUzUA8/hPzvFijQJHka4aMSrwAqwhC
GCDWMZiF82tp7jidAIhYgiz0XeSWhCsNlHuIZ11QL7o4fIyyRasIqm2goiA+tBCwOnADsVsaMm1K
b5tAjW+JKwuGvuY0ka1aBQYlZmVhI26Cr4HLR4hJYJ167hdkPhVrCTSYnQQStqDyWScNflU3xRPc
J6P0xOoTK+ERgUihUxy6+f5bsgbWrdvpFkjxULoL8b5urPqEB8pje8/Lqgv69LhKnb0UX6082A3L
GwaVb+xIWLG3C6r+RwgBCaJ6GQ/4iL4YquHIoRc5F2a99uioIHVACrJFht2VNeYhhCxOJSG8LyPY
h09DMo//4bbObatWtHEsjmRUvbMPZURx/f5PjIEeG/smk6JB0mYloVGDTB4XUJpbtURbIZPest0q
k+heXAFcywrZsdijPAhUxx6fP33NxGzVarmwSy3j0d1n1uuHppWhQ5uIwfeD8dGkgI/66rweWR3Y
22NrKcvKWmNVZIoUNa8SB+aV5V4wkychLbBKqYV0K7NT4azmDM3wREwCQzjc6/j4Ykab9J9+xZuz
QBiGuMs0B/n3m6G7SbVSW3LMWe4jJtBBA/gAuBMeFtqpsSBJSYfNeVcytX4mrlKvWFMTnVCPegkQ
gr50luEyymZalcbpRp4SvwM9AWS6CYil3TjzHmSaBYHzn5WMs1F8HRk+pr/IN9+OHAFcqGsncEvS
0I2i9OfinLg7n5zdv6VO5eG9tIdCRbQiQ8/lz117vdl9UDUVVyV8DAlT7nEtaerHgFSTmB+jejMH
Q5JV6XhvVKjoSLYaTsDsuIHOYIAZ1gEfl7JX9GJ5CigqV2hTgQtvRIPhBBxE728rV0aH0JNe2CK7
koyfvj0Jq2g6qQ0H3TWfpIgtWVqrt9XBPQc9RaHIUB3XDXzrIRuEyyEbA9/XNI6jBKIk/nU+w3HE
BtYgmhJuOa2yx31FMMifkYJ2a+gx50BqTHdoPw01ToTZJI6NlB40uYHKwyaP3fLn4IWhtw53XzK6
cm9pu9+eGm/lFUznfmt5JP6YmmuE/ChfLRKMofeyd9U9m2S8HKpH77mm8POvweAFG2rV5PsfmrOV
Fj8BW7Z3S7G8VEnhgLh2m1Lt0MfRKBFBmqHTBkg6hqHO9C04Aig8SbanV6TUEzBu75+xJGLIgZgn
636jhs5ay94XlYvQHTFJL3rKVNDuR1mPZ5wM6Ewil71+KEcJeIj3y6KJo9eQq6SOmPgu2G5VFa3N
tyGEiKhibWOUdUEH6EySYdCnQ9SRkfKBaKQI3RBtN4ayhuhh0OxPNn7tPSWsiMrEPiaXcjtE74s2
qTiBR2WIC//bP0qJeVY6YYWmezdJBvadt4KVNu2CGFIlbUNl8TvlHUGiw9j75a8jX8jlkqwa6XaY
8c4NyJvzOu71c8S0QAad5Rj0F4fBNhbhuMe1RtmrNQ+su1UBh/tTz/li/W8hC+hJ3Tm5DpYYzt/F
tcVo5TUrwYEcf5cbDsrZztNtY4XzO6PQkpa3LljJRE1cGbYbfZgwlkVgmYJdfUlzz4e7aa7/TVvl
nAlJZFsccxh2mdsmly3FzQP2RoJrJKi0cf60JPrD6ymGhKgetH/GQ/xK8+r7ca70NwUnoeyDOqQc
bQw0eJAr16tv3aIRgNzpMfCgJ4td58HwH0/pK52mwWpPJUuxHDfVfeK0IluIw93XjlF8L3XHLhl0
qkcoaUJJZtw1T7Ce2w/380+rjvnzxk7xKbl07PhKHxtPyMuVJgDL+1LdaY4NB3HftCZ1vUzGNg4c
Ez35hnEqm69JdBrwmSAub4s/7ph+i4pBjmlLRJHMZ4mAhSdQLmOhbCfJ0N/bqcT0FcOfsmPskatZ
nEDgyje8gpdyteznvG8GxtJyd9+au2jH+r4gbI7Ruk6eTzfpp7ZgMiM763HaNk28QOkdgq8OzudZ
xu30snL+UQ9esjSEH21kWZtjM2wBvDTHz72UHPfK8rZI2PmN0bPOHqsRfmGZHCd+ftVNFZKXH350
Fr7gAktlSB/Ub8un9LTlSUsUKUY4VHnAZaRqqhFExDkTCyuazzzNBdBn/C6K+wYwRN6pAr1fCnvR
sqnhhjRdfRnL/4NbVoHXvh8WPlFjeuj9eml96ipM5CmBcmy5fiCvR8WVP5bw4VQ6iNZ5QlzvRrlY
L7vOrEq1seBfXVOjgkb7sHAbJV8YLvlYHlt5NFir5jsYdUG9X1GiUhwOagInSTZStrBG0jpUNOrC
4XU4pUKaMe6TsxeRgB4MIYCl8CLou8eBUlxnZd84rFG4EhiyV0EecVwdYUEhpddVwLse9KvNqsfn
42ivuuoqsBdv2sOBp4lLeYguC7SrBa0UUtqsxvtDZj2ZGwuPqFPMaAzsaZI0ANw56y/nY2FiRzhP
BJHgTYMIFxCCgKKPFAzVJgv+72A8O3sdyh9KEPF07zY6bivoW17BuNwnWxTaf7d31mnI54pygZif
nnL5p8siYJOUlJ4iLQFEL5jmB+zo9q8CNjIgX9aDpdPVGfRD4JHtWtriRJ5Q+AYrTHE7NJMWribG
DUHkg7f1JuNKfyZGdtVN+TQAFZE6YxOewl9jYCD3PWXvDkztgaKGgph/oHWalQJAWp+Ws2BuxK03
uCWkNIbevfJ/DG7qdmg1gaQ9kacp/4P8ezhkyW7QjvNaVd2Gd12IAcKHeWsedIDObO002YlSpdyz
WQfArXEK8yNZ1YGAZt+n6VVhPoBhztcicDQewXxp8VbCbNV8OU6TApZhTXU22re15LFBIYdrrEI8
6Z3WSUi2/YokIH690MAPOqfGIBlKuaX3K5Uei9Vkt+zCXnDRrPHir3ewhv6sp7TCdVq/AYAQvs6w
o6fsX4eFVUpkGCtl+XdbKyffZNIiRf37qWQXT7RfX5LqPQ7fd5DP1vo6VibP0TqK3Qj8vOPLbHEg
0Qae4QEdzi/gEc5xqYU/Cq6CcZcQ2gp/LQvIasTabPuXZPOCPm4nVLH4Mp/BhnZGwm5QAifokSNj
QMedxAMWNENMFk/vrHzl8NDeTIawCqrARnmm0Nfh2Imlx5RIMidJmBQY9FHpsR/8gqjVL67qtqqE
caqOAq/uONDhrJHpvhlo2R9QiszrgNHvhrxo/IUjxdV4ht8qis/EgteK6YtemLVLY656fjuzjqoh
bIdFtDQCX6j8cPHreaAJtAu/RwI1vEUXE71Hp/Y/g/vnX1I9DZ7Y6+XtlYYDN5IsW2FE7btp/VAU
yyv6npBpSfGzJDbs3YJiKk2h3H9+jEjsdQ5l2Tz/xNe/Ens0Q0slKnYimlaFgmgdHLFSCWMFMMMT
L1N0Nu2UAKVXL1XjX1MtQA1RI+skeo9W0h5jNzcFZCCqV5xrf3VrgxchBQsUWQ4JyErwJ76alqsC
VSDyt2dwBdYA5h3wduksAcCh07oV+LJRDD7KcEGwAI4jbFFLKqGU4K2leKu9WmVdrsm4NMk3HUgJ
HqunPvjVLGTjxDgSR16Rp0wfmk2M6FeGTgD348zYSy4m6NOiEovMTAqrcvFJHRERwKqNRDdi0bL9
1ZIbQvldlO/phxpX6+eDcG1QGT6k4ZuZlwWbrabBDZ4fWn/+Ud7X3d2HBM9PIVKI5gOcTrstz3pU
LcLTvnKVQQzx/EfwC7gd7VbNBLnNwpHdZRBjOZENIRxhZaXVjR/UUUQLV99iZKKRq4MEwGd4FuNA
mAb+2AXYdyU9bn8zD1+dkwQQoeDh3XADNu2uXCC68NzYN2oqGJ7c2rStXsUT7bEUaPjInl5cGlIu
cwtk4sUpj6qovbwDRMDGHGLe7LMjr2q0krHUUp4TjJg6DebWLV3YENY/R32lMY9T0g2SJPn1jU4k
NZPLAyQwfG45XNSz6b/QkhmSbkIvY7c+AZwFdBTAAscd8k7naUAKXZRoTiAaBdtabuLj74VwCybp
A6+pAi3Z5enhHUCuphkLDk/96Ql2QD+jyRtt78YoFDoowcOPJyC5IMnxPwhcO7F1ufgRTPXRTFnI
3ZPuGd0IZfU0SetKj91hqfgjBXZ4Z35LnAYbymURJ/6Zl1T/3Sr0s9gHbkbUgWbR21Zaq5mp7gO1
D63gUIuARG9fY1MMxUJxG3GJ1vFsbzh4xP3rtvWr9qYyNx46DzeWP3MpQTkdO8DM4BZRxj4njHEb
6F81+VPDIIeC8Asol3M9sH5gIknPWtCChQBPXzjlPp1EoT/4DhRDpo1iSb1ym2jB0WwPRiocQTjQ
8WL04kdeH78Q7dSouy3hu7MnbJrpC94MxBh+uV6cBGCA9btlZbFQForxQ4lknMDC3th7JhAg7+Jc
ahpD24nno6m1f2E2sxnx0O+IGhkDOHHAT24tG8EZSyQ4HB9+AEHxonBndM/xYF+C1h6eLfBPKYsf
IGzhkkL1qw0rk49vKit/krgORv6hqp3sWwh4uVjTFcjpxqfL6sgVszBZpFRQtBMvTO737+8frHBd
NzWi6alFlKhZi+SrtahTwmbKqahJ4dHbTB/sUy+QPojw1grc43HrhveRth8x6pOzoKMK/kydpSQ8
9U5eliRAk2g+a3HTbVyA2Eij9q/IbCqgkEhNeUNiTNrIu/v5dtVmJGiCt/YbGybiTA5bWsI7wcwn
wvJtJ9kJEpiAYZPldA4uRzqSSqOBwehjWiZXn4ce4H+NZlm791JtuFxqfR8roEVP5W0rlLRWt2ps
zcV1jkf2pxxAqGfIHuI4Nsyi70d7zgYWmqaVo1f6TWcRZ0F8KUj4YQ0oXmER2JzNGTWlnyrl1JmJ
+IycgYbsWuVRy6hBB2T244Psa/fhO5ASvgGXQda+q3JaHJhLEtcgvTg1QzhRxB7vOPHRnNwaNcOD
iG8Sm5NhSx1kB1fZYYcInNoSed4aEGUOnGi2Q3sEckQCaBtqJ5H7XH39QQgpzC1Qs4EZocCuocIK
Vdq3cTZCbUOxDpAnPLw8jBZXDrrnypJOcZWnKaiD8Fj3xUShYV9SOjyk23zYYZSqxTEMkCexy4cs
WgYcwOwphp0x27hIxrLuNJCsQKJSilD8OgCFjoD26RPn3WVZqwAINESLg0B1mIe2YVIHtHNdddq+
BRqJoFE6L1PCg7nQSOk5CDRY/fCOZ5ozyCdrA77MRjjF94xnTBPF4UqlIDG3HN0MCWh/SVwku3co
ZI26ucXHTu1urNzIH9yXDvpd7SQRT4clsnE5oFPAQSYbJZhvAXcUu1xVplkRoYSmt3y58b1vPoOl
+qNh1SwTfcC00DRsI38/vYWLyd1+guPhDbx7zzBhrO3hBPZ+7KiVHYePMWFFPgMI2NjMq9RaDsJJ
0gYvU7RL2ENCyXzekYRCQOXhzI81VscVye+ajDa+8KST1zQozfVHA+zilIsh7btsWxm6XjKEox09
opbjTX32PxbaNraXKHVwOWznwMNFTMGlSAVeIR6DEJCklamJHKE6yV3zWTwb/JJ6CNH0+6UYz/l3
WA+k7N2ooJ8xHf/OwubfuxZRrL4Om9OiG0/mgzLw7rbhmbVC+TPdGv3TSfz+oCkucE/55c+pwP/W
JVjHsROnRRNJ4+ArrsLEVCEn0yS8+axSUr2WJ49oqup1bxyMM7EtwTgTTPAFqugfXtf/786luY2b
4B5BScdEAjt+uuRp2hGrWhwD0qFrs5vZucZV60oC2QV+pZzRsWv0thk6YN35u3RlZJ2a8Uam4kuN
tCaQrXf5phHiasyCPdN4PKppUam0sF4hPThuoBnVsj6P6lEUc0ZZWfxYKkykbdxKgRXYjobqSK0a
jaSspxMPlCAYqpkXSFRmp7CAYj1aJ4V012tQNRgmd3yzUTdFIwHbRe/HLzyCLb8txmQEPVdB9TC1
O7VIJyhusYkfJVm+Jh959QkzURT9hcWlv2nzMgQ3YimxHTGWqQxU8Y1WQ+geYztjrWldidoSoAW3
Twnz+T9jf59cPU0DqN0qgxh7lYk8VZHhVgmWHGOAqF3bkhNp9SyHyvBKgUPmFnTdcH+vDUqWcryu
mvB5nc2OUr4lfDkf2a3IDtIE74z0iT4SbukquQy2wbAa+575ylG+oxDPCCW7KtrnnXRs7rFosV/K
ovn2PwZCEHDXXUp6K21695xhawiTps78Cn1+SM6h6AOOg1bcywuIgmuIkvQtNqdnFEv8QPbmT5b6
YvuYBRUyUyGK1059zemVlbwFkuN9WmUauCp6UMAc8Gof24hSY7NB2+9iQwEQgsg1UYxuZ01C8r2P
bEO3F/E5Gvrw+7HmNPX+zvjNzZ2pV4tvTtOgCGOGClu+3JyM8xY5Isn49b+3i/ro8BzKSNpNq9lz
egsMQ40h6gWG6meArqxJUux7L5mKmUQn2oq2e0lhPiKTUrAcHuMHdPL/hmnIQQSoKpZOuLjqk708
M2IGzsFGd3Yq7dLk7NDsgtPsXhVBDJLQF4xcCYt8d0eTd7BUheiYfGfaDplhISfnlGiUCdQKehx2
Q2Meg7bXomDI7JXnRwmcDV6H0lxGex0ixCXX8TdU2Mr8zB5b1R9ENyNLlaJlTV7aFbfOxpnLkc3j
vo6CzTLtNrH6iSggt3m/UStXPenspqvNz6A4zYQ6dUUpQMCrnKCx+Jn5oCEMx2LqeQNVQtq1qCBn
HVC/3rJVrw1SJg+6OGo+xNrorXL6IRPoJRmdB/UQQRR+vMhPyYo3rDoLrWD1aR++3JeBWepYtbWS
UEbrsBQZJFTXf3xHlH2Zr2f1LAGpN93oSkrUw5tx5kziNnX0G2rMeJtzIOdvEWJbqDtXL643cqRH
SfpHtoGrDf+8/DS2RerJ0+zahOzomVcKD+LtvU0a4acmNSO+/zvcA/A3Xf8FP5hjik+yxA8vAYy1
Z9Lvgb07Mpq9EoWW+oKM17HGEvrHvIUatGUf/yiiOS7yqMPK8Ax1lyDs6ULOL66W/cYRXfwUP8dV
Y9aHt8O1KiLpHgXa2p9HZWrz4kRjRwmnuobRXttHCmHImtWgFS7JYiVnsZe0izIUaafqcqPdlV74
bTo8fhcRHoct0qIbiDb9qmRhZkaovmZVaY0MZLc0XpuXzxzIC8oyMWi5bDDQWTpVBesVtdPhUKGa
9z23TPFQ/gJV+185lpZ5RyRf2XKFB5DFUCZ4x6tY/TUMkoDnV69riwTjVhamYEfc7PZUH8qYwVd4
CzaSyUMZuobHhobJgU6N77dmXE73G9tIAildCMsvV6NSQtDl8d3cms+1MYHkC2ifAk7pelt4fPN8
d7svXVCLakuWfJ2IDxl3XzY++9NoIs5gECb19GUvm/ljbT//tq/uzlqMfCrpy99o9dUfoRle1FzQ
49Xr2DqffnijqNMLKgyMqSdO3+1SNcKJAU7okTgmPLJGdDOIsYdvt7W21XNvnb/Utlsm6/WVcnVH
VSswY9uhEL0fDBDdWdnaO8TaJuKbCLSP63q++HVxKGtaxwktmOIWzwcGsYiYjEKHSwcl7mMExaFM
RW3veFoWoJ2lZW7h8567fsXvxLU/ByDyIlEG7ZjRqN/mVItOYdOmcXB4Ix8kIIVErA5sZRqIqCWs
JF6YCriDoHYjvORa4eN7rqZvDir+EQ6USbDA+uUpmbKXR+iBUkuMUS3v0diY8rkNg2N4IGN9lSJv
bBhlWMFvm03TEy72/QMuhYpP+p+2eR3kbRf2WehfKeaRbK3GXi/5vS9ttguTIDGqxorqiMnQKsMD
cZJQTEMXRRgzTCCk5xx3dNhoSyUMgdwSmk60dPjRSfpKLHUidoA+OIeVaIg+SSbGru9xKREgUL+q
bJ2EKFweYFYv3SVAryiRahF4/8R+m4XjrZ/xev/iMLZr+l38XO0KOEEPq0R0juP+e2DUaQa5Lyi6
lFzCvGtggzyli3H2Y+JThCgdfy8r6hPY978Jzgm6ugOxM/eRmYaxucOjGS3df1aVOfZasohyF3SR
2+7pzZQfNx2Sny5c7GEVTLjZc+eYH4MJJsSO+78gLv3Ok563GCRX1P3471UFejKxA5gxMwZHwVkH
xK+cYbpojcDypUuMBqaMG5e8Z9lV07rfE+rTb4w0NNUHnCYvIxZrI/haGmMoBcdsstgJu/IP2yov
MCbj+4VQgAFMdbyc5zS60DIpD7yjmtPWtB8MZRGd92FtXCGF/Fh2TBBoMe4RZ1pxb993WNPslzz/
ikosOC7V5EMmMq5x27V2p3a+5kXW5gw+xUu7Q7g9wKzzW6UFfU053ffbvedDilnNXydAc2Isn2X1
voTI7EKbSZxp7GIwmLtHRmUphmpArv2gd+WqSa0yGO9v2zE76EkUTubSxNe/TRzFw2iMYYdYs53F
ZnIUHnCAUEdMqHNf6sglPeYrrGSKxRsqP5vOSFu7qHLW+oKSxmyNTeTbBIbpZr1EUyDEy5VFJnbW
BLx7h2yqXZoNozPBcXn1EwE2mg6iELcmBOfWBnSqJrWlXTUcqpKlEqeKAJNjr50eiz1rliUrk2zS
q1qUccqS3bBPjA7QFI+AVHZmCe4pQyJwaJUIl/c2isT7WWXwVfpNJoPO/kHufbQrE43sRcGZQvCI
pCv+qUF+HxjjH87O7ERh3543b8K5GffqvZW/AH8506f9hRbgrTh0zT1Jul91IJOmVqBj35MwrlxT
7KHa+PMvts+bBOs7MSkJDDeI3yzWbLbl6dtgS/HYOuQWv0BWVYos3BX1oiY3NHmd+wSOrTVyCewJ
imc2SjJspKmLjtPHYECBxNMsFtecRqivaGHcTlxerRVP8QrPBuQqzfXhrGg58heaHPPk199CvW1R
oopVj5nRDp2kYoDzuyAxNbGxIxpgQ7s7BTcBM/u/68Ti9t/AIMfCNt9rEwq1Kcib1ffjCzE2RNVr
QpWvQvihGkj6Q5Hh1jDeXztnIu6l6iFfk1Gq5FOUI453SSjvvuwJ/k43Fim6ZlICw5JzEIsO65aP
lvSfvhI0dcP4jAZnO0eR8RyczsVdV1+zC+f3syBktEv7JwiNsYHEpQa1zm95p3AjM56+uzhp8zmL
Kc/fQzPYSY98iHHPdaGxXnQUopJGrw2cInOAWJpjWTlAK/+99LFkfutf4owyBk0XUg7DfY4cnz1b
ueEjAcxFlztIDj0PodWTC/9h/KJ4OYU75SZZjZhmmgX0fryqsE1/cj5dgHvsS7QkXH1PrcyVrFJc
25tIze0bo9Ow+ZrXIzWBs4P5T+hLl0B/IjyOaHJjHx7Y1btbc5FaQchBUmeY2mfUg+b6YYhI/qVP
PmWbOgwg2qlCr7B/UyT70fir1hcPVp2EjD6mxj/REaQQDCQpol7SXAIkr17BbvM6cydNhi5kSMlB
bi34y2wQXlEF2hh79o4+RtPvicfm+eS3AVvor9KPuSbSm/eqvoTf5v8/4df2Q9lw6suEYs8XcKId
7+TX2TqsZq5moDXud5MJd90Z1rRjA2Cb3DJkGTCYclcxPU0TMGe3bMqoffD4er/m5RZEJqr8njR8
SPPvEt62AvbAUobrAGr6fjxmCNCo1ONUc81jCboIxSy6qetpV3WWrNKqdXnctuLolVd7TvoVlb63
CtoDppfbqMtx2Dish5tTBGVJLj4EK0MlCLg5Q7wvm0flcqoyekWR0tAtPkgGbBHJLh5UJo7VztA9
Eimhmxwfkrb3+tsmqpeHOGBacKsN9aB9gNp5/JvBpgxjfnax6F//eu1mxz3lg4EBxYL1zCze+1Zi
IuGjZQ9yXdvJeF+uGMDo1Dg+V9PHnkGA11YGIvkpo/ueT0sHxJEkqs4Al2CAj7wYU9ovmZkWV9Ra
mN3vV3dlbMSt5R19G+IuozR037KM1lh7em0azLVExO9+bgqz4cp3iz1VdNvp2AhyW2ZJBh7snL39
mxTPxGMarM/bHOVWuShP93cXXcPF9D5uRvccEQ0AnLiTXEqo/tczaaaF2lN8t20HoVWYn1uE1mUB
aOjnIpUhFtJ/NWj/bOOqYYvdHM+jhz919c8/4WWMKAc6MxXRnIy5Z52KNMObIiJb0brpcmXRCaZ4
BKTgrz2Aj9F1c6dku50srZZIQA2/11WJrVqpfAWgs3vidWumG2kWsst8UhqF/wR2hu1EWi2veLku
kEHaagyYAqJUetC0SmceqTdP9o8+G0YGl1n5/huSBhkIkK1+jgdSp2yIcdi6fuiecgO/QQNU2IQv
8Q6e9Shsj6emKoP37L93xfu1czE23pAWwL176SqD5Q1cqF2Ego7LVcf0YNScD9raRwWQlefYmhV+
BDvs7UZGg5Ry3D8bhdlDIzFSLzia8pOS6zAubC48E/ypVyr3FpA3gk5yTZydQCDXi3iSFsInEWL+
8fZx+ZbOqJN54mqWZlrGyu+tR0RtGJBCQNJxwLXR+TRKdG69wesJt9no8tUJQfy+XMoQeOGDhr7m
jL7Bxg31G4HnN9uzPmKB7PnHbMAA7mxBIV4aLe5ku7BjcEVW3un0KzqJrglJS43F7GEYglipauYF
W9lO5Sgp6qnodU/1UsvM0rwqMFda2EmQtbhJn4XQol4Cw+VfF/NXaO4z172qqR1j5QgOHml2qo+y
6qc8jpWEF5XvuB1zntpKcYfst00UR+KP4VMN8LdUE+7dHmy2KVHmMg224Bx/wTqpW+WXZqsOKcIT
Rm9FxBpF/blGkJhOXMiy5H+QhEx8LkiX+i0Ej5ItfEHVYM7OwowHWsa30mW40No8sVgOBuL1oudn
jU0GZ7fDLgp5S9WmSmxsWN11i3OyEutoCEVGutX6l5L/ixx08frTPu5kNeA2A3w3aYqS0gJSZz8o
HrQ6tD4wL2thpQvCnX+X/drUNp63u6vcOV+2sPkLekzJd4s5eIRjVopOOBvDbt/Z7aZyE2zlWTDy
8kg7hKrFqqdO8RasJnIeEh5A6iiQ1MbEHDZ0sTN/LpmLz+buAXTkFpnKEnrjwwvTtL8F8B8pm3Ju
DDYJBAgqBsYjf2lTa57cpl+ljcxkGaylqV9XoJtiOMtbc6LLeK11ZIDLIRV4EEzx36wtl32EryPS
gq0AAaNVYWSjX/m6BjZgJtXK4Ligiss+H/4I+DVDoAg7AdSyR6JSdQ6Ls+eVIlvsjU5dhC1QTinc
v+dgdQpBntb7KCuoZ9u/wA4OCb7JbcKWPjFOvM4RzMya5iQB30NYnv/9x4aHD5c9X4Uucaf2wQAF
Q6RAWytpICsLb1OMb2LuvsOTe84aDvczgjTyOTqsFH719Uj8nouFWwRbFM3aH2Ig297qk+W7qhR3
eIgHUfQGoibZlhbkY/9+TtYwUOGuM3ESO9eVFeyySC0eKWeeMTpa18V3BbAq2Mkr+W3h8QtyrRkU
nYx7V4MYYcbUk/MyiTmehzkbSA7bQlV93FpiylxSKBN6+0z69LXsTuiXhvAK/LtFLljOsyPspJgs
P8WBQYY82z3ZcxdNUSqh1Es5nzovHNYjqqYTrTBjuhhClhKQg8oLQob3UPqU701itxQr0jQMFooc
6HdjoaDm9sQnnVSAKWt6HGfW8sZMi2YfrQIDRrUSDxjIpc8iHQx6cNGLZTxGaANv4stH8aTwRpCH
akjJY5fJ1Shy/0ywM0doVtAyt7zBWarqkDKOYOFPlzYTAxUV1bioImtq8ndLxnoq4v9613JRMIi/
ieiI4xiyabxYRn95+1pltvLJb/rD7d8T5SVb5P1f4Wemyy4UHueaWdiXnlq/Sq64XxeCdVI1pP7d
xYyYWxFkkDW/LdZKXCpqSoY6YQWYCo5vGWcl3Vbl670NL4RzAIInQFGIKzLV4l/iveVSRqpotYXC
VEsin7VyaNDPyuzZXzmNeVV+dirgF0MDN0LwgsKGQexXlBkOplg0EmAEo4XMZy2BqdMs39+g2BiO
/Uhb5/yTrOFSiD/B40H8QKIjMX7l5u2XYJZmrbe6zF3ji2zIW99rOL20xzcKPLJUKzFKVe6DwnSN
8q6/Nf3M/4YP67zlLHMG81bBQRkfQo2IFhI3BsoKj6Sba8ggz1LtG1VAVFpJh7KqI4kqD14Fi5Mn
7B22yqEUreimCxpX94kOOu6jfd8ICvr70Er2nHWh7En9KVbbbXIlh0Whyk6FaHcKbsCzA1HR5WQc
VkCS66/Ww1NiTSpGgTZY/RqyoSHsF0cWGnI+FxcHaqiLrm0tdP1QluxgNfp3KfHof03W86RMwUbE
UpfZ9tSd+oIiR6oIu5E1DQdCGZt/x4mXTsG1B/xlH+egh9fBIaZsmBZHsUIHNsL6xiPG61Zc/oJh
VlLq1isOz107ES1ovxY3BOZoio9IRDC/njaFmIEuPWfF8q+knKDu/h7+G0ddcYuSaNUoutEadYEV
3CohY7Eirn/vGwiZXfLJ/XtEZXBuATBb68Zvi6uMC+R1KKZx/RGNoZpWeoUOJ81TmJPbHIUJ/pX3
l/X/Oeoal1BBZFlsNfLRoEcdwNbDPqDv+x3bqqnNO1du8n/pqHEa1Zcpsq5PTMUzAqp0NJ3NIfZh
Tz2HLVH46iYXKHOpAhp7TsQFOeeVw4OsegcJVf4OvK3LO2ybS3XYnDqGK4R6EnfY+VcajLPcHh57
RiZcpJBLgVpY6iTMrpwrPA8OhVnyui0Coo2XfVEZNePR/t3jzxyi35PqiQus3pk4MNNLfA5lEDRr
MICiBiDYWSgJfbehnWhe8dc+911hC6WS4nqdTFAtktdDlwGi9r479uQcgT7uAiMroNrpbwUykiva
Dhqe9C9Qx9LZMdY/57aPyPecfw+wd0GyKhQbA5zhEN3qWlDTDq4Xbn3z/aGpU7gCjeNRj6YOEX0u
l8sAFboGcyRwd4WRtTMlh1hQNtbUvgNDHr64BIVs4saZ2qdcrOQrDFSsWXum2BHjsTdX6YWBI8wD
SSKyM/dGZ9vsCK54lvYwwQy8m7Yjb4LA/mYXHdW63Kq6RHsLI0/YPG/VZVV7lOW1OaXyT192NFmR
k7iAqznDy+MekUa0/Ny0FQKCpEDoK2fsEHgPDGpxWsY5aHW8tFPN4SrhYuQxB27ftwq58/XVurNq
Xu1Nyfqb0clZEzIzBx42jxkgYA9xzbm/Z7/u1AF2TNegZ/zCpUYhl3OsuLOPFEhWImseLOMTyMQh
Y5tzpJXo9qV7KTyhcHWOf3LsepUcHB3pW8nSdGmyaBe04D2EzeOG0CdPnDCPbn/0C6t9VbOFN+mT
G3nBVxwoMypitgdgurnJI5Ev5ShZshsavjWCqNl63euzYAmYqmcNAZSq1Kb6zioORIKioKPWh95i
N0sPFO1R1rJsm6OJAVTmxfyhoAA0iKXmjzXmJbkcl33ud3dNxCwy8s8SUrVu4UtZMKyKH41v0F2r
v8Wd5uxy+djv/8HHsuXOqGLf0hL/h3LhtYFlWTjqmA4xjU2AlpO4SQOKKwy7FYT1+h5i6fDAp9K6
3ox66KI4/2O+08c1XymuGl3CNl5ls72smMo0eX2lWDIcMJHgN+Ly/UhJBHoTygqWbtvFhGZWAYfM
vFaXPR25GiqWFi6QqYiOxgRLcQfTqyivN88w3JIBQhYlwRBLnw9o0lnHFW5i13YZXcx/hwutOyyy
yqHk4QY3BBr7MvFlK5OHl1+BbAU5HeHGqxQZDeL19JSOko7+6/qOufZ9CQ/YJLFY5rTS1zrEihtz
oGvfXns3wUvnbCcBmPfQ8RD+/XjnWo2ONLZ2RnhN3Ea2jNCQv0/JAfU/P05NX2A0kJ8gnEFVSqqr
pt7ZZESh8kVbScwlpq7cOS94Csrs4Cj6Ub/UeoXp4/o1IcznYuHOXs372hBFs/BD73o2EXrdiKU8
zetwz+u4RxP0WoDSwihBLd9LA2MUM5LalCIrBuPwr5efv05vUEPus62RcutN1KiNq5L73qTe3yh4
dh2dCZIkoj6QjmoRhoasTVJCMsJ7JtP5T5viOlWzwZo7+Iv3qoXcpy6eH2p0Zse6aX32PNrIP9XG
DioKGZlPCa6zvM+Nb5tSGXBPkwcP+bT5dR/ckvfO09z3/xfBD7zQDtyD1ktgP7GhT1m82Jzri76a
s3cygYVRqITrF7pv8odEEe2LmQIfWNWGm4ditzx8lj5ePF6a/FESViVmfkU1VX3NJ0t0ReyantSN
U+EvUwh5D9Wyx8Ytadp24uljdUyahmhJqWFBJLPeMZ34fePE4m7TPVwXO1HHV77q9udWsDmoWScK
jVC4A2/oWlMZrwDdIhnr8uIEP8rf5UpWi4ejK9VxsjL4dNsJEKTdAMVJQujmkr2gYR3sVwKQ2Ot3
WihpmOOFO1+R1FopPpJiq5qOXmtlHdLtgW0Kru7lR/uxi7lxhQYdYgv0KimqoCv6ImcvXjGM8NBd
dWfViYzJFRrELKIJwpqKw+3C8IqvIgv+/f3xe9dQ7qNkaqYxij+jgubYzyJ+zwwP1BHzj+6B3y3n
6oamLHhvfEBgmH9YTwoLGjYtT0QVSZl1mAVi4q8GBCUZalOLFrEUpIovdltRVqTVepciJDjpbNY+
iqgKY/H7Vj0EqnNFKlwv48VLyKrJlLNuzwOsAS4ta+rckO+haOXhHGET+D/wxiTfVv3x9gSTCZ5D
/BEEY4CYrLXdxgnmiQTdYfZDqlyFBsRjBgF83S5weHjuBvcJGwSSvPOqY/lfg7ijzW+5/xKpDTb0
HzlHrCIVzRyCsZk7WQ/vDolZC2tHfEKj0KE+TyQiN8TaZmnyHNA7DQvG2DOtKa7HK4stNE/yBF3U
iYlkqiRPWNdmvZg4XO2NKvG4Ixy7kGPghdjspHAgQoW2EpGMyYK/yb1ZEWctvST1Z2lFAqsES+BO
5j4pbjCGpu+CPyUGJf4XL6oBlDhdFDksMkzrMRqNue+Q8jQVKAJaChkOoZVX7955PThMbmM1OUqo
srmnm+lB0UHva4tuHiPlJnB7qWE0zy6RyGfuK7d6JIOI5tkixLU5Z6/jICmoU4WDbiZWxbx6lzya
QGRVYusw6XHONmDrD1g5dm8HM/+WaQmkBsoTXQYWlNCV2ieTyfoMB+lPl0+8BPxByqfBSo8j75Df
ob8n6iIRx5aOVF7ejL6epj7ke2BnV/Ur3dnPg06HxcyFiJAtpKs+gnYExnfo4H+Gr4KOe0B/+CmJ
OL23FhcxVEdahNr4afbx/h5JMAVFexpkx9eWJhfl6x+pJoNHiJ9x+Kap5dFQEkRsl6HDDatnhWwn
4wee/DBivOQ7V4+M4Pg1xRwKT8g3PUeX/GTs27aXt1RtBhA//P2Nr/tStfQPPhJt7AKOmH5Xbzy5
VIGDFFApDSXEYzBbqRi8AT0Rgc217H7KGRjpQq3DEwd9WGC+uQg59AmhvLJTLfb54a+AyOozPs0u
o0qSf2UfyvFpaMoFqTnOW5QWXX16Gw2FeJpk4IMFkgsLRCBlwZTvapM9BRFy44x1QzIvfzDIidXv
5uo1Y59iGodtpgxMQ94bLoVOMiLtaCOfUZGd84F4C6rfNJ7onjDgGk+IRs90hW02sLcDUWJkWkgG
9H3gTbH1UYjhd8Ii8h38gGaLhRb+X9NHhFJThJoknqnOqA06orIwXLBrd3CiR6GsXYMKAIhjtmjd
2ukao0WsWRW/E2s+qpE0qt3l0bJ6r7fTXY4Ou/1H/wCIkGYsl0sufJ82rzjhIXICssLuSue5m4pU
L21s53m1u0QknjUxlAoYX/WPkqlPFV7wwQ/OSlXR3h5yrv9mNQqPR06NhzmJyGxiI4vuYMXjNIcj
vSd+19rjNTQ9z3YC7nNGuRPLikt4+JFnw9x49Yk4q7UXC8iAcaad/cwxfDnKKdDpX1t/Np2xY5HT
PJro5T9O8IM42UhgdR0gWnHIZo4NsphQYnYP5pk1bdK662FN+I8F7DcMIMRCcY78D/VeYg3+QpJJ
5sfMen39w37N3IHsaQWll3djCcW/9OXXu3mlNHLXHv+KzrZaY5eYF+W/rEIg6I1ug+WJZo86so/F
GY5XooRaO02MjszXritRGHyL2dyGLtiQGparFpp3cei2fFOi4092xxI4iZnjI3mNRc2WWz441Ikj
5yezZ8tYC7MyzC+vW3LhCPR9PMgjcyxIlGbJtBnWzGK5hfIyON0mkOnOzV2WIEC4lPj0u/ovK7ix
Gyrj4aYBvs69SGhnEdf6mCCQe6xLFgxg/A/lnea/y9OeweKZUnbfYXCxBMbLPVmwTBKE6lq/73qt
uuu5AaTDunqIe/3hx160P1cDAevXF7Unfa0IdjE708LsQkTm8E8GOAFq4HbDL6G1NE9KKSbsqHEc
LZANGCvw5QZoK+7Ko4eL57ave7bySv4gynoFVtn7TUIgjhpNI3jWLxL5PNcODYaeusGzAc35gPAb
zI1wK2ILC66/IAvImV5dXnzH2sF3ZFoOwiF9/7SzcIlGYces7g70OMfPyKldioWmgmxUQXIPh6O3
48F29QYAt6B61ipNNBoUQxUv/w+qdQLYsauLaG3KBkGtMiMR4GP71IlvqcJRPp3D4TI0JwnzccpU
Zb9T3wktL5dUR2AXvMKOJKbP76kGK159K891n0GqQfpSDWBqqS7hSwUZMQT1U3gniyCbNkuT9lTH
LJ4WwtncAgiRl1LL1OpFDNR0kBASuz+aRKvvEsDZ9hU6u41YU3mrHcMUbd/MQchMqNZKVBa2EHfN
ecTXHriiRTSD/jtsm8QYo9+rbUkkNJEWlaul8mEHSoWLgX9e5xi5OldZhwzvDQUSfJ3B2v+S3kzk
h7m2XpmgoMf5mxoUh6KOHy7MEqgOxCbLcLrm3rWRDuRPvotQO41XQAmVklGoWUqCotma+VCr6uHQ
vWZK68ZNmUmi8XGg82rwX1XxnHKaaS+bAUUVSH3J6b5TRuXxys25ihj2752qPycCDb3gYpJGjaaT
jsHbeDkhviZVHYKtNdCUnpz8tVJeNj+oMzm93/u9Mc1Puh3GzzrrhzxW9LOdwp50syGC9rb0LJwk
3b+uo7PTBe0w0l9JPmZIk69GixNbLaKl45xxPEE77Tdf3LXynah/RHavM1ZRpxcFwFO4qNVrjwsT
DD58nRe3jrQnPj8+Xk+68C81pRxc81Abz5zKCc7stDl/FzEr3Fu1GtAV/O3amWSPQ6RPLKSoTubu
9NUI8S7cu6kvQcdI6T7AEZXFe3yL3FSBSq6YySgOdAjM2en9Ker9azMniWbeuoGEd44yW/BOff7G
49Y28WSeB1VYBqg0X3CNdj8vABLI8Su5ET6r6kTVYh7BFi/akpQhObkgvH74WW5ScoBaLcJrLFrO
GeY/o0SkQ/as9tifdtZyKX4UPkBl2NtdNd3O5POGB2DpX0csF/yrnfxqK80ljtCVngKUe+uvCFZb
3K8CfKnD61hW4nFaVv6i7yefLNkltT2aBrE0FCT+r2cxDg67h0QDqzyTWJUoVHTQoqJMNt+ag6jq
zEq4JbEdqAGZtGL5MCJZtRbvGHjX650B/mHxqIi6TiT1dGn1uwQ8x6+Cs5Yn5xNpBLcriiuUBlUB
vgKxB2IoABN46UC3HsEzmEr1QO0u0lQ+hRf6OjGzUwlYBDjrwIqT4rSTfbTThEde12nnd1Oj1+FL
oo0fjc7QB48XbHp3q2v12PH7zIH3v9ZXW/PE87IYOVYs8QRXmENJTTKR9LhEMhfAsjVIIfQtgBd9
JZnCGfUbba/tC7L/BK4of3KNPe75fZpa8AIeK4ivY40zQatPOvrr3IyN2SSvCQGiBivFs6gozQ70
4HrTt7ZqiTQM3VyOYwj+8rb1jMHgS7zfaS664/VvSAMHy7CDfWQoSRQObQq1QeTvgJ6fokpUq+Yk
pVRjC/mfu2sL4oyVlf/Z0TlohepUSaIlQKFvfuACCJAYt4tc/E60YhWLGt0IFX4+j1pGmB+T/rnW
0gua3CL25VMP+Y74Wwe1gbYwOJORRbs6Tr3WWdridC45gWGbCWzC12xd55d6+SlfaRhglEMnAxNh
k1oHv65JpIjFLkTY3MXOj5SBns9HFCsqAOK7SjTXoKuMwh8tTqNQCEgMP8b5RZ+bacZSTkVHSCGC
kPQLBRMTMkgI+fuAzxBVUvYfs1hmVGH/Y0lRRsAE5c0r20e+3EXnyEf+eHkBSq1w4lZbG7SeapqU
ZYGAEuA2Bj4LRlGw5AZWZfhCKHhOUHerNHuL6fsMpEmrrZVnkFmwk+Ak2Ht8ddkWwY6n4OqJN59m
MysG9ekwDA70BChcJ+m26Hwxn1JS14EWymg6jL7VgUmqSp0fyEE9aXNuZFQXkH+3A5YJJS2nAe/f
B1WOLSXPosIOHNTTZ1nf+n6RPaFfArkGNaY0uRCdXldQNhZminx6+WdVj2zMKAitHX8/xqPLyYlp
pzV7j3j/fBx2pbO7oOBDIGpSFTDNPtRNmvd4MlMKPf/BprHvagP7fqrHaHijuwbwMMUff7CQrAxp
mV96AxIpiZ1eckgtQ3Y2gEr28zspJT9K8DXzpPhDazrTiWVSBhu3iVNwrt/Cnx1PuyS5tUgFNK0p
yJyIExIys6Gs6Ka16c2wDmEIw4misMKUdEEuPwGdFvnGVN2ZeXsPGX0T4EpkZ1m5gOaZtbMeud2z
svSlZ69ERbCFUOuOxhxfB5+K49MrIRMDgZAPjGE55GokptqA2DhYnJ78aJfyJIcfDazSMkZsFZGo
q7VUMouscuGo6H0wZ/NVUWo5ttMxr/Wp43vczpE3AIgX8F99dXEH7KtM3Pgxf5IxVd78wVZYvnll
IRjJxaK8fYoJ3MZhaDVPQ9w7GV0qE+qorY/otsGXJa9L27F2xawNM7HD4wJwXH0vm+gOMffj5/ZS
/S/COYJ6J8I3EGUjLfVqgj3VklfVc6V8sReNO0a/E8x3nyr3FmiGKo4ohZWBH2bw3ugvKcmcvwjK
AnkIEmaEMDfaBGiCCWKaKCpWEYz3DstN8Nlkw6KeIEk9qTEAQASYcqoqdviKpSlQ74Gb4gpyUP+w
LHVxQKgAw0bnBAWQugv05wLzyB3X2MJM/TLSG0ad3N8wkksQiovoewtrKsU7UN+6M9ACu5hJE+5G
ZRJL5zzxKyvzjS6avNnxt74eMW91hO+7e/Vbu6x6hsA1p2tt1kohK7dk547HA8GXrrXtUk7te9zP
NuWpCLTUfalG+LAV+cRLiJpqe51Y0NGQrBCK6anzIq2aCndXf6NfGdbvjV57NJNFFtAxv2YySNWu
78MdF2cdEsud1ECCKoZtaQsmgr1GA3cGuCmFWE5McNlydy6GVcxfwy4vf3Y6TRbR/QKrmEcURxMm
KPk7QOpLMee4kUm7Chx145zkhuFvPI0o0aFriSMRpRCSNrqbwOuzwXC32r7gvXchbyEfGHChy5e5
i7pwGAxDPpqBJc2z79x3vIlf5KpVaKAmRsiV4Q0s3SLLI+xAGzpFmDQ08ec+D/GJu/43gGZ4KzSv
Cdc11ye31Nk4B0jemnGyPRypXgCIMt9PuToVqEfCIAuVEs38I+n7fC046uNcqMEwLBnpEUE5XLBE
fNsOkx5mI8Yue8xVb1bF2dXNzpthPjWXzfckaWIHlxt8/URh718X9jbgI0xWEV7Y5KpLTFyjsAlG
n2UFDffZZmCyTPH1cfsVOjNgapVUWe7k6MlZN23CoUDtk6QDa9QtnxfpuxWfgmxS9Gd6Y6lvUqhN
HoA+No3Lln44xTr5g0/1wqMXmHr9NQIC9WX/gnd9z+F0EZvZpx5RQoqx7blgLpNUO9uSis+nPOq7
mnG9nhsFx6TxxbihQetRv7rBtz9t1QNj+ldiBWcBXyjw0f1erfDSl2Wd45fg3c7e7lTFzpoIhiXJ
O3mIhoKilUf5+oU5GfWHcUxTzVES8g5Hr3Az2jDW5rL7/nHNj8UN7C/YuiW6oqEdn2DbxTElHoYo
7YGA5UNcxRjThJlsP24p/zGEiHDsoiq6HefXySZS8zK+EPZamvPiLmiYaDEPxtwBfWM9LTgdMjN0
HYA1HBjGIWaJWxTTZDm54IPomIOnECm/PHuHRY8+kGODf4OvBiLI4dg69S/7fo0a069i7VSFaSwO
8231MFMfBJtGEsBLpv1DgfQQL0qUdrKc/j2oh6Qt5sSh++HaeWvOJjzGzLniw0uTGRnEoUGfQiba
zELQykhGjnyevxxwdmHpoin1HxVojyd7IQM4YR1m8s2FVwHY00YgMrgrPW4/oNbaXEwA79iIK+j+
LJX/Oj0E0Z6Yqjry7ahpxfxwhEu575ehIw4L27sEHn1O4zLRWfzZ3vTyUm4Vi/Lcd79nL7RGc7Ar
Bs0TU48TDiVoNufWWTZV+gdzmbWA/P0D7TH7R5ch784kMVzlod9Oa+lbURPz42+Q+NuX0iDbZu6U
EoUyUxX+20IQWcIws2qoejkyjBNDPcBRWE23F1P0GM6k2J+XHaWLC8Bi4cGyegpmYXNzDlpyBd53
p4e10BG5t/GI9wfHupH2cz5LZCUQL6qTduDjpiomxb7aSSekfwEjIkM3T+q7hKmV0FjiVgzT1tip
MwyMCKNkpGfJHAKpai6NdSL8+/d0MvVdzrjyPCPUJ0J+f77tC61WbGstsyqHb8yUoQPS0ibClO0t
jn/r8njCnFE/BgK8GUUiouy6bYWdNNGLIoHLqbX6phCh+gkeZQ7uJsb2XUaXd44NtpOKKo+ynHKT
oX1pAuSwjKx4YH460bKj7TVSbj9kfJm8n8lu9E808PBxssEItq13IcO/YCu97pkT7Hkq6TodJKQP
/AEmAhbN1rmRQW/R410B5a2JT6G7vU99l790gvtertlAYLH9m7hjM6O+Wyt4G56/GWgrSQq4f4ZJ
PnDqpueYg8oOM2CqI0UO+bUIQKGj5LOxYyRn9bkf2ZVvAgJZzFuPUkgBHrHAMbHpHHYmeT6+F7ov
eojRSFpxzzZuwlnoSGduFbKIFjZSJs9dVc5OuQDDFihvqBTBzrqT9J3yfGKEY+Ccxfzpjh6IfiQ3
C/wWXjOdnm9A0/NWGRHzZfYpOxUBlGQZ7iLVsn+dZZuxCt5w5ex43LJx9uu1S1vxAB7Rfwr3qBJi
IWtZAG7rcrGS0NtgIaqHjWhgubuBVthZxM0E+4aNx4WOSf7yndRwf481pWu06iz2J801WMFELZHT
H8t2wfGzl8doefdl+8pCIl311YhCa0HKeo6tkCVQQG8hUjrARtw33WRET/MwSV+9G9BPorvqeK+h
ym4q28DCvw0LmwFKb+1nqgkPvpXHFEyLI0Kpaicth2+IjBPdpFKT0kJe7CoFI0shI6BMrEnO4m8z
w4+KTDyb0poXZkRn3O9zrGHDiKIv2mPf6/xfBgcMDl65QBEhCHCYFPJli9ad7FRKJ28qkcDsMOE2
M7XW6az+zMzUD7X7Jjo4Ff1jYt+QR8BMmtgZlVUQUHbZLAHkltPkirj2Ime5XQUjMWLaDM5EJnQe
a0Jod4G/SZGYNMNitBKEAtrFSee08snXZmXjEnpHF/pLUVdBpWgqpq/meaiYsWKRAqqLHxxrd8Zz
5RzlIkyoBuNoWCn9lqQSdo+yotg0MH3vleHaftXfLqp0s3smtuy25Uvwfsi7eSmINTahFIOiZ+Uh
Rc4XQ+DvX7mpY848gvt2RYJejEIVk3gRfTyBB6dAzVntK0bVxs4t2sX1QdZKQYdRYo0x+aieBXuv
exFuwi7Ns+YdJqnm52fXCxO+x7QIH5Ez7N42NTmxZHtYTb4LFKXYDAOZpAI1liLqof+g+Dv04Ner
J/2HEreHvofiE2B3AVwtYbaUNK6StpwZ4DUYUlMVqLEz7bOxKZCMEIVo5ao2wwlAoJCV1rb2NCX4
Qpo9IldqBnhdQjofvZnqBb/FDUZIJ5XOFqP2LCou/HqVf+j9hoZmSmUhy3cLCixAIs8os0+Eg5/j
nY6iCa5ON2x8HAezymw0+eiIq8wmQJ6BBNstJfMCiA0KWZelFAI38s65Zll1Ms3CXLCzN+QkS3sr
rSKDAk4SmuU0hlYG98MzeRAtZDn3x+Bm6ym8o4+EqNMrt6qdrBnLOjEKweDZvfwj+oAo0iDYQ4Vv
4VjX4nUX1zWM9kVZTiubReQUQxDO2oiUUMgnToT5uX+WarQyTecTIjTo5BIjF6vxXnYwm93Yf1Xt
W+gmFpYp1joXcqnOcGpbFuKQAjBjZlGc+EuDuANTHFD4oJNPL7nRwUnSuS22TuBOz40j1CDNb2e+
i4rJdXMKyxVMJ9msKFwIxhsOYX6SVtP+SAw4b4Qec90g5epUT+LrQwPXD0lb5d3yTxaXcLjGx49X
owy3EBbRl8udi7MjxIm26QwZWKv0Ou37PUHLoC5UjKF0GW1uFlakGzz15DBFnKMQpLxf2FUICzsl
a4Oka0iNSRD6fW5x/gXF+umYc5yc1lDaJXakSWX7RJg4XaZImxsS7BS2G1uz/A34PBPEACGkYtDD
1W2zDpgy8btcClo6Qt/fp7ywmtYhVSWE0MwFnPY8xqCtjtsNqdx/9igLV5XtiHijhZ8N2qtA/EL5
r/VP/MGsalDC1Y7sdQ0uwkDhAao78U6/2GV7ZHIQpYa7un2+wKWHDAGUxvTnuRQLKQsTHtYyTBdz
zsDidZ2P9fTUrsAY9tkT7avcy+cPYmlkVT9Zji0G/Psnlx0sTanq452wJly/64HYxvC7+cSulDKa
gnL3Adr3U7gMcsP5jFIr08xRlh4ts0FVfPR9bMDXLl7HJcFt5Prs/ombWo8I8tX5wnHfp2ovguio
Af0E9t35GkTNQh2UoITWAwFieS4Im6tYMY6j00IE3+v4MX7DNzsK0Jy+xahG+6/SMYkeD5CNpmIu
n3IdDXBHnz5FMEDHFsORifPbOY3TDIa5LYNp3SKLKs3Rgbz1/ZyJsP4H7YCBicmp0nuNEOjRWKA6
DkX1L06JtsGIiSI/OxaH/E3JkPqShutFTYJeOPnYaIL1oSDnRXAkSMzqeHF9DzU4GPZudcBCitvp
WCbffhw7N1L5uGLwc6wEtC8go1/cG6NjjqlfJkEhC8gHYCvBse90PA+LcC/YKIaKOGXVNuYZRSF/
NnoPWMqQLtVigGSHdXBSOJ49zNSvA6n3zSDKr6gAxFj5ueuq0KjX7UigMZQk12RNfBhwslkC3BoL
3WFgTyWsTOVptYRpyINesSieTfQrHYvyXjObNn+LgVsZjLn6EJV46ydhcsG5iZDfJYtKXW6YQOF+
BkaBX/JXDSydewDTruujAxBfXWCzKTFawgXi7+tq/iVcgWj9ZlQx9bqMdJv9iMoAyt5kgVkHy0MK
Sf0+wMFcfeZOCPWEUGx1rnhciLubLfnz953mNdYFzr5d7r5CEkC7wgYiQAix8yCfmF/YF6FEGLJ7
2bA6N+AhtHjJbgIHmfI1UuX87I2DYdmY2ENrROmLSVcazPAOVK6KE6aIoxQ5aWWimvufHIOTpACH
6WQE+uSWpHKwwsw5fXdfKVZTu21Zf0fbg+txewiupTSZOXUIYDMTKS60gnLgr3LHYl0Q2nUjYYDy
3sH2vt3zjDK0L9iMy5UBV5otkx6cv9pD2coYh9jDkIwl3xM3NXI9liWvU43SP3L9REWu3ruGD1hj
hgBKUmltwhJpRmjIKmhz9CJ704uR3SOVu8hiw8IQH38cZJYUX9bOQS+1S+34gIBFetedOVQFjXXf
jGINzhInPVdvt24foXdLTyh1i2rWZcvsSPMCh/SbVDD+YW+62Gf9v2ANwn8+FY6dRP1uy8Ktb9/a
BN/4Jxk8rrCn7yhOcJOBo5Z2W3a68SCUFHsIBExuBkTaV3qK8BHX6taAQcDjvbwpiJ6/PGIzoK9Y
WlYg3LQztBmr/mm0sBYwM4yP61EsWmXJ5dfOm5F6JqSYM6DJq6KRjHHAJxptO1BiwzcB5XDG6eAv
M3NJMygBOCCTeCR7lWzutDh46JdnmWSyeOrGSEzW31gk/fr1otA0rYys9dfXwAfjKsEygO8vwrCK
b7nhYLyV+akKTe1LNSbdRziSC1oSwd7LvdzmRawO5AypTWVn9kKEsISQD2kqc1ccjtV9iE83tkB1
Gby4arS/FpqksDoLNtZr7uK4M2sKaTKOBKeuNUlhpzIm/1t8dCX1RlVRgUBhyQn9iAch5xkEUYWd
jDh5LbsED8O17GsMo+AsDLbvYi1lYJhA1ZP2rcqhEzjXsnkcAYF1/NJnMx1e12/AY33GTcupgBny
eKUvaIyObCEy4xearUJ//dKu+VG7TvnJeFg6i9+JXGhqPgh1crm0m+t/+KOBlcJRNAMQ/in3Rk8T
msgCWfdGYNH5N/wkBCCR0nX1KTjMfvYv50Qhgj+1mC0krDJJxgf7cjAG/0pbHOCt1T2aYhl1R7b7
Uv4fHd6br+hLdN9/z6h4tMjWzuX1knc4U4udM12d+cUpcHKyYySRD5On1O4/je014FC5q98SDPTv
bqi2HTLXE6KkrkicekNplvm/+jn90ZjsHUdF5nIlV+bJew0J65xf63CNAvicimQkl5kS8NYD1y4j
AGfqaHzh0XtON8xQ73itisVBlh3M+xWJinV+eqzzh9veA9zsnLdPZICSU7jJamf+b0yScCAAZaV9
D0N8ahpJ7bOv9gw03LuYe8UCTXoTYqtpEIxg3/yBruGexxNU4jmq6H6cure2jV/BNCNPJoz+GeJ7
148uWfMXwmlsSG4qlg8fJHMRrguRcNLC5sBbI/+SF900hOsgHroOoLNWpFCb8y6c1c37yEaq96/s
gI0V6J2h3c+0uSv9uFb9m4kuFYtOoNlXk1qplX/fh2tZNrQrIKdvUm7WrELdxgjIjLyx4O736+vY
8s1QGRtBsxVIkRcxxumthl7LTuS8HGsVuu5xHHEKEzPh7Hq6T9WZxZMQVe3ngzkjgIOnthkKvqa/
c5ejlRhGdZ/EvhybkklRKoKQCpzpCeELxuZu/K4hk+spNrTt5xbsW3HdDqpAulw2cWXUnn8QGnxc
N/q2UTo2oaJaMgCRjzjbyQiBDzx5MDQpUZdSpWn3Hv7SVs/Z9zdbsvk0D2VGuJq3jhllsqpLKrKt
2FrUhh2dPb77OhJ8IcizJlmtgQBb93mC9Pz8UfdkxlfetkVvjOWV7tVEks2NwY20g4gDSYZm/iec
2szLIOhYPoXDPEA2mbBmUt9D1NnY/RETHcsgq07A/5HBUjEp2OvfhUXJL+hxHan0UEjqyMv09A+G
l4y0NeVhfqlwDg+Vq6MdIFTSbYfNayzI4OKnaYEIorAL7eWALzxJGkYFAt+Mu214Gi7GBQuIpXP2
P/5ufy95bb9vx9npkzNf9yHWm0Mi/czKkVEpFY9xoT+pK90xVgY0IBb02RPH8qHQZUQIqpHoyIiF
Z43654QnrPMV/dEjs3sMZcwK36zc+JxtDtcnv9Ix9FsOmvVCpqA0faJ4WI7wSzCAxb+1PRmLpYcc
rhy8mqMKH/nbFd+sXHct1WmT/SpYU3N4Tky/9W65pE/0ALUzsJ047HNK/m1VBZ/0cvFnxA8okRvL
POmuhiUzyumM8Py0BFz0KYOC29e8LDKjZwZks7kyTZ8O7yRV+j6Tp2SAoRH4SN7iQJ9nMpc6oED+
L6C6L6dMpMqNjKEs2JDIgT+jwc7y4Er4gCGfAUddIMwgUXDB+xMzAyJtG2XP9PNsarruJ3qsZlbv
AVYqR4m/vhy/KF236MqKno13zvKQJsV//CG8TznqSGOAglPOmwmFYtSyIGgX1z9qlmwiJMM1g8b2
tM02Y+S2SipFivceLu978TEBqI14ggPNGfa4R0iJJdv/XIa2mjpCBTKnF4FEDfLIs7/KYNetOovY
MwWU+E9CFiVMpf6SVtsqE6XCdsIs6/l1kT7TYkfl3Y1QcAParaLhSGynN7y7JrUHw8tnEFqaNOwx
pE7McOLpeSPqSC9dpGXcPwn//Qq953WNH3+SyAGZXFK75XZwy9cxRavjzHeNFhs3ZvEJcmKWoX6p
VfwVnQ4gofZbyl4cnUTH3QCi2KAXr+vfC9HomPigWUO3zkWz9782BmSp5bwvEJptMweq31qx7/sI
RTEHXoqmO/Kb+OZRg4xlc4F8LmSXjipJhKBXpJIIFuo22f09OPPphjqwV2EZjAIzsjDFeTyIWtYI
QZT3rJUsJfBdPWYtE9PTIFTYtbi88zrPHXSzUjPCH4N2GOZfdHf42cBiuj2Eha9lsan3sbbg7AVc
YAkIK3Js9dK4Pyuljj4jszwWMFc8j7HSWfBpO79QDfsi/qSDofReI1P/rtymNxuH/Tj6HigJ2Ee0
k9+CBR466V0rR7iFBtLt7rYlGi+nbLtVPZtDzFoDq1ngn2jYxCeEq7VOCuCAtm3Ctndx+kLqhm5+
x/eeVQyslvWLfVeCCTyM3uE3/+vtADm3GCW0MIVxeT/IQqYRPlghIlgco0VXAEDIUoFwJRWq9uAR
OYg2luoLnUaqL851RhXWU/WhOH+CJJ7exIgCf+7tD0zspBg3MahH9sWVF+wnPuzE6qY2zt7MhmXm
9mM1ENWFbVjHzr7Dkg/eDd9JbKTPBnLxoIwBjsVQzYgHjXAWTBsbrb9KUyh27tqsi7qL/sNb/4LL
ibhls7WJBgPzDqpAg0kEhGV+RHEqPRWWLn8eiK08fvSNmHbEM1WnF7ix8zPLMU6mgeq1zUXKAAnt
2BhMNTgYujBxb7yJdg9+V7NiBL7recyCyzIKP4g7Zxmp2NFIqj2pkjInVzhZgjAefwEhH7coTHnz
7avVGw7TDtQZC4HlLRtk/OEwBc4yOLGZ/8nNXppilXJrPlKqg3TgNQd2WB9rQaSmN1tHNz8J8INl
aEMSG/fWtbhJ1CUUYU3HL9BTm0FPTS/oHD8SlE6v/ujBrmG5+QZv0a1RlrJ1Bux0lv70yr+Gu1u1
bUhdo5C9AUBpE8e8rFT9WDQCLICjoPbAlmIxPg0ah8UfLIBS9pV5U5tyT66Ov11k8JXcl+VgZhlo
b+brkBTsBnR9RYWNNTlFqE+jCA4/ZquNYB8L+50W+5MsvWkqgIRzBNY9YwtZvV4HfGsgtklLXx27
oGOKLbU2la8Q1HabS4/o77ErHTtMgiwz7g9YaYjS8/J+vwATPaJ7/V/mhFPN8hXYpkyf+VOQJGnr
++0Redk2Sv+8PCH/M3zr1oYWp+j0FK8ihFsUqeld7PHfr1ikgLwKFAIyVmxE3QKUCntt9q6FYc/L
e2c0r4RyxD8FfjlQrG+uLIm6vBolqCuJ9TK8142Z6A0xOG4sDRkS3k9gj2iVWIj0GmaOzkCWB8Gt
sYrAtH9o1SGzFgDKnBYSGNdGO/WzQ9Pw4gwQWEeAINWzK0FBOihFikzpFsCXqEdm852KJGPyhlgx
EoE1AMCh39JHiI1Wdj8tkU4LmNYa9WNOKSCpk6h9nnPMVeRJIQJL9gdXXjWSuGedD0JraLxncAep
E5FgkNSxdsdKJ7jaBeSZEO2JIyz1+waa9ExaXU6A+714zXMEtsI/BWkfSgwh54SKcvq+OsSmRvZj
xaAzKsyHS3xpK2oGiy+nQiwOy55mAZq+H9HHppaWFx7XZFzFMK96arceSGB+dc6NgsrpnN0rfwgA
Qq2MGBy4pGpj/rk1fHjwxdSvWAytugWBMPpAjw77w2AbpmhFIQCfIfQ8qA2KvypJ+1HMnlblRZ9V
fND4iVPBiA1urKunxikKbxD8VdZddkiRqxwRAY0rvYEsuoG9vsIt9LzklM42w8/a8RgCij67rBmE
UKsiPYo4IVINq4lfS7OrssiMlR83xMDAsnRZaYs13LU3mKghwMTKW+QVwizVhjzx6MNgQ3YX3dkF
HakiaS+chAf0JVlLSMYSfxZO5vYdnJnCZPquJ1gPOn4WyBCitfEpyu6R4yDTOo6/z3jMpa39rWkB
YXcVUxHLBJFvAt/lNbGW6n56sq9N8bNA05yPLLz18uBc4H2+1cMSFqC3SsUsyaX6HpKdJRLdNs1Z
yqGlU0R8lsxRBZQlweqgQ/UBORxQwDSM9aqvgKaL9NDiN8leb0slYrthLRbaPpPoK3j2sof3x4UK
A7z4OrxDpe5jko8wNtHevwwsEa9lSgT+sjizF6mEMbcs5p/xLWPv48/WnriR2ydVRc7LtMet5bxf
61pqNkILW1lEOtD+hBm7rIAdede3kZx7yjJqQy+kvf82pzuikE0ZnIZvZr/8LpxdcXEe9TymM88s
vcgMJQBE8r+7su8pcAeIZUZ79cObXKXCc6042nPWIbqNnVmPpeIur85kAbKQRHd2ww+aIv0q2gZy
iloLLT1SZ11hmau2Zp5ANf6g+NwnhhBnsfeCYLpxW4erFct9miFmG93qC8sHRAUztbU7LlvnjsWA
hPuux4V5cZcbxNoLTh9Xcu0tduq2bMzrZ69b9NGYtvbFMyU+t2XYrAqbQxMQy3T+id+ohWf5uCUS
BLP3pmWcw5/ysLFuLaUl4c0F51l0BjY0+fxijBPXH+QhTHDayCkMWEZG8ithY3KWo7SYOX/7st5k
YD2uCmlhQ0nLp2qWEsNjBjuWf5gZRt3lAJ69mFLlW+Ypwyx3go2IzPe2GmJPX3oWRCLGWrRoTbWX
C0W/bcCKYRmDiFT01+ED7XhhZffqeUp/Yi5YTLunYvDp0hxlvrb/t+MS3pFkijDRic4Phvmi7q1N
BtnQnKUZx83+Xdhxv8fJXWunMz6/fLPsB++7UYIN/XuKJNIu9qUQAxQpqCVvEPLlE+FK+W69o3k7
tYC/K1GcgL9pFJ+fOTLiSlWc7bPG0E6k3T2VlX9piZGtgD3bOKjII2sExsGcSCyY2upQKgHpnvhV
nu2Y+n5EyAoGPVOb8BBlx394iXAcvkCXRYj9TEP/vv5z4lD8AHTUmnY8bLIbIKxKk1cGMudlxCBK
0JNorOe2ehYgFrPyLNTACzvI5DsDXp3FajujNCURp0qDnxIo9kmJD0u8oWAnBnVjBWt8A0CEzZI0
/udg2RmaNh7NBEjOJuNcY9aBEFLE9ZTWS+Uf1EqoP6kluSoRnZZotzDYnxoW0tLWgCwhdC5uJix1
8Gsr7z4uhaWJMgfzam81XnHzZmX8d6fuVS2LSLYs6zYY3+vfdLxGKktbCEFuJJ3Scd9T/VixiUKD
rNo5105NRNf6k4mtM/RAcvhLuWHliU4bvlrbfCAeeNII6eo0NnfykbLgcHzMJzYQv6jKcz0rdB8B
2gprloJZsfCYnaqkANTUSMC0CiBEONc0cSkc95NpSmO/rdGp2WVZiOdI5qjSo7Gka2LWQaZaDLmR
NRqkKym2QN4vbkkpgR4Pu3YZwynqibCBWGudoenUnYrtMa0TfKnhvE2Rq0ibTuGavCjQjEYsl1FE
Oda+0xHkxNnU+kHhc1k7+DRhSVlmlDGsHMZqPAfG5b9cYWTCYIZPmOT53/hkACzdzPD3R83N9NOY
AFRyAWzf6dZgzOZBkEw9S5iGpVZRZK1OKDca302/OegsIpF5SOx/luHNoo+JhciIr1H4q9KX7XOR
OO7Aaxem6mazZizFm+5UbWP0KyWgwDE+HdYpgsGe3FwHeqB5ChA325fCC914T9QjGfeycFl8Iccl
wLho2Uu/HD8FMKmsd0ywuiuZxfrovD/WhDqYuANzvJdQ9QnuwqOII53/wsfttl3VxEui9vomiga3
umb23MIPLVsDYJYqud1wDfPI5lZF7xgC7bjl1NlrFa1TYgVakPIGLngSGKxe2Co0rTNT6XfDZX14
LV9j7e2ZpcV4GO1jOR5b6a80p7gyEzmSQ/Ah48ZGt+n4TkJZrGldIxIPJhYg2KxIdHyjKPySY+Rt
7Rc8fIl0eFGv8qSuEf6p9VJU+LSbjF9+KhdUw7sZd2y5xwrX3L/vD89YjcCIHf+VMNNIxPOF8eqO
SNLyPpRP1affvB7wt3w8gUs1zgqIFvDAs74qOlDsfmzxdgwnfjMQcbySn6go88VgifRyi+fxUdz7
Uv07frgm55JZylPiS4joydYqVIsj/mVg4Woxg6nMZ76qJAWZu+m82lUHiEqqRXE0ooFxwKT9JfXp
6AJJRevWqYN+MQcqI4Bj0gG3uglzPHmTIT2DcZqAJXFoN5ZcGa2mrHtrHPAvjgfI/+9G4g7Gxk6p
bC/Elvp6RhoEI3PjI6KScxM7s4JjDCKL0T/FynbsJ+r2f/xceEXFPzmpmOeU7VjHPLaxAMNj2089
PB0xXUZ41V6U5aOHOR2NfD/aCGYDQqvj2brJbIv8m4Sp6hxhkqp7luAaHuwJv74ot5W2GOEgnfNp
fWSm44xDxvWSEmmxcJ1zqTKFg/P/DnMKobdCyQBxkBL6RJBQOYV51Kf5pXI4+Tx+uj9+rbs9Cerd
Y4jO2QC4Vd0y3q2F+WJzShDao7AIto3R2YHGUzA4wcLKaPhMuSAJjNPDqpw7qyUrMtpgit76Ai55
JVMAMVVrWgcYMnGhzVirlODgf/ENbrwDfInS/iF6qQ/6wG1Roz1Ghgjogh+H5EFSJWWPAOu0rGw+
YSDpjuROLv7KnoDhALrG9hfP5gFeqxspGmYair2IOqn4Oisy1xOTsf6CxAATf1InW0F3JrUNisTV
NN2zEwuyRlO1ZRyHbgWYRPl0VphSWem5PrDCKWieDXnko6w4bTFSmNyXU4FbVhEwQr78soug+J47
jTc63Qu5GquVkztx36tHkKa/mT2ND5hLtY8bdl1JxTXYQy3VPqoyHHomwzUUlBbjhlg3Q8WTAjsW
e/rLutskv96Ckl1YIWbtkwpmFQCceGn74/3/hOOlh/DunmxdA/OFrebXUSNnWrFiHLgUezcCqjMJ
gm7rgFQMzszg5JtBWN6Bk/mP3KlmMPnVqFMedPuXI1EiXG7QH/6Wntjqo9MWqiXGSeN0651slC/y
nbiKdgRcDls5v8ky+GWiM58o1E/hQ4nzLWfQl1GkIAVf7VapZf7+94JsdDYguw3KCe0IDHYPAs1U
wxWxm6cmkajyV2zftxIexEIhLpQxG89fzymu1Muf0kCZgtzsCDnOi4YZe388USQaIqklM3tRI/nC
AE7v1ZS7Ey7H71yWCFPPTyws0DrHFan1fLa3GOdEbD8VZpL2bPFVByl8dzyZJcHdv4boOMDabPrR
7Ef7kC+fY+MBNtdCo38gBAWlFTjeIbPjtZvio7D3m+f5gyWMsh0NMIBTB0uj3NnncNH7W1L4tZQz
S/3yXlz2BMXycerZPa00pnpV7pdrzmfhckfDgveW9Xfhsq2UTMx8Rymt31SfdXzt82KdKeecRY15
x/f9Q6IQgffbgLY+WeE0T4GJk22X/B2vrMw0c5ME+1xsukkf63eNImq3fK09LYCEhXTqWhVVkisK
T7xSkNoxvhO7iysXWnthbImRijn4g5xUWZMPIBM+ISJJg8tuJgiw/o2mVAJRQBhACMhaFsvEcF+6
JlqQVmzJd0qp4EgAR91SluaeY+2THM29hMILeS/Vu59Ilhry47sotbIv5hz7trtth40dwOkI8hrb
gECNakEYkp8+A38vFH54PNH5CfxfLs+ItKs9jASeB+7W2e4xoRhLLGr17TIJTez5YceT3xRrEWxg
0T5dIpvcZFx7dXVMeF3gtKjDsAMddioE1OglGe7Y9N0M52xsQEvNJQ6qycjm178XukXIQU3aCoRh
fTynC/jIBKlKjDUe2MQiYgIjA0HOh4Gha9rblw6seNvAcQszZG6Hv4HK2EfBCWO/P8lyB2TzX3P4
xg0dybbAt3kMuozMUxlAMl3bg50cAnnagn14T8LVHapcZBnONNeu9E+sQl5jpI5HmxbKjOTv8WZw
HheYTKbEj9tok9RPXvlvQwLMcWQMXrJ6e8/c94iVJPuNwjwd7ZlrGDD+bnlrMhTk3joREk0i6HOq
B44CbYAy0uMmlWJlyta10DNeoYsPSoWpua5I1TK4CjOtjFTv08ID/Z9SF+nsvOCV8SYfZXnzSGlf
dqnqjcZ+X5F+/DVztuuQJ1MdEVZoCu3U3tr4efmTQgK3BrH+FnYBY0sqmGDNmQGPrTBR6dkofwoD
Y65yX3s1Jny/QOTptNQHIIvALjsCtAnOeK9rn9dUZRvySCocSquoaIkerofhRJPCeyTBVFoVDszZ
ubqvxMAoJVCQpIT++rnrUN/tpzUZilHE2Pz8UrlAKqVgjzFpMBcfHgBuW/FgJDGsfd5fnqrNzug/
iMA9RtKgenJEpIsq9MUlZZTAmviCNWdrYkyA3Hn6r8hILUvgaPxMmP3bkh4gveSBor80YfV3AKHH
MTU/RmFNUyz7QfaL9Q2B6P/L2ESzEo9q5LxjOp0NmRQlKDdyAJucYTFbtenv2o8qYQDKTVdtMwFZ
7U/gJb2mpSGRZhS9Ncfm5EnPRaWXmQn1h11PaOBlDgyyX6Vr3pjc5iwsAGyzSJZxul69w4BP/6uI
7zriVELthnoSH0cchtL3IxiYA1fZhaCj3/ZhAFTQFTIUtlHMEbOuk1Ra5JnE9OToBYuxjp6+kw/v
xUtnzOdtbfqkjTV1caBNlc1vh/M8bfll04JbeCTp/hYa4MNep0apghN90RA7j6fhHYn8k/Kpay+p
arHmPQOjVrgCW6GtzGvjLf1194q5wOixLoPkhgazXj1Bkv85CZhssEIJBLXS/FO3YP85WbmqSvTH
/fepDDUf8fbtkWP+Rcv+Qw1F50yv+WxM7EAaiTCwKeSCZFc5U4TjyzG6UJaKYZB7wz4nkT2gfvBp
yNYE864LZ/xeLCesh2Mrd/MET4DYBgyKfaJQEuWZ6iRygf+UTyYw10zHKz3idum3Ge5hFxNsPNqN
4mmxRxgFEJYKkaUT92fsvjHMXltZpeezjnvHo7wAmLuwv75YR6vHw7BkjW9EFyDc/OOkQeEv4s94
pnWUgtmRUobH8C4+frpdamRfV5UEyyPrlkuIf5uxvTqV7TJY7eG4zKtidX7CUdej6Hdlc//mqY0C
EhsCA7d86GjXLmqDSPbEC4nvwGC/Nkhi/I7fYtQ49YpGD2WaIUQw599skCpFYVRVD3Emo+kAYdIo
mtu7FkZFxib+8JRd8bGlXB5sZpeTz8ItQTB50Di/0W9qZCPTtJuxcEyH978ztMra1GpSiChguLHf
N7GHObSXdXSn2k4EoMnHqJHGccZgc+pHDEsc5ibm6SE6cqBmr38UbJTk8MEXdL//lDgtuG9oSgmb
BHRaiTEUvQ9EQPIG7XqheZJ7mTpY1QkbFIebmCJweKUBiXgfdp/AAiWs59qno7dE/qYoPIc9TO37
nKn2tUSvqjx44qi+w33zNwbctwq6viEswY/l/H278f/ZWr69Et6hf45c7V4iIyQIc/P2FjM7lEmG
qEZdy/ncZdCE/yYVrODVeDlVCqbvPeRIRogrKf6gLZ+dT1EnnE8GYu1p5K7xlW4qMAP2ewC5LPXW
N0x5lEzqIZYMc/XLmtk2u+cwE5FiNTr87q7A8ULBklQ4os2RTsXyIjhfgA5+B7uCJwv6GfePwa5a
IhRO0Xl6FTfzQgPDeOXfekHErFwH6lxRhetCD27e+yEYFNX7zIrfGnLd6nKW9hKismYuM8rAnHRy
LpVeQpKUuvQ74lXsXGKJKjJySLCKMKDYbjguzjT5U7J2bgjPpE4RDM+qtR0URAI0p7xtdUPovxni
VIMo7EKajHqCTR1cqzmoP2vDVchIzXXnga2NhcOIlCE3XNc/kOxb8a4XgfmFeFfYtwtHppsYhuVN
lQnrqd4hQ4Dd8QWiAH15GRa9W6Pi7V06dkoJofHalsBU/ax/VUiuJpbg62Vbr4SiNPj1Mco7McNK
nXwx7uw4Or3ohMLISGiezgaDPP5EcOKYpKRVyPcsUDn5dMSUrtMVWJ9RN1vxQJF/1jMUtNS3lfQe
dFEmID3TVOQgaDV13EneCIUPVDcco2xcrx3+QA7s3Yzz1zboyAUGl5nKJJVnE4+2Q3uCRvEOlbtm
5qoO5uY4qpMDKwEh0gOCuMraTZ95h1KRuALSQImlI7YsSwGUDqros1uluf66z2YbmxyGWb6s4nh8
jhgbJ1CsCUf7rSY4qSUr5ujNI2KSwXR4hHDgwtrEVpvIMW9M1uLM9axnIAziFgT0PKbTVwoyghFt
Fea8GDy975dwdwwkdIhGJYvNfCAMbQlEI+mIIOFG1U8se4NL0PVEZcqV/ryJipnKFPLJY4ogIM6c
MFu+0NLrIgMbuD2PlfPnr7GGW++9MxBZG8ganT9XdxMBpvFeLsJlWoUvrvbwWb1NCDa1Rb53D3tg
b19Imp3Uf5U+xiY9hZGtJV+FOpaEzNMUnS8ieN2ls1ltUavfSL3+R/qaTdu/N+dN8OIeA+m9/Fmo
RFKWus4xLFJJtwsxgdxmL6JFZ6IMrW5eUVvZICkgEBGFPNFoFDNWdQCOlpN19bCwALhoyiZpGylU
x+jXz7xRUIMi/ZEKK0v2NtzculynOmqOMyVNcuqhPOQfCyn6ccx8wiK5rHvhBwl/v05RwBicKuWL
nAMAoBRqPr64YHxslLJYHRp+u/NmL5JW2s8OWyMoxAZbIaohCk5pPe7vhbuNPSNdsWjDw8NmDlgV
QPFwEBP/qLnJmhWjjKK7X7dR8wOTwcqLSm8U49AJ6ScSQY8R9AbBS5lwL6ASJRB2fEhDn9/DgNYx
r69VRJmqE6n98+9XwbA/MoSrXyYuJ8vwfwBeg4fEDVL/EL4Jvl3kS39Nus3Aq3xs5TYvqmq+MLmy
gU5/d/bMFldnRyU3Imet2VWi22Qr4jjq89ZzwBIEVX+IEgtJ6/5nHX8sQrD5WteR4BioZ0uafLI4
XsAG0hGQLHidNYwRiEkxAAMiwulfqLDYFvbVobj6prWdzzc+ZPzjY2P2tRBkdzcZXIMm/oP5pC7p
84Peza3z1aZDhVWBK4nTXI7EkR/xwVwGwKo4xPVwexv+c5GQe9EqIeccS8Zpp8dEGYNSVvnVwDHq
8BCCGlfDyqDuTNdxfpkdJVdTnVU0muBxszVZ8uV/j6m5ZAZleJYE8nfEgAP1fm6YmynV8wYFafiS
eJPR5fYtYujY0rxozMxbd2OkLuS1t+Buy9/JwkIissg8mOyQNufLPvOtNxX2ynSPFYC2Ld5LpmHn
cD21z75+KFotVlysS73bpGl2SWjmH0g6KveduuY33pTwF1TeA56feYmhPXD/abZIIYLy6+O+FzvF
s2tMHO7P3LuK/EOm3iNeVjXoWzDpRgWFUUAIhsXpU0lDijF4HGBOpNzXdBx6ncG6iYVgrR7wJ8Wj
IAHqA39cilAmPkW6POFqSMtC95KOjgf55g0rKptox4ejwO0gdJL18vI9Y2zumuiEu+xeVnXHxIOl
obPb/uFt/yy40G8gTzhXLOk3XxPy7lWwkyWMnO9SAGqOWzl1tzB6ROElI38Pd5vXSd4Z+nRFWWW5
Ipn0+F4XtVKVcYcQpoKPeznmWVutj3h0vzLPoktPa7sBCKMnGn76zH5D2TX9lWAObaKphJ4CZxPG
IvivQipu/+twhGrQaN5ihoRN0eNOcAjaVW5Zrylzh9MBAplpVrPDfYZYn5W9X8OChJgq1jHHkbEj
/JFO1/0ooajQEd35Z7VG9PJbuJukgVymIJK9T6WXMVYMBKb16w0AeCzVMYiJGMux/9X9dFRV80Yp
2LTb40scqbLGYFBQuZO6IYOGIuvvrpY5djdSDOq8EmHYdgK52d8H2SBTzSIefDoy7bpUF/O7Bd30
bGnmFBJABr7AqxDDn38KmNhU9uJG2SCvr8zdCN/EhthzHPw9lmp1qV9mjDlUNDI3OcroeUQxIHuJ
EyeqTkeJ61pbOlpfwRv5c5F8tAKQoauZMh+zGABVi5Y6ZJY7KTprVchYYA7ruK3/BpvabQ7Zr4ab
ZWpDUDPOJvNWJmS47GsRt8LjpCr0gfuMAOWSmPMETDXXmFKB8RYQg2SrlSji+PkL65PFYBg5L5jJ
DhvSybr8lwlrJ7Z3Ingn/UK5LJXwLqq9+m63LLl1gmKQo4EZoXxSx+7sfQsqDklOgqCZnWdkl9va
GXp86YHffqVj390V5K0bYe+UEBq8CUePohyuGpF1cEcR9ot6XLZuq85hz83aHbkeXGu1YvdrFDm7
p3/P4p1P72xVO2c6XmBOFZsAC1oZOGSHZb49f5yFwOAKnWG018uuEgJsCqVBrMd/00MjE1hEIzz5
O4+cplgnppIBuhb4xbxiRsiZmdd/3RIm6MnUhCba3u5Hq9nmN/8n2hU7AevY1EUESdFOvOi3CoxW
M/TDBYKBfMDuhuEV0oHiiixpC1aAHDN0V5d+ZOiq1uO6P6i2mZV70A8uOAo1cwJnIC3pC52Q4yQe
dFLoZCOpcUwDibdNWI4OQLpkfsFMB2q5p9LD8o3ymoUKp1bSCdBXjbiitS2IWD8Uhni3JKjml0wa
XOcOQIB7akOZt4gatTtZgfGQj3fcc52TDgq/U7U5X2QuCLK113R6GvUQZ26LKWVXnsbfchldL4q1
bBvsuaZ3GxLdVlTJy/r1EX/Fgc2geeujG/HfXg/UMeFL74yzZWHsQYJWQOnIy6Z59H84EE8hLcBw
5hMTYAmCyqIP/mPjBsyhFDrhG5rQaf8L8KbLzAjEU8wwCp/tWx8bv8u+YsEqUSSjXupXcFttRJyS
uMXY3SJpwRveXjdARXvjnaEgbnekImSxIj37Z4ggEAy+M7hJ8xavBNlAYOBSuaHJfW4A7PdRmPN+
4cQYzA/dV7EuAJ20uJnMGFH6iXCNJPXkluTV9z7/Ixj3bNI7ts2CcEVbtvcvOLn7WNNXjv8++1Ak
iRLvEeBmpiGRDkO0Ana0AC7Qxde3M5K9/ONDHyK5tAQxA+RibD/Ok61ni4TZGdM6n+qmYalKpX2Q
lPuuF6M+/X0K8wxuTw306tNgzsoYRURSmYPL+nRzyM8IEiFAgZZDpUrm5AausZAlXdimKC4CUmAL
N9Plgkh/Ab6NneXwaHemlRGF/4ezx2oO9nklS+61233nt2zecU9oJXz5EZHKnIFcwmzmuVKX9oCF
FTOfgkDl1LpLX7ANA5jx5ha2LPqErucpLK3tlfsBMdUGKIXmADMeJqljBY3r6oVdZrRDx837i+V1
R+/Ws0ZhcbMIgHjmjopRvTOH9KSkd6NUvioXUHWl00AIqw2o1z6Ic6fVDk88doCKluvNIMqBuAUm
79M6FnGlRbboKxIb0TI+cldlFKIw+pdB7j7ZZ1POSqK0iGAUCVKh+f3gKm0t4zRpFKda+g46QD40
dSkHN1ct6oD7xzeWH1z38Vu0rg5k5vBJptDDXYJucqg6xj4m3sMU4uldLZQECF2JBRQmvMscVJrA
v4HiScYTBS/ju5BfzolGgJbes01tHYZiaA6+xIMX+ROn1abVNDZQUt6kVzdtJwun6t1gWw5ZrzZ1
eU/W55vp1FD0qfypJHcO4yjqfDaZGiulBsnRf3lbbUGvh6uzrt0HX4UZS+djC8Ul/FoOccjx5WyL
WMzxy3FdobrCckGWz+5Tp+6hxn7VczkX0xJmC23MXElWQJdh5ZO0PC8Tb4QFnvzd97OO32dSoNoB
GgW1tKNglIvAVsO0aBfI/OIwwrOfs298HY0hel1hdulEOJ8tiSJJTjeMXkGfQxgcPo7imxknOGLm
hfFfxzxvoJTFJ4iocsHt98tUqDllIglI4Lo71WrxLz921Dmgcn+nqq1G7OMkh72froHchUjtfgZ9
p3rDeuGCmsCaTjsmJ9IZP3NkgBaIlniS+T5muwwiNr0K7UfhDvK1p9s/d5x/DY2xMu3cEROUF280
dYmLXQLWpIOgh7weAv+1cI5X0MCx8my7qBaL8n3iMkdYzhyRl4uTihkbh7kOtK3b/4Bk9cexlaeA
tz9FK1JfakgG4lNyGjmCYJl/5QhXtKIk9RLynvACYZPTokBLyhaig6cZNcDxs+9rxhE5H+XgLifr
XAuJztcwKHi6YqDMKXLwmIWnN2XJudxh7mURds3+GOfuiQYjQlZtScsGslCfotsi6KUBCUBKQODb
gjGyPrEz6bfz8bV8+NQDYXd7UqbJCRRSQJMSTl09nDfiPGXUgaOjyUHymqGcJQVAlo+aGd1J0wOj
P6SQ3OYBHIp3b1cvgKsSuZLPCq6NPwRs7U7DSwmQXasjB0MEan8yDTFeoOQ5VPF62Y8kunF96rrV
g1u3nMbrMVOLkvZI93zkF/mkSTe/Wr4T1H9k/HS5R+N7i/8s1UDQZivJIf7pfPa51S6kL8bw9NXj
aL4Iiq9v0Y2wszAGQvdQWTw0KwXqu3QiTW3Q22L7/cNI99UMWYb62ESZ9micGwKJXIDNq4639RYN
mErBmcP0Xq7zBwMzsn8A96vQ3rbfoGqj9sWgQf4t7SMgck1yxoDbCH6lJadC6QLu+d/Aq8At3qdH
9oW17kTW3dHKYLG3QnmQKYvh1MPqFGTFrt0pxOz/5erN5Qvz+qkK5U9GfR8iXu5pzrkyNpOao5Xd
LLKJpu0M0jHi3CI73pDOYuHTvcpmd3oShmvNRDimAj7yvOQtnXd3EgGMUQxsb4v0BUu8kCvWWS23
x/cHqaDQ+G7QqpqUmgm1S4kAlSHqoUCAu+AoG3zSRszZB/kNzYVLtRxPlyIgy1nnp5TH52pKSxyB
bt+gmSRG6b5DTfKJb5mP4qFSUu0y0sERK0Cez8/5nHVeCm8mT8+yCoZcf9d+2ekABUwiLHQqgTY2
IlYBWPTvdFoQElCIq+NeGEOhm5gsy3CudTBmfsQEk/mH5CbChd6YJX+7XaNnhlMo7NG+KPOQI1BE
YDwM/fWM9OneoLqQOWL/3sqpX+kg1yn6WiICQOQzqSIZ4l/fqrcCEDPSg1p896ItchMd2X54G3nX
QK7guoXJfnVLfh4yOSbWVNslU1XmLpwWrLCVgNWK+Tido3Wd6V28UwjApAp5td6FR0CI9byVSFlf
lIVIgkq6PMLhzCGEQwIIuYbVDwGkl7zv2PPyKKrikJoUcajQHGfORmIk3yEOZCxDvcbTFvrXVBGA
caJRKlnVve7MDk2VJ3qMw9mC9J8OB9RH1MJ8DqNRfvweMfQBFiA6dFF4ybawTdRwbFUPtsyXwIpi
XQAaE5ACycN1Udj0SVUX4Zu+gMTT79NoRxgMwNjHJ7NtB2jmNi9xWZBlS6j0HLLiHC0hL3lwosei
dCssU3/v5aOh+NXtj2rO2iuQPk3VKPjvcVruE8T09PLzF429F/gK7UQSFRl/76ZIM94sSuOPZhB+
Q8bxpoZ7KbfJu1PKSGiD1ZFEvWPTYi0PO56C/1wH2buFu4tVbR0m6KdQTrCvQLiEY7Wg03BKorRb
iTouPOGJhjVhJf14nxoN1KnyVcfhIKnxlsdGVYzG+VmGWRAh2cuPYCIsGS8ZGidizU9izgXEjjK5
mXedWlOZfJrTLKaw+6TCDBqP7o1nlpV1Y+DKrQJQNfEGmc0iBpm0UiwcQtziHg5IiftHVN6QJASs
Lz7xp/O+bkVxSutsyE7tHxI969kEwOTWmYO9uW5UEuuLyrn4gqRkPBTvvhiWrqmLCvhgExchNn9O
I33jOxsluHRsBFwNfXbqOfXl9IiENzfAku4QFHnWmISvnOYevayPwjXs4hXZwRfdPLsK8P3frEru
oWjPcyOMVlDc2CuwK0uje/cmwl3nM4jRAQtmpJq/igpXISwgT3jrLMlr0AE3xzfZJLDVOvo+qyIk
/RJ8t7iUpbk6Pfa6OoFtD2oeQllL50zU9QwoDYwJqVeR+CB6fqFZ2lniO/3R/0UyiVyzYlxX5HuL
oRoDM8ztgPo1ZeedHPPuQCeYqjq+V/c8WwLSx+mNd4ACj7regW7I53oMpAKJKzAtf9+2EIe17kPZ
b4e7za2nzIptwgiLTvC8q3LMtPnT7NrysIqnq/WcIxct1A+obNtwNV7lVcnprsR+06AnR8o/8YHJ
CIGOzFfDWTKb+xK9J8uXhN5m2eouP2WgAU8fswQKNv7RuHh1/PMmahBQ94Jgkurac/Pb2ccHg3Dl
KzdyiRGJGx5dURO1jtWnNXYf+c1ORhqMQM+pZtGnGIrTuEQL5lnCIJy44O9TSog/tKvVQqcUMHzB
gpeyweKEpfC4bBw0sAuivTbPRclWBmHBlR3w42NWQGdZm5pBjUbHM3yynUsTN4q6FW6iB64M/jKG
6uxpkJWAX0SoLmDnR6KYDdKN/c+nVltgQhDeasmwGS1TIrjTbUxrDmDuOn3Hn4NukeWW3JrfMwL3
f/G6Qb2sJztcm78Duy6dKFq18Rdhz3Wi0QX82/N8Q9/UC/j6allDMS7LLPm/0n8zlcafTCtJlQtp
TzGmPZ0wJ64dvyxGc0fAyFz/2usrAwEyCveEW3iSXydZM6G2TEMI38rEbxG8jEBYOqv5BQeOiCwu
wpg2mnyjbkenhvbDWubUeZOuow96lxBXQ8WAC03YUl5na8Fgoo26KPCsAuT97ss2TYSC1DG4zGo4
60fxBREyaKDMOGksbVQWDGH+uTE1K0wUyQDvAE3x9zFXb/YWNLTGKtfQfp+U42YmJKhbyb80JzH1
ohE40l/mk6N1DhNWTis2NYnmLhJRf/8t7B7tivvtozzfQFCJbQNZ+IzWP2W1l9UezjNVg3ny0E9L
UjccprVh77PfqpN4hZiMkfGNMragegGbaTdZf5HuGai3LtD055XEeKqX7kt83yF0uLtN0y/Gcg0B
PDv/pPC90RlArIPAX2z5G24ZPPEQ3sy6UqTuQs1YN5vdCA84g0rGjThVrrRwIfYOHMHBFnUe73UG
3YNvLLijp1NC19yHkf9VYaa5JGUMWJRZchLNr3PidtMWJKDRrjr8RYAG1b7y5EDg31pUfuWl0gFk
Gp8bG0iKgU8cbKRbnLQhYUf9rjR08Atz+/s9LnVRQz7xbu9mPTpmmJAHc2sZ2PqZs7FrNPGKczof
hu2AK2wRwmxRGdyQw1J/6bHnq0NYwURXwHCzPGnN9sNHwLTPnwngtx4SafxKmU+93xDcRPpIfRFL
lrofKJaFd8iYUR3Z6wYCK3diLRrWuYhSpDf9LRzyB1OyPG1/N0mCJoBGelaOvge2AWtXfW6Xc9l5
Z6qku2lOrqeuD4gZRVJhht2K+0WdSs3YPVcBjiMMaTKYFTQNbnJ2Jij7fhbJ+G7A31EhW+BIjHMK
Le4BjONRxwP6p7TRIpidXTSixpJxVITfGvWHZ6yWMWExRg45Wo/g6gUGqZYqWCGshu20EqF5BsRL
mrTKjXU94xJBZzU9pyok4TbOwCvdcGEDG6yaUDNUGymZrjBQJ7+IO5JLIQxzP/akwzUB8aRXth6g
Sz7rDauFxYhhkd/M5vYbYd2uaRfvK+k6mMh3+Refots7Y+Ij70Xo5RIuZ7nvob3LIGFA4y4nWq4l
J9fHq6zKWBGeBl0kyKOd3XWuIHrIwgJgonOao0xiO6Zv5ZvEZkXeodEoPPhR8MH+JIvNvX8dqeFZ
7KKqflXytFnv/z/f/UgErviMce+ix4/FNF3ybQl1l2lRlnT52RC5W1dmZlehSBmyz7BR9Srox2Xi
nf0BB/um7Anhtq6+P9s50B+EornTOPB9IFTBC3ljYgPUXCWKKk2d5aKRMQmDyTsrNF+g/t7IFqzW
r5omIM6pmVdsITXi0t2ytfuS2P9k2O69womoP+2mI0cK1MJv0hqy78h1jcmpnMjCwIbzL7MAzzzB
sesDHKQd0RC1wXH5IlrhXYnizBQkMeg+zdotSI2f8mcuyfTZjdD+93UPIEe4MQJd0MVP7Qq+6xWL
FV2sYS/bEgw6HwyDiwECM+39C1fZv4mFFPcs3yMm5nA5/6f6/2lLgr+jvZtLG/7jzrMo3Jcj5m+E
7Yr6m2UhRzGVIgXFBYJ7h/8K1b8owEOE3kWd3qR9vBkUhWQVq7lvoWcgDNT5FPS1uvIvLpZIDpeo
MlpKwkTAFFfwYbtHTZRB4H+8BC78z7E6h4aOxUXk+05Ah25MkZsp5ickkZPkb0A9rhQ0SEA+zwBc
IIl5lJd+e0P3ADzRVmgKYVm2EibbyCusvXCp2SO4wTRYiHzOTxvU5xu3qHaGnPi2oc0sqMRoZGxV
b6ybFMSgqgxqDdx5J8dTjpQvgOWjtBT3Qu1qGp8fnBeU9SjaNqoxoMPEBqLOudC8rX3JBxIas9GB
nXcFLTmmQLSLOCV0QRiMF5WGt5yfKMvGo4zRplerA3w0JdHJt74A717A0aq0GzhezSjNVfMLDt0d
bKcIDMz+9aQ5cJ06eN45HV/1SUzcT24SuArpBOaffYZcECKiX914yYRmY9Up33TJkANVqSTyB6tF
I2YBkreDnUa4Gg9wWQtvSM5P4pNiQn74MqtGsyeNvr4mHJi03703XFcrsmdoKUDcZZGmVsxcWxiL
aoAi0Wz2xAyZGcB93FXDc/gT8fbRLTUcfu7ePqj/3XcKxf87us7mFBqY4XVebiOz1ePDtSpe8vGo
YSAFS7tY65Io1b79FOPHCC1tXY83b7/kZH+tg02ica9jmPNZNj2DXX/QGgFMEJ553xaxbTFXdFwb
Finrt85N1jZct9soQr7kA0baQi1DdJTFNmIoS+aBseP15/wjS4JmKhuWjl/Y2UlAEaeuPcxDUYo5
cLV658WSF1ZWAroBuzSPXUxRWWHyL97RcDaw+2Si1GmW8oDaeQjHYTsY2s8BxfPDeqQ/0tq/cuKb
kNSabHsXFLHJF+9tbVF5iyMMhfqQTpeRMPa+PsEGZhy3fN62ouAW7AQak+2zCuc9eTgOESOb/ZxQ
858RXEk/4E6o7q/WdEEducAqC8+V/vKMwS1ML3BRn1u5HQ2mENm2RhDHvT3FIyvQExLg6YobU1DW
kGohweyy0RLZtFKO1MBuzxhvrcEBCAePD1im0gbKbG0Futs2G/0zHDffiSjyJxRHwcnKaCHB7hDZ
iaXo4IjEciyLIS57DAsLZafwldDb9a3yNcHkVI+vnoo7U5PUsvlTTkIVIl1i34QCGhU9EgZpRxpg
Id6gsPq5T0UV5EvC7lSO5U3ksK42ALXdgSsrtcAj1Prmi2BUKWu5UoWPbSTZMAQOgnI9JQBYWgK/
0AAxz2DPuStZr67dka5oJp78enApIQwNbNoPZUBrX5PyfWjGxbL9Xx55fcDI6oI+P8KUM4mZw+Mq
vY4bvEGHlZurgFl6yXuYaLig30exJwUFZMRheVkwUXcGg880z+aPnmBTl5Y6btA0CZn/Dk+sYF8L
WX9Xf/Zge5ZnHYIOInD0M4DmMidx91WPaQjOWNp4mxEVE3ajZClAz4izm8G45TYuja9rnrQQ6csW
3hB4+sQGQMUchE/f+R9I3ccr5P0LVmfvYxUWTi82aHAcldMB6Sh4/I3BziDQ7ryEPeeH2DL5tj7d
gJkqtXs+7w4fsUj8XpTaGaMWsZ5ROEs8LPKbbGAAmcMkMBzsrpbF6zHgL+Yb+gUImn5PjSC9gq15
nyp8hrvGO2FNh7i50XEkvy46Da3rfR9nPzOce5TlrU3qJypochUqeu8ZlsI9l9yo1KP5HccO0EhM
xDVNLLIN7D2aeAHr0G7bezNPllSgOujJ+YAft0Kyoh813KWsr5c/8TNukpDgkabCGgH+hQmzTICb
4YxvJ6TNrlZmUeiF1AZbcipJZ3Pq2Qs9WutadVLtOZytmaFNlRmkRs8ZDT7SscXFj4XFesdOxKCh
1ZA8ZZQ1tITClpnMoP6FgI0uzVOkfcZORB+jYyBaN94pRLd45fwzvv4Lsvf3i+yfvuHJvm3KMtRs
r1dnGruZA80eCEE4LyvXWA/SP1hhA85Ed+bfL+RYLXpzNd9T+g10nsoAHAg+yPukQ7Dd6P2xqu38
1ixvbPEYRO44iTqvG8+4I/dS/3NCtyndI8iF6ysmoe1FQ+iSi/urysMqB5xXd5kBoUuNs/oKe7pS
7Yy/BUvrj6AjpjYHofuJKRjcyRFKBJb6qmymkN7dTB0RXsscFz9Pl9c0yoF/CUYapP+ArdRL6vLn
eJxvVrA84YtvfaLUtKI/mP+W5HQj6sRrUqPf2WpJcPeszEt82O0GQWkWPVGZp6+rwO6Q7227uSS2
0II7T/hcX8alJgu63poiEooPwKgm8HG46gp71lG6mFq5+byritQnjKtsfwkIRbfnfx/HDQ5Fa9Mc
7gebQA5c1G/alPbSoUYblra1MCLkw4rorZvhUq/XPOt74QPrwhvatOrGNq9h46IrO0RTuLpe9arz
2pt004Whh2X+mBBpazrS5J73F4Z/0S5STukHBoBwKksLsJTSRgWUs8J3qTLsTTQ/pvU9j7fZpke2
7p4LzUbRjuYoVc7VfqnTeKFWYGS+zyl6czvANiW4g53Uutg7fdFKKpQWubKprgKVYv6xS+l9egw3
CJ8tcdSgwkevXpeuN1F6VWGrtqDO1I+nxD2mnGUvCrkAgCL5Q9G2vPyIJ4/J/kZdQung/v3I9Ree
KRbnTcUDQ/uD4FevExGUMAFyscOCErhU+n93eJI9n370Z8xsyARyFrUX1CoEbapupOFyy7b2vSF/
z6XEOOth2UpV5zFVzhhRu+kjLomkMdWESjhIC8wADuwPRe4vzSoFSWpdBjoOuhe9Jb22ZHaL7a1n
zMw/IrhBlaaTFLzyX7Z6fjnwpY+Yhsq0t19WgiHnWJHyTUcCgQkonDwzSbVHgWgWKh+yAzAZgjA7
d6O2mAZfUgS5obN4a3RaebNRBBvgr94qUlB3xDVKZU4qEpa3Qq8X3IiqwrW4Rnorq5j5QPkKzuzD
ptEu7xvY5XpdJrn8LFMNTEeJOFdoHMvuqYBeu0mNP9S115AjGhKIn6WO/+Skk5UtCKNB80mtkraE
5O9BjVlCF5G3+qO1ZdZXlKVJ7T39UaXRexmluI/+EtUxL6PKafyxbCZWQDVsMvLWTJr8EDaqgr8Y
KA12X7VQQ8fAjxTMFJdYgNyQt7ypyuYS/BVRTMea2+0/BCOovfJrvrz6IQvCT9Y9RL4Prhbi3wjU
t14FDeDbUBX93z77vgz3wnuAPfk89cFnemlm1PYimQcXA7mf6CDB4pBcPkK7Kd768u9BCylZYEVA
XGTFHZRupivrCfP8GPK97TbPy/iDjR/BPYWsQ0mhTU/wMgjOkDKKW0CfjaDVLL4grKFUa3GcpmMD
tq7K9peuzzvx+j/DKD9xKnXM6Bq11gRYlqJaquu72Bsy40iis9WspGt0lZRNe0VrCmsjPAZEgaRM
zQpOGaQF92MxpR6yiFqLuDsPO4PiQGSj83eR6Wmb3MmnnKnZaEWJGxcjnS3tEUFhhHWd+SVr3TZl
zri+161dH6Mxjw1LAcoqXFw8rVgHN3m0aplUUUeSN258bciXuSe3gYP+lQwy5wTnOCJYD9y4MVnj
PmwFwiaXyMg2yJOkZgKaAGCSvw1NSiw6LLlxb9lM3mRZVWIVDpZxZErSH6tBtU1f/NP/ggW7lEC/
r3No4foA1ZqZ638mpPVF/yf5rznQwmYgmnRcuDredfUikqMtkY/cPeoth01ccBTMJ+yICcXY+RyU
uoke67LKIV1RU4P3ZuF/9DIqViiM9W/ZHMvzdnbV+t2PGGxF9KBm7J/sYoGK3ZXgyyag0WOibOZh
hCj2jK8NSY5UIXZsn4+sqs7zXPyvYK2gH0y+mDZWF0IHJ9DSrNLsXg4SnkewjsPYzjmLyABvLdpv
/pGLcbGVp96NEq4jUn0gz0Vet1NPPNMBNJWJERdAVbz3egEBRrTbYeyCo2bNsHjA8M1RzkvMV5Rf
JKc46vuZudXs6ZmJOeOB09zOU+xPHGLiz4fOejAZ/NJKPAbu8pJ29wT2yFjWMNyc9ZiGq6ctKPiN
Z6vOP36BN1yQwuyBhRiO43SBsuRzrzTzJ6znDa6qAzsdLX8E6HP7AUj/8SRmWi65xyj0XOt49FH/
uUjUzcEAFiFTe7fiCN7Ju+60exAl+EvdYnZ7MSgAA7F3yoCIrOy15/Fb1AO9JIoHivHNA/dbA0vQ
5JCbh1+1N80i2dj8M9Ftc296PUr4WIVNL3Br1rQeGwDenmyhNB5LbYga7+qfO4uYAouBejaGFqy1
IJBX7pvjNk6LGPzwYj9rpWB2wuvL7zS8v8khWES5GglxNzUvl4KmI0Z7s0i1+uPz5NV+rBJ752qN
yi3A4AZH08R8Afn3S8g9qyu38IQT8ViHjp4xeJlS4MjeKISQgDFDBgoA0SOODOVD6VxwOVykrM2L
BX8QeASgP73v3H/d3scxsG4g3OF34v7Zoz3L4wf8LFpGo7PZ3pohJ9LOeUgd5lMZR/M713/LTmqV
BvhVGwD9+N4m8b4qvOXMWkD6xq1wuuFxXhwMjwTBk2qwbrXNkt0AvGlLUXxUPz43wsfxM4uHHkzb
6G+PH4GwYRYVWb6pwHW3sOrr8Xwx/QOnohmhES9SWlJhpHpwj9OyDdp5nQqp2WmmFSj9oRqA4H4B
xXRa7gix2wvU+AFHAh0R0ajK2Axj82W+XKfxF4swdTQnivlP6bRoPd8PA/uEKzgdBlA1ze1OmZQY
qpssEq4XNhM8dNWLe+AdjdpU86YNMiXIsHf1iYzQl81KWxyr5emsGhI8sTZ919Vr6UZsckjeMOaD
I4yE0HMPaCiCz4YgzjfAQ6evIaylCWwDJ7aoySDvOrRAXaW+dsa1ChREqjfhTZvX5kG+Dh63PE06
4455DKeR0e/kna+BiTlOgJfM32LZwFnIRStubh7tLq69aDj0t6X5cvEP1Bs/Ocidtiyj+/vmGI9r
sz2KjoinC8J7kW6CJb0YGgFtCIv2IUpr5BuhXcl830CvHT5GBoEVTX+pp4pdT8loHSzgD6EWUuHO
re38yzXhT14g2YmzqnKRFQvSJnhOZ5am8b4wU1zAGvUThslgK6792U5kqiOumyk3kFBH1WcfX93R
6s6SAjKzPh9VazYypt6yDenfHgXgWCqidLiOVDtIvuq7OFGFzZNksjmws4/WWuV3hcpI8VpiApiK
niJLHnvKx27C+xDi3WiiQ7lDFfXLT8vEG8xB3OFzl82/V1kEbimFPUZe1SeUHrFIssGsyXaNj+oV
agG5pTdlgAWvhESITQDpUwGQpO+aK/4yIPRrkd2cTwc2rOgfaQA0B/WDUjrgU1bJEeIKkQwl43pZ
YZOZfkRH7DOpsSbEjgPtL2eUvF43hHATHh1pWkLZH7vSf5goxS5qq2DO7TWIwjoV84T2xIX2eC8l
e9qszYxC9UhLI6T8Pi0f1J3zK/f2/FJEXjo/WMvFPpwg7HdGEg1jqMkZT8/AgLKI3EGsEkGX/zf5
+wSsJnTjfm6hNrxOXI+HkIt03ckEPfRvaWFC5+yOg7LzcUkgOzxzp4lPeEAe+iNRPeFc2nQ4Bevf
h93bulZKz/zSg2/KfvA52056NYVsRXiRplSd85Fc1g5FlM8bdiPMMBSiCK2jeAc1VV9TV5YYNqV6
oGL+A9xDCG8M+95CZUxZQRZkILATCjdNYFfymau57Lwc4Xqtty3p5AbPMv3omY7Mjm73TFCmfQ2B
EkajFxqf1sus9wlY+KQMPr8xYlb5p5brZNyCRqEuWNe0kz0HxQyvep4syKuZcC1QOm4LuVGdpMzg
sLHqPxUec/GWEx/Z67DknY35phHnIOQbvA5VGJAVROv9WqB2qqkcIVy8A/Nzij7CF/TPKqFWBceH
ujqHaI0CVHKVW062SrGqzZXMrMeYH9vF8QyTCyTyd77muMxxK5X9OP81qpH7G38fZspRzi8T83Ty
OQgLkBwJ3AAPf9IPlMi2eU+wBgSARhoQcxVbK3IkomydzywzhuARqXg+Jrcynxfxa1e4CmfE49Lz
Q0kuFqS7cekQazj5DoQd5tCGKLHyngIyycuVCsDT3LnVr7JhbKjTayFC+MI73V6RIUbnG/FouTIT
N0zqwX/To4BrlEaYXidx70EDsdAdlDY7ZniewVTUPqsXbC3DELceiE2ykdPpUGLQKHLsTgQFJuz1
BJGwHHN7dnOUE/ayp6uHvVEi2eZcY198UNLHAtcKAj66HJRFT4Y0oW+OVFLanDw6rdHUE4GwIJDb
10GYAKsI4KXaB4yB1689lLIYDVfUfB197EWMqm194W/6WSrDuG7Kq6NmzhuxIOwTwRgblZu5jMiU
YHYQF5vsdXdBwNWeXjhQxw0mXLvpzdVQ+YRXIBE8fJYeHZK7wnBoglhCB7ibwVvuQnakkRh2CRVQ
UuL/soJMItpjBqFrCr/rn9J+Dv5wirqetnvi0n/IJul0GcX5znmrMc/D+7iIV1jsstYU2ivmcxFf
UDU/ZeZQa8o/+07pnmexktId4S7OmTOzVUB28bREH9ot57HA3pHD0D0jQippJ21q4Hb/Iv8F9POC
rqBz6/YnMIidUM4pcHE3+yZqYNz6ZGdSBmrRVUkVEd+k2+j5Yc9vynCemk1K1TRrjlNfKmPI1kKN
lUGWTKgW8w4h+6F7bSnWTJzU3IEl40VltSVwIs84BGD97U/UKp4HEZgsdNJ2YJDB3JlNerViyxmG
m9HeYzt3+gN6SnxSVGBjGPeWRLNdWsFUVtuLx68kM/u62Mrbgx+lGeomI31tC170xbMao3+bjjZh
qe6D15HwmOrXV5klaV/3qR48nVYeJ582V3gtHJyLvH2QLCvqXMA116N9lxQ28Wsdv5JFba0HXOrl
lFJzRi5pz5mhkuppRhFLkW5HktocG0Rgdy5PQbEjxiwI9pEZpVR+kD06O1sJQ8lFM/JJxu+gDn+G
SrLoxCMgN590LtKHLThBgNSlVCNDK3vpraRlfWyeHieLhLWLty1icSVc5IQ3vWMOhpbk+dYF/1mJ
lwV/EnJAp5Y8GluypsRSIp4/pyFmkrXsRIwx5e3YzzrWKQq6w+FB4iTmA3SvRStinCjUCXWbhRnx
R1zp33lnGsenI+tVHi1HH5307LowJSQhnTIsQPJCzG8cfk+YFgzf5wEs4f5LzKa0hMfHxNnIMb/3
MsLpPIzkSw1SpYJwqLaDIcBlX6jo3Lxv0sldtRPwgyvJ523DfLKSY4ibYt8wGOCt8GAIm8XbESRT
hWyFXzkd8v/w3vP0GoscxYFP68f9qWLCS49GtQs+rm3lAUO0QQSAMpTG/PSwGsT3tEd6zaPuz931
CjpXe1bv5iJaHAqqSWv1+oL+BL3X5RFJRuM/2Q+fz7VgBjxOFayTI4X6UeFpwYL4nUZXriYgz+ij
diFUfS7UQGmfyeWIMh6XNy+U4DqeMgezYto0QzrJTJdwMVon1QFERPU3ZCAgOp0Pn8O6ASy3XHXx
u1EpRMV5DQS+vz2Am6CHAlT56HcLcBdA835glvajuDngPAc/cKhrg1w3lCQ4X9Faxdm0tQ5Da7Bf
oTqII8uT9bsi6pmQtCnfLNODoT+Q+9977YnUQbrfRoOSQJYDs23C7Hjg0yL7gs1H/Id+IQu0E0KE
dwqbyjPMSjR8ifM6visSJw6z/D6w3S3LbvA8JHmbRufyIXRvWLo/jv5BL/p2oGoaxkllvmutbt2G
EqiK4Uy/ddLyU+VBAoq3v7cm4SCdpDzUbBNNY0dCdvFM3D8E+WO1DVgJv4ONOHAPjSKkUdKfHDVt
OODtGFAYtgq+i5qWNPD220NDYTilo7IU1H+T64GRXQ1O0x1SXRD/fJS4hSjXmzfL0Imi6RUv+6De
XraMUSI+UZqGH+u4kqiltiaz614NC8rTxoY6EBlU4s7tnOj0rIzmGQbEFZ1JMpiUT+512wq4cbA+
gic12FMAIAfgPPqjBV7Ad70Dqa4KJD2iOVwDGrBVXCiii5wl9J0hC1eEktGA5nf3ANEwouEnUeac
rJGogojGfP67j94rrKZ4bU7QJ2Jyei8tMX54KM/EX+ihirauwJnAFh3TKr0m1biymIH4TvrTEAAP
BoQfQVHtzLgUrg4UQRb/ih4qJSYMluiLckuQn9KotKGS++yBEY/bkkkuw8OtdDDRM00bs83ugW9r
zH0UGcCYlkfSd7Y4KkWLrifPp3S2jfpz3M7w0zEGsAM1eJsiBb+5bVk7gABSLPIp+ZVsW3U4aQcD
c8YhhSAa1aLXmigZSLAG0BhEHSQdYXzBxhCsHo9n9WMw/uayKqMyxieaQn7h17jV/Z72mfZtCHwL
MJwyoGmwMTW6l4ycO0MP715zHyjTmaI4g+C/Jy8LJyK8mGTG2326OKXzHZ/Z3QMME5TN6C2UKXo9
HUM2066/PliiR5dKjZTZwL7El6WXumXjHFCGRds0KkipNFKQn+zBJQiBVVIuF97C/AdyRbMs9Yz6
tMzBLvBNsVB2poIsgzFc71+W9ggFysoDgZ/lu6nMl71qWbtvwtq7/3m0xDUvwKZe1ZRSwHd2rTqb
DH+1No5hRXjxKqNnclYt6BeTLETTB6HyE46o63G85x6BWNkICW/uSyX8+DtDRrnO4HWySw6BrQe2
gySz58MY+dnCf0zUDRVJBof3JDzzH02i/z1ypQXFa1wFiyqg4dkQVxcngitMDUXTRx4W5/qstxIv
OTKKVuOSmhjwCF8ED/y0gUDFu9DWOoWtdhAIv9lcpgD02t7UZ4Jan/0Smpsk0exNG9objNUhQDGx
dOpKn1X5TlF9tv2auRnrDPTy0KcMCGXwbpPuf4lolsDAH6Rlpk9yM77vyt6Zfiq+Mt4U5QylcByY
Svgq6LrYkY0zI02aMIcI5reiNlN6bGO1vMOVKIc8e5Sx4rQmU9VM42MCTimG5wvdbeOcWQtq/6ZL
N8l5ZmpD58uu6kHWu9MSXk9Ik6W8NkcHXIJ97nqyKQD3bjxNU/RTDtR4helCzvM97Rwy7mX6VN45
hfJRC2lgeIIiWvIpMi1VlAf2Ic/iA9orWlvPvG1sU9AzpXe/700Z8shcz1MCNZE7XPoIfWMv1/19
mR87WopuRvGqHr4HXYOy5wQYYC5wfJqQwUSbdq8gODff4pwVAjpNzs9B9qM6v4n25qthfhd+EZ64
6BjXqAjGY/393RFRG1XPI5HXZBd0OCaf+UwFDZdVt84tSRR7qmQUW7Z97ifhQEO+FkCC3d3FYXu8
UyYC77UcKGLHO4grymIrzs029F1SPtCJMqDIL2HHo026NGEInkonPAaAB0g5KBitHcQNBdW8HuNQ
deLVG2SY7XascAO+yrHT4FsTyCYxp/AiyNRBOQ4bJyIg1tc6RXxr9K9EyOmefoLF2lAIA0tk1U96
1QhWkhp/EB1ChyS60vn+PhleNczsLuJSj007SuuV/GHF21t+k01+/sJ3mQe0OYPb5RMkg3tIi7WI
clhixaZGcE06qeSf9UL0oPNdaWPlZO/Dx0RE6c5L2nqn9WMvMtyC7J8zBFDESSE6qEDwlaI7MA3B
jtjM40+jSvVxxytgicFpSgu/d+4EF3t/LtGsQ0LZhOpdLi6591CaxyxcV/cUCgfZY55C2LSGbrtY
KOrE5zSPNRXKRzwbPO1OwZlphr4QJCGTh3vNloaF0bXiokoepvyE3vl2e0UBXUebCiclHurKPVY0
/ZMs3OYTTvjkqfcIMUiY8u/3KehmdXpayR5PFvhFoyd+5yFqA0jv74E1EZVzMAjkXnGJfpOlcoDl
tSRtRoovhXAomZRr6c5uRcjRag4Z2hFqoG+NtbcN1dAupkwQDZ/yQNOJFc6i4t+j/RDFAGtZdF6F
5k5/aZWzHt1B0pEWskpXLKVptdpTfyBaXRpQ0Fdgx1/tCmhaXFaWd1l5I1wyO2DuDFeCi47u0yj/
+8Z06PlWWKRhdfUpVpLQiYIUGX4zRlZ3UqbJ66h9/NxQJ64llNZs6bq+Ykf0XiG7csrJcrLxM1lE
czKiQuvxwig+FRAMgl8HqDfiIUvWnG7zANYWNVJMdKsl3R0iKysx77dpm0z1aHJN8xb3SO9sXNfV
hx6RCc2EIlcyv9MiacanTeel+P7Tmdnj2TyZgbRZXky75xbusCb2FtbVcReASaW3N6Se9Dz30fDY
F4lZCDp8KohLGCeQWse9gL+y5cWpfsN3K+DNSYd4eipY83Ho5Ec/DAfTLjVKon2F/lwmOflCG39j
JdwTixWj1RMZmZa12qX9XMm73QbiX2aDOzDw2er2NSQIH4KV6hTXjNK++67XktLRMUMlV3hKj1vd
+1Iuy8hxplHes3vXG/WhIuTK3hFaR1ySCTehIWJWRZLTAz1tCR2FmcmuYkmUChPrdZg3UJbcZf9Q
QJHtdnHqN8yf6weg47dzVDFkkpCXB/zdxjnw+KTWkPQblN4D0rEaNnQ2Kr6kqkEs1RgOH342J49r
HB0unRHVUDY4WrWmUlG2P2NjbR9bF6eahSRoMgTfjzwO5LIYtNrj4zgRE7tPtPD36NG+4aPH9c6k
L/nFcLU0Jw5i2v00xOXI3UKfCnU/50UXRwXuNh/rCa7Jxb/VVjKaqsnspcWUsjsmPsYDdjcKBDJi
yVZBpcDLU77vXvV9dxWi92to8JO+o5RHmv3hrWN1ZTgRW9fW7ObaYNpjuxt7htocPrfPnfRktjlI
7I1pc1fmvwv4TNP1sXaKD1X0hulxlsg+UXMmkwfc4BaOpwX81cZWpj4zTc9poIppnihWmCvVcQ6X
iRVYIhebmJbttWv7qXMWZtD1gs8oaDhG2eDs5LW56CxFNexfgYRg1hmop39PSgV7eJdjY3BUqmFE
Bu3BW4BsCXIJNIDWT9WgGeKNRLM+9vQZlP9vp5ZIlCz8H7OHE9cc3AUcl7HwZZexeUBKlXblxm8s
ZqNoskZ4Qkc/Q3TdoAyqWWcIJrtUZSQU3HeHBsitAFB8TIl9dq2jXGXfpHDqsIMbKFxdX+8NNrxI
cVZ8ekFhqrGW/qpAquDah515YvUWWKB1Y76fnL17Q48EePVkVW7wDEHaZ8EeczWnoo22qBUyYgF9
urg+OZwRbyukDL/5M4es7jF2xUTigsB6HPNdt0BjNiJH6KKnOJ5X7Aq8qvJFKGIFeGeIaT/XSoWt
RgXXuXBASGMdJHWYKtgtpsCLQhNgKKL2nNdcwusrObi/ofblLdMtWdwK3PZqjASTVTk1PRSL7DRo
rzLpsbBKZsdIlFpJnxu9tLwyyEBf+KqV8jC2oXfySDcNwPPVFhlgWBSaKYsCpS6VPqDdmJUUIowF
x45kbT//BIhsx9BlJbOPymiMybmcNnLsqZj5o5tv+wns/TlunCeLL9pt/D2IvJP2bMgHpYCN4MY1
axvEtTKcgNZ3I42jOqO230/8ag9gDM92+QG3tVCkgIsafCiKXzkAQgXSL0EmTlbmTi2c1coKbHc7
EpHwkaYgcSVOIEhUecqpKChaQ5fykO1UEp1+Yh1u+JhMxbKx0PuCtnVncghx4OCa+zkDYChYmbZ3
Nnx/bNQ/tg2CEC1N7ZEugwSTE7QgcFIH1OOFqcfmI2gGZcp4j707mrAQt1K046zMvnDpwO1Q2Hyr
oKK6JAeMmgg3A5KwaZjfMn+wAPA8zzUNCNNnFlLA7GqaawciOm5HC0C/XedzdySO/ZaS6bwQUeb7
Bwm4H9LNzqKnXrRwrLWHuSF/XCTpKwNlt7uqaXB24kmPslimI6nmnliqZfagDRgyvLpea2wqdF4w
C7TMgvKsdFS6iHNDmdtWoWdLw+M5yrFAcqf2ehSD9dwXrldLdwIICh75HZjjwDYKM3RRmALVkVOW
RpShKsGonQt1M6lP4u90ReNo93UJ7Qw0/9gMAIgwhiKFGxjBDssPCIUhpBHhTJTTwORQ2/WrIEUd
T1538sgYSbu9I06dax9nPYKM8voT1lr9r8P0DrR+IlResIFaDW/WbSeY3UDKTqL8hJOuYgfduVqF
uOQNMSk8hU9x5+fC7Wfq3aMIhA6PPTzs6iNu6Jkrtu4POOedY4ajrorB1JYTFF9qsb+2n99Vxy5/
SVSNVNrQLw4GeiiM3CeZkPgQQMv3e/QVXjkeZp4kd8jTMOHcEr3EerQhQlo8SliwQqMVaNp3BGAg
k2dscMf9n2TZX5CoBtS33PrUgJ83S+0SCHAo8n/eXo16eyzDXVaeqh7HO9YXwwyPC8gqqFR4BDFD
Q1XJuS57d31Ba/8OnfbC5lIyq1DNg3BNVYCxAlTg3hDPlZ4s3UVnDVmbFoffI7RgedVAk6Wmf9Bq
YJfTdVpuBW73xBGUe6oLNRpQyz+6s1LdjWwshdomYYHO2OLteeLxSYuHbPtof3ZpbnVcJazxUtHm
KbITW4y0/4ffXhJOd6mnXuarteAOzgldBB3zdvA218DxvBdes7PlBkgiO703VXqPdW/pCtalbxm4
1SrBerrD6hf4+yu7bKRPnImdbiXFRJUaw92t1KN3gL/Z8EkVa/mgr3e0+gp1dMCZXvoRi8vd2Lpd
BSaC1bX3k1v+5MUXZev5FJhDlYlhjXnzbK7iBZAbB96qgoSusWqJLbDVN3InUdp9QXdhhXm78w+0
pSJfuFHuyax5OI18x8aj1li4PdD4gC00SDfa/+IQUDYvYsM/hTlwozYTLPJDiXZg691K2o7IvHwD
SSazsV0KZ95ikLWjBFP9FmI1c5BjD+aXwpqvU7dxFNcMDdBwi1FGQ4zeOnkVoEElJEoBWgDhIiSR
LAlrY5ZYBFLBLYG38AxNfdoh0UKOUomLG0Gd6Uyv/Xm+CEdOZJMkliaBdMbH1ADRmlaq6TvnH/+R
VSyk+8SXijC3LN59jyWUVm8LWtsHaWnm4eDL8gnXZWZw3sIH98+t0o1NqQ268F1kVfsbdIjeDYjD
A0KYzgosyzaUadwIYM42Dnixl05nDpypmJK1FLEpuDCn9P0Ta9Y6a1dqaqWuieRV8RDRW6tNIFcq
U6XP19whmKWyJBm96wkVTmmr6c1osyWSp3mozEsUPW6UGtdL+BZWe6l3li3OB4g6MC6ngNGoWAQb
o8nBxtlui8NZ2EEVFQ9RCjQ3wrhJmumT+nnKryHBAZbqTeS1o0nwEW+9UcPc9d475UGPvYdxr1fg
59m76LyBFPtFXD/LEMlIp/B34rPVtQl0FoSgTlu5nz4AHuoHyZNowJSo2PeKXWgf24M3yjlfzVdB
qjOzTS1JDX8GdMJNPdy6RLcDOORhj5jHd0tbo6oM67JOuiLCOrJubDcwYU9sBiEqwX6iC07I1f1D
nZe/tnqYtUmOEwdQUxm+XA1uolgTLDEdnt3EQbEdomjNUJbNczsxJE2GR5yr4U/YSjavCZpAzE1d
+CYM/TrBa+h3/MebHHDqTG0qm+swQtqwBHL02odwjNmvABuFtBQWr5qo1XVw2pP3Ieo+3KS+lfbO
xjFbp8iqkxPoG5d6ak8GUVPI6wPMlpWiBBwufUCdpX0XUjZ4/bVK3k1A3EfJGLnJKZ9b6iB6N8bR
d6WcIGr3U7o0sJTELNiIZiuO4ZcZfVJHYlrtd7r30Ts5V+hEzNT22e87lgnEGfRO05824+ACxtPp
nOXsdneDCT0GVFXMpyBrm54Rt4ybk+E+ZU2cOwBwu/CPUhOLYTaq5BQE4tqP8qsm6DQphrQnkpVW
IcWhCJEFFzaJ1utk2k3shEyWRmDk7LZFgbrpL/Ku4uAojePL93p5zcSnt/OHvdjspdkr/WuXoL31
baOpb8WgVFS25kR7+2t+nywb5i0iHJewZubLzFlqIVEikzFhFA3JpDw2JKIfIpMvB6aMXGx5uI/Z
XaVKtclpR8gabIiRCv/7xiqCh3yVWQ58DjXyfe6W8bw4vBORMpCgozIJU4gxb2eoZPeoI7E5VTQ+
vMtbs6qDeFkUj0cw4k1ZA6JmCyC7MFiNl/XcyTcuVnXwqydqrwb76/pRNt84uH4OmrRqfGivtqau
u6Q6WeLzNJW1c8CIZNNlHsjlchgAZixsDZB0MXz43V0L4oTv8yJL7xUOuScf0RUORaq6lN+VGFOi
7YInwbCJmTDgWH3M/3TL6Zkp0PJZT1L9aw3Mo1CsLnihSSHJb8566di1pJi8PdPOsHFqQMmxFUQt
k8vE3QM7H7AWeJ7vtrpmuf2o8jO1eT84NPOa5cb8vpAxUHbaRrBZ1EKGiOIJYTUhRHE+SfuXqgYG
hchPjDOJNkyT7ww2LRMxLI7nruSJDb2lGd47faB+acKyFEfyj4bQlbumwaJ7JREMxk4O3nO2FQpK
rKV7NOl3lQvjuhOaMPhSZnZ/SDaeQzrKpOHg5AFsi0i3THei6xFC5sEp04r7Z+vv/kn1xl/Q/y9u
LMrFH27FcqQarMcyqXC6esLSbYaMAwExkTwsMaK9H+PMu2r2CntKbU7UX1xfbTodLU99lmkKCsft
qIvP69xmHz5zZK539us3TBLpObWmzl5rNRLfhUgUGnG52E4TN3HxJ7wU/Fb0pKhgGgHjlXFlhlX0
P5AqL2MvgHkJXgYWd94rxijHBlqLY+/3gZplmSuVYnCjvikd8Y0eEgHvxuz+W8XrKTU3fI1Uhhgr
hmezLi4N9ug+i2w7AVo2/oJNwrUhI8Ej5GXjTWomHhkZs3V4t9bqiXW00FJEnL5bRqOiFih7BtVf
Y7kQEKBEmOLD6DQAXGgC1teqI9bXzXWlroBc0TryFxHyGVCuAfnXZ4eJCh62J9XM1kcjlV7P1dxR
PMxzdnlESGgKnFd5hQTzrJyM1qxHHXbwNWlnn1VmVHk6jvoFGlvS6tcvNpzfHc6Vd9bF35Zhv8Um
H2sNOIHsvA/VxcVMjWMk9AqMvxzNM1hWa0mmx2r+As8eYytavu7NqJ7euZ4RvZ6LTcoscN0JWO0N
j3hx1l9QOzO/FnWFptOT8CkOWq9hC+MUUctWGLKeDXrGfAa8KG9s4o0Y6Fu3i/ah1wP4s8hjiRPN
BkIXOoklJHpOHARom12ZagZMUduK14yOxQYCsaXZnjZP0zUYeIG1yuHjgGM2A+kO2KvdmcKfw78Y
Ux/ijyV8PRZMC0efuC/hHfIV+TiTbuzQMbHmyFKXvQOpWEcDKshulsD8BVpME1q48/n3vs1wxcq7
/BAmnRcakGmGaXXEpN1CyadNPTveJ9Udrx8G07pXdohW0LDLzDNvd+u2BXmrjWpMoTYOeiLaFD6T
t7k6rJn5kaYCgeJ1bZDbdfNyC3BvbjzCYLGrRzw0uyFkrFLgyY53jPGkvt4dYj8tTDLGjkHJBqtJ
lsMXdYp13KWtLnK+X6mb8tUAwVYYXOR0VHChBJlKEV7ODHZTKOf6jvMG03Ix9xBvd6Nacx5lgxB2
FFENWUzZEgzpsGr5xBRRtQ03QK29oHvN4Ss80GX5Zex1WPqhhvgexb+E0Uco4cZg5BNDvGY/1mTm
J9pFx5B5xPSWw3T7WLFUXXi3RClzMXIC1Fwk4zcIngF+SiUTjmwnUWBv5MSnc/5WwsPheHke0Qyf
/2nA33DldM76KLD5wFC9h53Zb5uL0ZMay6e/82V7Sz8lTfuf9XoLuQeOVO3ta8evIHi5lI3vzr2c
L9j1llROtkT3uupAafp7JGPJF64yId/cmVh1fWd8Vt1/XiyS/jB2c8UCcc7+Yz8W5gE2H0Bv0OOd
RIMOZUtMqbyKtRTwfvXJdpDCaVZTUBvgWd0bcwlNfwi1Bz170eHTUOo/MYKQjRRYv50Ab5inzzw9
dEIkGVu3qLbGzLTCPJdmq0a5ioZFeWZxmB6q1bCJT0aixyNJWdpE/jBV2lil4tBqO8K6Ky97tcSh
RP5vPOI3Y425aj8ekC8AlN8Boku6BAA36Xs0hUYaRfxigdLfcthN0cCr999Ujh4Fznegm0g0+Xwg
y9+NaxVs45btejX3JKjO/xHUdx9nkdZV+51jGKlPZC3nIK64sRcU4enUCV6D4/Gq2yHa9I7ujPSJ
Gra/HDxPAF9i8oQWkR5pu8FjsVoj3XQDQvpL2/qVYpzSVvUWlsuywrmNnwXaN4pEp9iL6ABTEVYv
sBMWt7QTjdHDs70O2GZl3GIVcyosjDKW8B5/cFCxVphS5G007qMVvSID9mC6jrruf1UaCzSQOOiF
WuSfiaExdIHTtTDlKK1jsW+G3V1CldUDSXfRkQykbXffwq5mj1nI+URBGOp9S53nNVNbhnyn9fan
N8YgVazXg9E3YypZQiu7l/vrDk9Ff8344LOujzRvJLCjiD7DQyjcC980bog3ele7PhB3ejDZdO4P
LzPEruc1ET1GKBtuDvrFZlU9qJAqvXrR0CBW6ZW89lAb3qfKoX9YOnx5FlcDrz6zBd37uxEOYnQq
TA3+C9BpUriL5a4guH1Jk6jFzzIAUzDYKb5pPI787zQx2cpe4x4ninn7Ou8I1HAvy9bVtdYqEV4H
tCOz2U12fk9yiVGxNN7o62iEvxLkAgzHyYfWaOxfzRm4J7226HJhF9y3LE2Sl6YjLq3pU3YRX3bE
3eEAnwgPvzADdZFOqK4yKAxjdi8SAMBll40qikePUXF1yigC1PS0grnCEpfT0woPxpbjEK2FIdB7
UU+6PmSqBSEELD+pnFo4jc127ltlY54nGE1m66rSR8fqmHzW0jkzzCG1Y3sapvmYPZA+7LUb8p6z
2AsaO/dua/K/tXJA85D31JhmKekNt8GLHo34EjZslJuNssgHCYHAhZuOqfVARgAlmKBmMMP2b1Z/
T+2Uh15m0mrzuzG0NxuYzJBBa7FLC6jXjSv0H4KQDRDNwUVek8PvkRzrzaHTT4flGFmPhMe3NvOj
Bj3Srb704q4rIhpZ+YC5UpbGvYiE/B1gwaKCjl0wXqn/1NZ1vSu2/qz0fjnK0BQ2KiDyEzOo1DD5
5fthp593feRR9O5vVl5lutxObT37WC4kvK/D1X1JKRcnRNbyc9XUVhRiMfhed5mohv5j18SEZ/CJ
Y3X79Wg7Y/a/qdztHrZBhtYN5iJ08fLsNH8ksm0Y3znegCm5FkWXwrvBtTW9o25riuWxxCrf/uRV
DHW00AiJA/JXvLkv7mOJ/y+znKaH5uwuM//KfWv/DoqvIHgBXkhL8zNSZDWAq2J/0Py7E9OgliD8
r57jwWpxyv825Rdm6zl1oXoQHknNwwrFQaDiS+v1sUTCdn9ipFhPDyLg6AvCxsnxLUNM2ZZPQgOP
vPo11aZ4hfDmJS+u1j+mL6YEuV44Ysw6fU2REfTIBknyvGgHPDDQI/13F5HZow5WzoG20dF5HLR2
FHYnaDIxZP+ZVER3wmvuCLfdOO+SDqsm2FGHQRg7KsBg0s63nLSBsuSYbctEXAqFN3ROq34P+Y4C
X6/+slkHFRiINkzWnXmvK/dF4mh2zMKhi7Y3II/6U+0d52ymDtcGO0x2QF8a0KhDGD1Aq01KAl0j
oqAx7YW4ER1PkpR5hbHsfsILr0981sYwgl8j86Fy4mzXt8KruPuQMpGWKP8cByKqd8WSa8RTZO7/
fSoFzdFNdrukeTPjliOFLjF3C2L/xMx5kXsZtcewPW8v2xzOT42wJGMjyj0+NfRy9JyunG3imifb
Tt1ry4nWnQjcwZu6ATMGVPDNkOkVvbAnG1DQDuSdWUJzaJaTaNz6mJvjAqZ68IDe9Vr4gepWuwM+
W5K64TpxNeNPG3bz+QVpoIBVOfLIDmm/BbLDzoY2p0K3RoOn+CY5VO2AwGxP8xaJQdnM6MV/UN34
B0e9fqC7MPE5znSHH0gJNCGILDmBLPveCWUdz3aGWOzK16Z5F1fbZyIwpBZnk134UvhryR5mJ4Vl
ahAQpTooWyW2hXlhud6K6nwW7QO1trIgwGwWS6Lzq5WaZTG/maREfp02dYEaxoJ8QU0Mv1N0CDHw
VsJyipK7QCkZK1PWa+AbHKGgyXXi63gsUVRnCFSHJvQ7tmzVjwdlgvM3+mO9ntEf2BiDnwFj2K8Y
lFGBNcZOikYDWRR1x8scb8j0cl90nZGtbE69Uh3S+7oWUWqHPG4EdGkPUNPZc3zE0h/B0RLNXikp
hYWZnrEBUwar/Zx48/F/+f75QeEpVc7IWK0zhCW+OnfHgaOkXElu1BIXFivCaJAHEQbqXSYQv4DD
3sa4EljWVjEmYk46+R8lULCcBZ3ea2C44cI74HJvnhIJqkru5wzbj5o7TtXW+JQOWIDmyPfhalhk
/Z2MnXHPWAYVxvqHX91Kntp+tXMyvK+6sO7IFsQgI5up9B5FNwZx/f1aqKW9uTGKXE+3cGc6dak4
Y8O2cxT5JEvNK0Lz/7twJf3lKPfDE4gG8U7vFxlO70tSwJAJrBDZJ9xJ0gahW1MuOS1AF8jGELpk
eMpZO8vZ7AtxeU56AYxvP/qL3fey08NXK20jPgZKOHBE25y6Umrx98qPQN0EPs7mHf4vqRjUwwfo
92awukomfYFbeRluELQ54pDK704MiP2F+JFQSXi6razCgopcgwrUCSe07XfW38J55JMZMopnorCD
AgJJMLQk59qRXf4D2/moYc/RC1ONGhhv0ASlqMkYa43zGXZKyxevVfgmIhxhut12y4c43BRaPqdH
Bk1Q/MhV83NXG5MZMFcm4QUem0uFRMk0sEgDcoMfrBxZBKzgL7X7wLoEWuXlAraLdZ5fpICWqdzc
kfIkCZioxR0db66IMXdgJw/WYtn+aaLiPHHoNIM3Mbs+1cqiXMOjUU3QvULCjRY1CvUMJNvpwJTT
jVDClBvBChxtD3IIel+j3ZpO1HY95zmVBbcxGA2iK7IFSa90N8n/2M/5i3GdisfLBK3lIEQ5nk64
b8T1fXKUoineE47BdiWcHBtC8ZUrz1ET7+HbDOz7FTfTi9IM2wMsg8k5jRpUghMKOJ73/AqAUmXV
N5PD0m1DS01FqXNgozyg47f1GxUaMqozWyKNzHjUQKzHgWqtnYjaZq6Lbr3kY993P29jfQxkoUYn
80YzFwouYXmkj3n3JvV4i4Lz4rUt0i118a1Xs765qqYA6amqIXD/93yTcPkQSRihdzZQ/C0GbHrz
OlG0oCFeg4jw12KkiaBdfFdRif0BMX8QvEu63ZOljopeaaGsCRIxe+lrX9Rms6TDbUCjYylRxlSr
NKKCfZWD6E9k/JO5+BzORAq1lSyp8t/RR8Ptr8X2uG8BggncJlY+ubJoHJlWrPD2kZ0y3Nht991n
iAjOhWyIpB7MVCdzOVZqDjk8ykA8OafJZmqKW58Ad4MBoF79heCFaVD3akltZ3WUB130XQJSTY5Y
iBs3KI1bEpxOVP8Ps9bgcishvg//FBm+7xlu2ie5TKr6LiEv6JdwaPZxlZh5nG2cW4W4c0SPfHDV
s9HaL9DZszJ8TGnmzRAT2mbNwoyj3JkS0kqxL5okLTP/1lzNoMJhxEN3qEr7luPa1wR1gGSTWvuz
HPYIE+3HEQE5ks24f+WLAAt7/UMOrwmUtPSW2BHvVgUCLMPvQi7QqiZ0gVtjKA3+MgyPHDFqELXt
FRd3MqrcR1FuxJlNClrN8ahxxYgqrNY20T+AavSINrcsRXUa3QwSmoTYIgGowinKXeRHWnpJL9gn
NeunBzrtp2+uFlmtm2G4KVP8+lM8tP0rkP79L1o5FzQ5XnaZHuqz7cJChKUQat6eAU9gIMoNNof0
6gyDrufCT6UsTMRaC8+0NlYtVELusBhq2PPf8GKpsJNw2Rb3PutyxSIf1vVIC4yNj1hS0W2+KB6n
I2jonS+/rGrouPWkuwNmzns1yhMJpswl8IMDd2xX1JgyvoLvOELVVcmOYehvRgTN6bO17rQeFaHM
tChzgS4syI7pwwD3Umb595mXDR95ChA9M6MtRWcbA4R1p28MBV/0E46zop3MNpCyjSzDeL+BzaHA
bD+Uo9cX25mNuxFv/9ME8kZHg9nYEHXbYXKI6kvXHtpE8Q6QGkb/PykEfFO+4TdnnJOArRT/Az5Z
uw55iCeGvUju+lf/swIsS2vBUtBC0z3uVFbTArJM5bcQCpEJg4p9LNdmTVw2vVoM1+yvDHQPCO8k
eAnerLpIWNS+7bpGheZch7yGoBUW3udFID4sx/pOuT0g0GjyVe94Pk+/RSY+IhbvoWvWbzDPYQEg
tZ3WyHpNzolQuXI2jyKpnzix9egyWQYhG5/1exceeeN1MplN7/ULqJz9CH/XqHnpGMq3XmgkoSNE
2KChvQ/F0gSLkz3juikWrViTaOt+6HejGnG3FbphU6BNIdiWobgJm2vl/R+SXHsjWfsaMV2FymlL
PV/qfMJwVylkbAJBhh1sfEW3M6q79m/Z3WlboVyA1YQyAtPRe31l+Imdzflo3Vsm/Hr3oDlNq5ro
5UePzfuCYoK/kwXpBZY1p3EMaGaVSx8bA5TjdOBiSv/hnUVrwPMV72ZM9FEhXg6LaD452ZTmnRrf
ElZ4d7xkyTZILYVU51D3HDxIV+ebWXlqiTXs1Pitd9iN63l4b9HG2Hbzny7hSS1AovPcKclfhbeO
i6MAK5qcRWxUhIAloJUAlRGswaNyhCtZqCIRk9Hm1xEGG7JRg4iV1KPjct84dtx5ZpLeYdUWW5Wu
iQyvqqxivzua0/RSq9UlHr93YeGVBaKlJiZrA6AggNWrLk7pxSPlJNmnnQhd9aLTZhU6pHVg8/ej
xLx0JntFJPmAx6hoGukYulxVghonJKSixdlj+gZDGCbLkgzxQf8lmwoXAlMGENeuyTIKRDTnEDa/
Njma9s2I8GKE2QEI/4PZ39OJfULnNhTx7GKIwu9c9chpQfHBbpfUVzAondQ2SceZnL5J75U/SdKi
ellMGl5QuGe1VqVbxQz2RIqbSLPPkS9IHHvrmuCycYowjYI4I1wD4echdkNBj2Zqo3Bl38fMiBNy
3eyjOWMLO5G1oqng5h7zY/7pVq3bJ+JqBGj1tVOPISKiq3dyrKY0g6MiT/KC6QHxRCv9igmT5JDo
36//bNz8wZRZXpgPraOW5pzz+DovBEuoREbeF+JqfRsMVAtSc7qoHAAJeiBm9zJ3LrIygydOvnRr
Az4HpmDgVohZPM3cSZRswO5ZJLMZbQG2b9mdc4ImTFuQWpv818zqturkb84XiwEnd8sbcZ6sjI2h
Bmypw9A5zFndyVtZOSYHXdPiKVJFgKA/XZGgrUHL8x6oHITuoh+sdFfaYnyepRFjp37M06NIp+Ie
0BG7KbGBLVnKEEINHcGVYEI94ywLLtkdkR339UVrGgPsotPTFC0ntglWqzfbGxvZXhwkfxr9L8wA
4o2UGVoqv2wUdS4XSIDvTTWah1Qr0QM4wOweGcjf3vSFRWTaGJ+gU3BXQVO6BRY4KF1xnqkLgOWb
osbzSn7A4EjWreomZ5z6SOdPHygjcxRTguQQD5drIz4z/u9MuXux48tiDRBGKJHKgNaE9ckbHJ+p
p5w1TDzJOOCn2mQ/Yt2uL9YTBCy4TmsWuotPOwYlNiAeTbfhVLT4B796J1tk5BHuxN2LLVDRjCEw
GWH6oWxu7Inwt5Fha6TgYMvFBMXabVa7Cgn8gqbvlKox5KDxSKLbQTKNjKG1V662HYazDWBSFXrs
rU0eqj57Xngo8khvYhUGJhMXIsSaCS7gw4oYkWbYPSchVtMhhTQZs4L+f3dkXRyZmgwjTqU69U89
tjpYNtDMgWVdBgAJ4V1WLh2rTIsK7etVNEoFlAKTrXDlnBE5QV3LQKcS57BzKHEOAOcTI5rY+XCe
bDxkHAg6DyS8OFu2pP1Yg1oOBP/ebfCwRmQ7TFef8KuOxffDM69xOr8Bd5w34NPvsxy8rfHcrKh0
CzjelMjpfM7suOCMEranufO9/X1uhZWnHm7HBxrEUKe8DcmNos8gXR06OYM5WY2XOmFwTU0h3Hsh
Nf54D1Gx5ptni9eWQY9IZyeOP0Q3ppDs/yeOQLTCOoPeDSDjSG8qX+MewfurvihIwUfBuTXVvkSL
/xLMEemNY6UHTIBVRz+FQ8j6ADKmL6t8BrP1k+q28ZqGFReDFGqJnQb9bit5K3pRuLEDmRCSxmyR
xY1erDpk/dOKpZVyQN6Fxr6CIiynELSMEDURPO2/gXvVbqIV5pBAJjFX79EgK99ykSbPsiO4XHcb
Pan1R2IP6Mq/V77yCdRRywVIHp53CPM7d8IMwsTDwI61DIt6OCyMGz7tg9wsN9BB4qXlmYJkzDit
dIcbA1TzjB54mSzTd9h9nYeB06cdJ9kRLW3edTfgxmuWyo6egnoFg+BXuT6AXnaC4tWGlMC1ZpIc
D4L4diM6HwVecyvbezOky/Oglomd/7IZOcvmazJ/6va4IbQxLegjeu+j/t81wkTXfb3aLprp7wFM
GPR73c0oERgMSlJHPXcUiPBHTrfgt11xFdnjBVDYzSN816Qzecp9AwblMWAXtxxQOBT2bJjYBxWt
syDr50HB+otJ/YFRyTWPVd6DTcFB0WTqfrZtbrSHB1PPGJpsCYgDFJS16bHG1XAJv2nPJRO1lyvC
chRTMlfFEnJQ9W3/4NcYX7Zzeewf5LZ48Be2aPEUXqm2pUEKGfpqmUQTpKr1RaljRPCcSrKhcPBR
9HD2isugsOBegHJGhN3HlSb+bNPdByjv9QyxHoY0bp+i6BmBrbMFGwvaBm50qZaqf8UaMV/jaruM
AojTEfiyXVfr/Qz3A0zkXmdnRkTqCitcQyJbN14NMa+P3vaWT4j4aI4d+w1+ERIF9AFUgG5y4YSu
AH8kIH2QZB4RuEl/QRfmC+2DHlIn6VNFUgUYLMbw8z46UHVr4G60bn46xtIl/sdLhp+KIWUGC7+o
7WJwCUIJrn1QtGJoozlocqK4rKoHUg79tYSQNHZAjM6C2XUJcrl1DQtQSy7VXUALJVr41K3sm8dy
ENnL4sAmLvvGoMCy06ufMFwMS/1fEfGNknLPlGumJpSSjs/hi+taMy+YB3QyJvz1daSZeqJ1mSP/
R9PDStJXLOouUHhqwbFMVUCvsHg9HSEw1rsMIFg6PSs3pWzw6pUpxByPmdZMf5Q+0RnBDb1U/En4
Jw511663auMOUSHCod9O0qnUAliOpdmmu1yk/wTfKPJ3PCpAazhSrLnRpwqQ//v3t7NrNT7V6/0W
PlcRNhc/+0bj/F6ysk+hVuxC8OwQOqQuPt5Nyk/zrkytUWO6XmwIqU9xXuOeE2vNSOeKmp+uZnhM
7u0JNjUl1M3Gsblg9yAvAMorvbRFLsrCMaQcHPMcsWvPe7bBQ/AEz/FtZmBiGAKyxipHueAhkmTo
g3MaUSBVQB2nJIlMLeQvCI4lvgpJFxYRhm0vfXjbbDkNVQ+yvaLNlA3cKw7jHzakWjiRgTSdrQZ1
Bic3saiMkbSKK1Ld4dpp0WuXCiZlH1YNKtLLIqsBzBVJBe1OKhVuX/6SPDCFtfYIBy1e/00EC4lm
BEFjskcq8Lh3+hx+JHgvcMggkPLheBsVY3INjGLY/QVlyRsm3+eIXX0PVJN7AlFwB6eq+5B7uO2A
L8aTgJNcPLYbyIRBGa5gIdXZJImt8Q5twiFRuG1OWEIzdaQVmiEzUoPsAcXyU2hPG5ORwYMJI9lM
BiUY9ZClGOnCtdT1UstS1TyK2Ox3x7HDvxyyLDD4oCSrQud6b/nqmUHG7awk8SStJmlKxYwOE7NO
hIPvoQBIFbNkum90YMIE4WqfLw7zFwo4Z/nvJQp9b21PlK12cb9gnGC8xuDg1hIOd394iO0UPJID
9JSczx0rv+4g2Nqx61cFSD2RyBhbg4LoA/JBEG8Ttsf+GUxR5sG5G1+uFPlQGgOj+dxzMarO+1uY
AelY+qRt0MSqStHDZ+wMvEXyYxiTcQ9MI2W2GXJwK4bSfWS81PzcbRFBHntFBsGdF+pG3DphmGgW
/Nn3lBNb1jppACiik+5wS35g8a/fYcuSzWkT9r4iFgldZT5wToDDKQO7Bo/Epu6OZtcQl1s1ga/C
SQYJEScKjPSxqgXPEyu+rP3cDwJeYpyGkIj9fO8ZH5I2zYlBXorZKBZthwyIOyRMo6nx+srIOaQg
5ZLN06Q/9MrYXWLjE7cWoXKU8NWL+CcoFgxA+ZAFBL/6mUYnFkKm163vs2d0RjHTHuOS97ZhiFBi
EeWnjx9vxByi84LzLNOk5sB9k/Ul/tQI4O1cn7sNGGtJ4/bSrLXMkaWDZb1WBCQcyS+21KDtmnS0
7AKeIWFQBjK0rihBMEMAAujUYN/qHpiAt1a9byXvq740qcpDjbhuxr1gGndfn2vHa38SSj6cI1sX
wOMbKT8HNE0xlcbQoUnqgSz3r151V2Et3oP455iVG4HxBCGm72Ru1OoVyVEFIqVF44YojGrhJ3sc
7i2uY4cAyW8XwrZmegOMImKFrb7MYOndiV4++5JfFvQf7zj1/rEaKiWia3+ROBtw2kMtFBE8Q7tK
MZqQkBlZnZT8dSJpQU00j2uivnP3d7GpDpx2IK9sD3+69fdyF9xPw3F5kpw9NsQp15YRDup0Guqj
K9wVsxBILvNgUJaox+GqUqs70GTVG/7fVip5ihNgTnPKoFedRFbp3p/Q2ynkkfKTHrn97fhLV5vA
ZlgvsWeArvlRyBsTM9fbCHbjV9PIbZuX0VVGmngzo5AMuYI+XhLL4DLtk2a+A015taZlJ7Qj/d+y
BYx6BSTp/BW+OMNFL4p2E0NRmowukUZS1c1sraThSDbDfq6WiQ6+AU2eKGPEZi/z1VRU6XX+BLTz
dxYKH10MUJ7UkNI8t0uVqjTzQ0XemxWMLW4SN4wj8TPZT/gQgYkPSegClLFm+BodMQV/U5M9QDrd
KLcsUVsjpwu0WNspeqf8hwu6PucAKjAq48VnGVxWZDTfTaqx2dnvOj0g+kjoM7XkEbV4zAWdVWBZ
2LkO+Y+BxyNX9WSqkYJdVs1v0c3l7nRfACbH3EPCKTYRhwfFz9SAgtkYxnhntgaWXSzU3CWkJ2nN
B/QYOhkRzuv5A1Z0V2D1GvwFFd37SUCVB8yE/IzJ4WYLmW/g8emK+Vw007e3gUyz9cvkxk4SBWBw
5Im25UJU5TNWkg6W88205plqfdI65mmZ0yT6+7i+74ahyYGBg3RE604jbOLi6d2mSvnaXNl/8LkH
DpvzRnakI+KI7HKD4PRzaJIdl5u5H4AT+LUU04UOTw3orqackpsy0lIMRiYlS3kJM3xX0cTLOgf6
eiBJYv2GTZxDJgiEjgtBIBHPND+X4S8HOIrhoU7rif2di9Wlid+24tunwgZbjb+pH+280t2Z4pP1
F3JNX8d3R2f2PWRa84tNN0h0XjLbVf5WQcpOnscc9jUcJF3sKN4FsWJjwOLMruEcSUILrMPhQJHC
vz/gEfBVg6kKz8fnTjrgVSOwViiHw4FyoEgADkAIYLeZewNtyTX27+b8wLEhCBua20xYhfaP6IpZ
iT+Ww/f4yorZZfvX7ljq3D7EdnwaH9K8cpINHlks0xehEcFwmjGimaWx1z0aOpcFZ7bwQpyGY4Pl
I4yiGm9oeiFU9Sj+2Zp61Hsh5ex+jl5ZASvU6hqG5a5gXIrMiut3q7Fr1z3/KuH0cubbOl1BaZ+w
JSRfHPEnvGB/xIIxdNRZE3TFyd1+EGBYYuCoOizLgQiVIAYcezpGnZF0H55t+nxls2g5+c7+SE3x
1+I/3k0Bga48meMQ2z3tcdPyWwBBFzmwP1ZBpPRRZCBrnM0wULx5OIKd+ARVLQBMhnnQSlAYjwCE
PYyJ9zDt5GBIyyPmY7WdCBW47rDiMf9QzrW7rrFZfB9yqShQ23qLbDTUbiJ5vW0QrRirE3KwTlFm
CruwSva3Tm1yoN+8jOj37Vft/vgK0J+O2U5SMN2FwJ5pm4bVXzMgv8jPjprTDGmAJxbwBeJVns3f
w2Md9njl8Lks6380wQ3DyqSZSu9wIksMMAPk4TQ2YwnQ6xly2Zl4yGX8V1NaPaMfu/Yp/iaszex2
fwbfzjbeBBqgT3RB+iiyCjIr2T6BKJELbaJo+0rMg8djsHDrC9yaRbyv20fNRGKgAIOdmybio+55
pvjHShApmnPQdRlaGlCATRF76tnizz3AhK+hqXzoyHBs6E0YYYZAib09iVcUyB1Q1i6IUKkIAHq3
KYz8SLD6sbdUJthiZCX+1fy79O0ZcyvnrkBlXyQ6HdzhgHOETfe8l4HyJpKHjzLhRJEJrxeDfX3G
ht3EvJtqG1ZnGS+HU3SWTCoCNT42dqWL9oyGBH/vRQ2ahqOKz12AIoYQlLQh1SntzKe78YPgmoEn
9jqeKNb4Q2rnlhB4iwPx6Aq9fQpzcaw8QuP7mS4hv7zEegRGkxT1p0axu2oA7AQKMFXX6kGNqKHo
3wbJzzcrQOvJCqpk9gI9vzCHK3i23zJOEF/qcV7FnXm6XE0ckSwLR+dv+9LqNd4sG5Vwj5IDLFaI
TTnLLk9QtjgeIbEQppqmZl+CzH3JY7HFL+j9GryxiDJH/YY8vRMDEHue7QsvTEEZMx0Th5Mw1uRh
HTNeL6AuHCFq/DmNQkHLt8VNFYrc+gxYXwym1dYwbSQTpfHvMeK4jR1oASpWU5OPRO4OBnMUtWvm
saNZvuvi2ZSxOOW7Z6sve5hFEPC6oP6F60lCueGwnAm9NtFgUL+1BvYnl2nswycqLiYu9hfmco9i
3RkNyH3llcGVoldHXY5pmnA5JdaPY4hvbeMEOYd5lMnxS6l7gnAq8fp2IGD9CBWDPPWM6C4srx5H
7q4GqPKoIGZxpgUrlEP4pmEHfmA7NDAyJAq1qVATt4a2GKWKtQN53vxZDQ9cRsZ/5Mm7oo9Shimp
kQczEWMV3WE5lEH0XdnlFrrQDNMwZ7RNY4sS5HMOuQ0cx0QdbAbvaUmUm5UWtZHiaPKFZ0CNBuUS
LjjsC3q2NGp+30QWhyAwGfvbWyc0BqQns9EOKEk32No279KyfRVAyDQunKf9sALwkUIxo8c9e03K
7B5pSjKG4g+GAOT4FQDbrF9HgGOazFKASGjddQWgk6+mZh3H1m9VWxHLk52XAAUMqsVwFofebShP
+XGiJPucz90jDMtn1I/KHinp5VMp4vl6puSE5IuSbyGGMryC2m/LqGHEKB+1oSVp6ePQ35SXKXM/
3/jwnZebphKXKjj/9uvLkyZdqCn3qLiduRya7A+khNMAMyGeegJCLDS3kZqz9CePSuQxviJNlKjk
I/QhPNPUVlTRuzbP9qxWTmQ5zJ0M15GBqz7+r04UU1fZ6RT+FmP/jpezgDodIukxuuvAx3//eGzY
pHOd6mhQ/tnMpFhHFLaihWQlWvsk6n6Z36IR1s4v2AytljTq+RCbao75pxId+XrtRsd3xrJYkOyE
kEHbMbEF4g7QFYNQsmb/1SbdmQtS+vFXw7u0N5QSfbicaiJeRaiwR4u4E6ADdO6Llx5vQYD/0Mpe
IQP6iCudUWedCukrFUkGon9eM47TANcHRIwND079UDrlM15mR9Q3C9i9UV4Ms8ALP3Jozce3h4hz
oRKTJf7yVSAC74GB4foS5IjFhf1W+gHhYa4s1S3+tpnjvweY/t/+HaTLTC+NqvM9hGr9jhq1Yz3z
x1zTjRvhGfohDwNXHMaNfRUimA+sqQi6KzcvwlnW2XpGoUlN/7yCO+bnMpIv7uCzNGzwtLpv3qH3
z8LIPB1btTmPFjJUbdj3tUtte0f/1RvKSVNLuulNY6s3CA5S6KKQN6S8l+5TBsndGH1thLWfr2JN
oXuV8Llyf+RBNTuM6fVjjzG1QVNbX4j+0JOqhJIBKzJY5xdoaOr25vJoVRZUYW0GtJGL3N8vi2Aw
/6eNkvAQ8mfCJqDel4BGDtSQ860zUYLt7ZsqcdNj8MDKEBAImH/zdT3bwO5olxj2gW8UP+TaoOJO
GzQGzfzNydBuMQlsfpONfBI0gjvQU+wJiFGxFCd1NbeaV+2yeGcXx/k869+5RkLEtHMdTTauCia1
12UkpjD1Dtw9mJQnOPVZJHs5kksr21wRQuFQjHkTI86CfS9FGOXS68yPTYMIohZfTE+mLyjub8ab
KHN9Nfh8knIkWDZiYg0fUYaoSqW/M3zqrXG2+2E6GfuCJMrs3g4gLYKubppywiaxWWF5WhqT/btK
RWxkc7Yl6bxkVrvOCXywmC9KOgIFESwtWKR8f8mLiMUmyVcNYaFoiCl1xR67dzYyTp1pq5QGw2i8
s/am7SHd7NVKVjcLHF9ZmR6T2EpzA1T9hsCbdUYjZLCW/C0YDRDizHJYZsHKboZt/VDrttezx9gl
bRPoweMWVE8xzaURQeUGapN4xcYkWVIE64doThUljJw3MI2G1zPyzwgqr2AT91rZiZxSfOxon2oI
sFeKtejlQQeZFU7mLnJJlW3U4jWb/ic7G8Fwx4pMpm1RxnGltlPWlZukTV2ej6LmwSMld+qivnS4
9NThIYee1iSNEVSwxqQ1vGKMCSIyoDsaXp/DktvjIPi7wPmwzH3ERjx3AiGBM1RmJ2KMpOIWp0U9
4DJj1IUlZaUtvk0meU+qYoEiExgxl7M62G2NJPoCsIA+9Fn5BmRY3SVHSlzoYXqlGXDT7exSRaq9
FO5o50TJRXnwkJe0c9+CngvNPZeNPoN89q9gQq9Uhj3hVeN3zJWITXNFl4qkxpX2RAjjDZp29jAU
geiYjmaE2qf+1Vhw3xc6SJ+5oM7/vZoGWGLPVFUexZq5HfBljzpzTYLBiflj7b7osqpBr+T5/c63
YZF9pp4JSwTChW2P8EI6yXi3nO5pacRXE3cD62HX1zU21sOnzfJPphye94qliWHcLalVj5sZ14Gc
RH0a1vemBPgEJ7Dy6jMe0xTohnD+n7q/mB+RSKzqcDeEMqObraTGEnuTy7NimvJUbps3cBQQq8Gy
JYwS+a/FkDBQhpeE1GWFSKX1gutCRlC1eRHmJIUMVJaINiQeHF5hQsBRGFMO0+IhblOe7HUg3wbk
q8SaBh3MhmYt825OkyMSxtBK5CkNxPrw4ZAFvkm2bxHVEfyN3k9QGzJxqJxELQEz+Vc22kvc1R2h
FUyk9OvCcWiL4XL980ggt+0nm4CDJLLXidEMFRwk1IMnnm8bcxclW8HI9QklS80obE904JOygrPf
WKmQwnKM+HLiYqR5PWUeX5t1CbSpyW3zbWT0lgmcQcUGxWMi0VyY0/arZl5o4sMb9laNudx9mKY9
ELJp24p4pco+6RG9X8WLA9I44z8dg1+Ij4XWaadj4ZBaC7KQ8wuW+8L1uwZAjLJU4bYrF+2x0Vkq
8AQlkY5ZdFEO3YaY4MWkjdRmENP3PvIQOuqKNvCNvvQYBtLIgnm+ABMGlWYpnwzgQXHiz9s7Q1JX
A0J3JSMuTbZNDWdzL88TA2003gKR0mAAEbqTYJwfWsQfu8q0TtebKh0za5e5W7uHEybnkoSFrDHQ
vBGAefCQgkELm+JfFBOUnA1QMc6jkekzcUrTyFl46OInEUtJ7bK+Fadi0Akbke19LllEq7s8bDTj
HT4KHHE3IWSZg2UmS9iSgNHPlU363i3tVa5cqWTeYhSpyp5/qDoDh29otmemM4qOL6KiTGSS5eDQ
9RSp6aUKW3JRUxGg57zhMSnkEBxI4O+gOCCkmQRx81/NtAOSd+s59FUZhTNAbq+/ULbg5DNWMrhQ
S2d0Uy2anqzeFUPtNlbo8iSXJmUjAW4tJ7wey0zH1pnsH1nAuflw/2fYQV7xd6sZX7WuehZa+oG5
ruf84AIf3FxyF2ZDIAHFZxlE5Cgy7cEkbKWfhfeK6GFmZ3wxuBWBXs5pPQzLSPrMbX3W1MyTcgvx
sHKcTYMFCRhN2IWo/gMD9a90HnxbuyYMwZtlIbyovsE/67KE0SAU2BwstzqQ3ePdjDj3TDBNJJEf
stkUJ5D8h3fQCqDzTFD17BgyWHvn41QIvGZzHws9qoHcBJH9rVrLtfsFrlMoNyuepVcLV7XdNR90
LxvRqtOwAqrVzEGnMGi9a7wn7iTtiMjn5kMhAUscC8BiesxfxNF7iwM8PgCW0kqc3H0HQF55bFOI
8nHy1kyKo2HC3+5zca9XtlrgjZX4/3QKVVAqJ9Xyl5Q4WH4U+twIVm0WsMwOJ6FLWzeAU8dMRVhR
KFmr9Tuq1GAEyEpOZuS8DdGZHvbu02cRwyfmI1IZtfevGgGLXDsUqbgdr7O6jyH2CmeSmV4E+D5Z
/Ma9QgeXTVX/7prGaevWcTffxhyeuQcxiroKBYhtlWVHASZIRQ+uN8zU+o+BWNjY+9QWikyw9eXQ
fFAlad3wvvfHVT2YxUcDGYYTK7UIllJuD4YJ2ZBqzpkyrFp5ei/7d4zWV5JiD6vYG5uDiAjRELmY
su+koSmbzCQV9x78uoJGEZhdmlCi3WwjNaIcqEAXE5EoS9SAAN7daLCwBKEJXH0AwR7a08slwA6/
1I95HwIr8o07p7018Yyp+az2tqfKFUL2jlfghJFD24MGLgEGyJhSz1T8/66JuIlbpSABjtH8tlXf
59rVFz83xalg8pxUpHgDsW/OM6aIaoUxpz1rAw3XHGrg6dwbmDlqROybYcxXjHEhr0LsjM4C4h6f
OJhfTr6fUZAJ7C73dJTYzJXXYo4QdQQH5B+IU0kbZYT07rQAV+pWRH8siLI5+nH8z3UHrPbIE+g5
mKJewuT58M0f8cOZnMTC69V6PSHmWh+2N6CkPhOXGWHVmfcQF1QCgepQbvY7CwoPVljAMAl+51+I
MgsoZlAocY4FgoCY2MXiwhp6f9N4Bo7b0FOBDgdp+URDXxq2uznFdkRZRNtrQdfJ6aZvvKjkaQ0W
UFurOFcZQe9+3XrU1LOKCW4VNqqBeWlf6/NesfoxueHcIo8NUecw2EixPGhAYaug4OW/bs4HxIng
71DdoSXeINS7Yx9smpZB2RgH9f5AjD15N2bKk+TeTv4urUK2jfCpVChb3iZkMyvlnzkt/XZa1mWn
ZQanSGWQkTeSh7wJTdY83fHsvwBZ/g2ROk34+SIHy3L6gz8z38w4uzWZmQAOg8sv/OT26wEdbiWH
hgbfxfEyUwcO4qKooE7Hxtrp1zKaCcw2WMWbgyCHgGzd/x63cnLg9yi3AV12U0MqBoa6hYlFswfw
y2x8HmYtrmXClsty+Br2tI4oXKYeQ4w8WxeRUJmY4cEd8wh4xgf/YmR2uc7EShEcSN2t6IUWqGbm
G+yk2N2OAMG9E+EtXN4VhMVr+zTBef6CpCHlyAvp/esS3n/TOjmQyYMvbhG+gXqJ3yQip7RP0CqT
j7iOM/0HuPygsagcbC/GG5zfe5OvcjesPxB5depO5G6VpZTzbrio1nCHTflxxQpugCu3uxZDfG6x
EVQkJPNEMB+SABFIZLBG85fok3r/3omsc7gtI0HNjDZauIKDur5htEJo3kzBtR+NtHL/LgY8Kfjp
Y/zj6o9Dy0SqayC6GjWCEbf4/A6gDR5Ot+EbJ+VIZz/f2VHBuhT8WlRhlq7tKYhhNnnVfbcvkgQr
UXdRfa8JNDiPuo2vV8KKtFVJdmJjEZkSzDpGno0eHPVCnVgF/i4pKfqSxs7nsRhBWnd9E8isrjSx
LC+ivY0xXUqezCuuJhbihZrsmOCd3Y7vxgalC2IB+h4iGBeQ2+nIMLuaEvIg9m11mexV34HfI/k2
hnLBKwrdNRW0JmZg7p4SXvQFby/A7Jy5lF/KZxjEnKjb2C7S/I//avU2jA+Gvw5TaEBID2oY8E0z
a/lOjJi8XoYH4CGiuy0iErpzaj7Q7a4GVZs/8rrprrzv2YRRUHUAwFr8nAICFhPbSoewKzIo53B2
Ufh9I/oSSSZBx3BI5T95FqfZgN7CR1qBu4sxM++F++FqrSArxM7wn9PxHPl5XYJu8U2azJezfvUo
Prj/X8SFSIZufGM7u4H7eYlnFCY3GCm4Ip4TuK6nWodBal85tGOyBuK5uBc4WMpCSqV5q3gYDjrm
tlWTEHi3KikTSeEgq6T5mFpskPERR0TkelMxF7pTQetnpEc/eWf65VeV6TdrWPTxG4rYEi2LkofB
oMAFrWfVnk4LcIzYrmu8PAmA/D8wbyulVbv9UPydbiA7Bb4CN6fi+7smDKLxnppaBTGHwLLvwQXi
AatgxqsAKo9eWAR9YerbR1Y4hEEOVrQSVKTH42+TpdD1FKGDYvdOW52ctvhjwR+nyxj82QecyqDe
IigYtirm5naSg3JDp4FKq1oPu/wi+roCxBVGm+8TEY0028NCUWNkERZTVCvF3JW6NDkSCltO87LW
ynp4MR7ktdOS/zg5X6ysUXq0T5j+YPJUXr+5hqu3UlUBQKgrdqcT2CPlmt5MqM3HFs1kckCRCnhb
NVMoe7jeB98sM538IrZNjgWkzrKLk8JcRwqYLPKuqXJ+Z8Ho2GdluxwQCr5JHFsY4OxX1aMmTicN
vu5C9uR2SO/L33yCA3mXXNWJCh02G3NTVhsDDMUglDxRjHGON6Q1Cqd/quTRoNuXCab6dspnzyU2
yO3d4snQzf6Xu9R6w7vFCQ8iguuDp8MtwcmxXHR57tFW9tc+AxX50j529hfiDp1ea7PxufgOSN1m
2KdcIRJG8Zlv2gG8LQXYyHchlhtyMjSH+BbnyQ+XNIdD3rVj3b6F9u/74Nahg94mSsaBeyW2KaZi
EPfWIfX2Ocw6FWsJAYvAxqZYP3CCTrV7owbduCD9hrtloH7l7AvnKM7cbCCRVDrh8TGBknqhrKrm
aEAmYq0XwMpXXnXhf/kslJnf8uk885cThFnOuma6H3MuuQX/OphuEr7vVajQIBTm986zp3S1BXbD
y0itVoc6jLucjU9akJJifUirXsEF7Ok9VpWmn/OYjDOKuR1wwkZRhMLsp96RuGd/QRVNeV7D5E3g
Y6C1CT0hN5VRWdGbmQevb4zZkSCnhamnjje5GMruGtUD6TOHAt9x1n8aNDnGmIRYKHoWTTBN/ZfS
8t0nM3lWVoedA0bhoXWo1PpeUSfD5UqkaY9Gag+6ODzdID6vjkawGu+HGgcqwOB3i3kpthJ7icVC
8sogQAX5eQ4g1Z05z8LV7JyPb7Z6zMCL7v2ersYXnDbJEAVUhUb0pZHCg2yBZB6lyTYZTUm2gqHd
D5xNss9S8/cnXL87wfmsNmE6jrDzAY5V9h1J0kCX5ikuwyFtMN4+zH2XFRYQCm/B/NIEcUZ3jFsD
tz5R54xneZYf+Ob2/hwBSnj5ElAeuEcO2C9Hh9O/jQ15RINGfnZzCuHkOaivW9QGTSnuby8/OPTp
EACu9L5/P5hSpdZnCa4H6Mgpy+fLQhppUfuUAls+qGao0c8E61wykz0L2yQmpLBPIFiBbrJjVbXm
ri2zKyatu8tqp6XcMAk+cqEwV9cPTEqLPxpXrPyccxNjA9bSo7ixRFHVuz+uIaTJSYPThWvqu/IM
Usqvr2OUHYoHMNzsRcf4BejMpG+jCkRV5YXEPD6Otz904THOB8RJHUSuMNH5ye8ZwTziR9Lvu0yQ
aiOoJDRKKMvxE5BJRfn/nLHKtzOCqUlrFIjFFtS2SOVw4Dw6DFu6m3TESAsp3/EQqgMW4wOSE2B1
pNz++rjY/kl6u0nTfmQSJDacjK4rI3zoKtwmmDMYXopa7sSL1FG8oi/zwWHYNScPdqa8aHRNV1wv
7RfhDEoAWbc93EjLvt6LfWVgmrWRo3AGvp+p/FBNYd2YZkDcJ662nsjuxbPH1GFziQ02wvVjGUrR
JEkl5NuadQPaa/31vS7GfIB7VElkpG7M0EjMrihG+oTpSw9K2GuEPe71sUeeNi6nEdMUW+wb4/y3
s8QXeo+xlRUyFzSm2vAkUYPqg/N23rKim3c9BPWLL/Tv4flyQKzoMpb+2zl2cfUoQVMS1EUKdmUF
D97oL2Um4OfK8JU72bVWxaAoyyUAE0wpnj/NsaeY4EpXzrVv1106U70FHn1F90qy6Yn+y99Q4qMC
yPEXTahKONWP4xv4df6bwY3bYQ4Ck31jT0eWed0h9ZvvSG6+3Sk4V1h6usH+tITqOzrPR7p1ltqo
tO7ic8u0UMPIj3TyOZxYCeECvalmt7maOUG5TnhVq8rOQ6U77ycDhgfTMxjNkWcAVT4ApAYXkOuw
XajxuCJJ/xeHU073z3FzSYt5DoS30NlZC9+X2trvrv8FfWShq8DzBWC6G28mefk8QJ7q6fpgE1e/
u6abYIIu/ib5AYn//cyUU+yVZN3/KZ4VEJj65SdGsTbt0cvZFkWBaxigmOIq+psbTG9KFxZ6Ij+0
vl0++YjTAtRtXkbWZ7wrcP3P64HobvdYveCn9cVaZdS2zJtbmr4kh191PucTiB9KLUStau6lt+Ll
e+cyVnw0nXFvNDGTDPFyl0YwJuwTzGysFn2XARYQ/amdIII3/kxJdcaMmGL1c4gzIJ905hwQyc+n
ELdl9eIuKSApuVf3WqY1IaEwj2HSan1MTEXdgqnO+Bw386GE8hipnwgNv0aFH92VCrbt5Grey70w
Yt8Lhkqkkrua9nVV7oBpxEGU8MpndULa6NAlyyItAElyZOsjHErsKAw1wOWNfw0q+2418gsqOt08
ugN2GNCR1Z2tXsHqxSLS+QRwUD4rNu60MRu0DzuWJs6VtU7xXBtBUUz4uZomMAuTpK03IQKKHnte
St6L3xG6WpVGp54h248lLDFj/3ViWmxqOR7GlTnW6Kgv8URYdh02Q/1yewiowvFyK26MqBiS5bM9
2Gn8GHv+E/zkZRIXUFOuizeO3+seDWJ9f+X0qPMqEUZg7ZuyyDmCn3lza+gyeIPlqUM6dtaSUIoN
SmkTTpjxIlQjbO9oXj/qHc276BJIwAcUzm6cw1N65+Q82xHGhE56Ytc/h0Y4pY+H6i4a9qH5x/jg
yYjk05KrNMCMRmcxl1HzldjlZQIuBQB8I4wF9J69ZB3BSIE5T6VP2gEzJScJWnS3pjTyIaR8y6sj
BqlSP/wt2fkZKyiclZxPYn7Tux3Yz3h4wevZo1zUBj6GKMVHhjyslN0B9rL+TbDl+t2mKmPYU8V2
8WV6bjgXbmP+oAU338/t5FO/43KO4hsJC7bfkxVZe6zXWR0So3NdRwsNKYRDtaU69uKLck2WHBlZ
I4md42J2R5MlAQxxPNp5R/PLrw8xFbf/iMB5EFjXwj0SCO/OGv0q8bFrCBmJy2xv3H6FcFuroLZ3
uvtUIz1Uc/Wmen82GH0G6IUEgxXnu43Zfgnqdz5hRYtAIdS8oMWti7IH6s0XFQQn3kkVXWJbcE6w
XG9wEwJNvIvZqK6kzS5mzTPpPg0PsbvDuIU7nCI5a7LwXuD9fX+4TGqWYxHg4sFk5OyxafqiJvtC
+pS+0Ttahs9atTkaLKpIO4HwamjeiV55iCt/k3EkvoklS4kLnHlMEj3l8AsULM/j/Edr6oNwbFD5
ojK4QYK3NhMDK8Q7jWYPL2Li496Yr0kT5txsCxW7vafgKuqpC+ZH2A6HeaOfxJ1ZK7CSP1gHpzlv
2Z20LatKH5PJ7HFv42i/QOJAmWUyakS4UPZEFNs9DJTfyj6R4sa2WoDqKQGXKLCxDwgscUunMLFv
vWRv6KUQiqaj6nN21L8ZAmUmysTlNUwoEY0Y5qJOvABhgq7lCNmW2UJENFcD0jvHAUzxO+HE/MOv
t3xnResZTkugWEcHC2XjGCwPZnlsc+6t75TJKV5HkPl5v/qr4G/tu135yVXIEhYR10LVuwWIkw+c
iHq84+96EWLaqQ9Bv12NUsIN/AcapMrKKoIfIsDJ6GNq2GcJbIGSK2J5So1o6eXELNbdFS5ziB7t
72pJPJx7M7JO4qT5jxrxGOhVgh5SMeBnXrH0lDrwQh10K9+nFDFV9tla2K2ASHNhqkD+ZniWTofm
qHbv6Fj/H5cMuWPgBpGZHqVOFRr0UyYhCGz3reft4UythdQLfqG4rfGdx8sdvgriS+aK9ObUe+9s
TO4CekTlEf2RgFtyZ9OwhQXhNcrvcjxU6e9DsqAEpk8sDzQT7d6IbR9+oQRPs++XFQ+FvI40wy63
AUlv1WKIOVeduvdM0jgwBhKOYVsNPwxhSQGUoHGWpd1KPDjp38E/iK9GWLEoNJjO60hRtnFqTqug
jT+BGC5FXhA1MNT+Pcq4vaSRNUwK7dbRXsUDQw1Kwt+hKo4zbJY/mMlqIlHpsjRi0u0s59xWfQUm
ASDAphEKnkJ3R/1b2oYaF9dZKt8lJvEZcwZRQbhNKkfFKD44VWUAUh5fMgnfYf1h8ccw4mjNDuSS
5vJAfOz2enbIfiYWJP9dLMXhSQ+iCXBjBcjs9Tezcxbm8+lCD36Vq8cqYlITQAIY4tkg1SC8KwBC
nJK5bmEPhIgT5xs7gPwI21wdsQzOqB04q1UAP0t64yYIIArIsYcmiTvyBjwr5OQ9A0SGgfaiA9y2
44spTLlNoZhj4fC51rNow6fCkWzsMOFYZ8FXXR1tIxRCwRxyFocobdytAYVYXog69/WW1koeheb9
0eXjPZJjE00xHfILLIc9IupdzBMZOX15Ta+lPsaUMamBKm4IHJqGpD+lehSj8u0VS+7bXile2J7f
CWEKxyQe575SCcROE2ASMxgZ+QwWq0JUV09KhiOJ05Y4NrrL13FitopSkxPFoZO+z6FLmH/wqj4N
6kFM4RSNvbW88Ju6EeeHM0nKs72ot5r59kCWI35DaOeD8VqrqyySfgt7VcbK+R40rcmOBhUcEmRy
Q9R352nf/ud2hl33mc0/gT2eql5Aqagm+PP56lN0x2HUqLsvmsvJ7COzuN7fOJ6Gsj2Wovut273X
6QbIddKHeS3Kl9JFfmOaqA5f9TdQT3qtMGemNgak4wnMX3c2LaZJqaeXyi48KrlGFxtAczv4dNlk
rr5+xAy9Kj6nlUFTGW1nbWPWf7xgAS4dRxocTOSSkttQbCfgp/40nSBGmmW11CpNT+LSbg3esUTY
DlHi+gVpeK4ZklgJB0GXbWAcfS8TiSDkSc4WSFA8Y3a6ilF77ry4AuYkokFSfpD8wS55Bw/6wVzD
WCaACO2rCcYMsBdl3OeJrNMv9vOf81Mq7MXtJDPlgzmk2cRNFWuhdnZjrUHJItwPYRJUMq5haSpo
BIMAeVFtClJzBJVv5Bdqdhbvy+pYGi7d0hEG1aFHk2Yo89kY8JitmTRs6HVDy1FWCovzSMzGHO+H
qhIXFi+E60Ppt/ojeLnHIajap5U+dGRNYxAuBIxyGltoJTc1I3UCLaxMS6rivcPtCGc6xSEYGKsZ
NMKy/PCCkKIE9Q22XcMP6yO78aweOvM87v8Iq7R789qOj3AqklNksPMeosV1Ev9DZabk2UzhWyN1
gsKFBnpTfTRvA5AfJzIKwP692CiWWAVKFlhn3Os8c57eRHJsJ/ibwaN496NLziDywmULCAWxsfCU
XvI+Z4yCWo3Nwr0XV/rmB2D72ptN2P5Xdryv8OoZK9qfX8TYYeWHMOiARIL5CN/uAb2ax1QNQGNY
47ypm0oYoMdfpUcZaArhl3oGywAPTn+P1XB1AtonlCfkGLqODfqF3d4JGfXwrzIzxYMQ1AaYrbD/
ExBGm7cUvM68cGUhXLAn3+X1dwEQVsniX/jUWIbSQohpKmANsgRxXFPMwMCwFHwj25DDZ6gvmZn5
gFQ+zfKFF8W4EQduzNflnt7Fg8r3llrM/SZVuq11ZS0nldXOAYDyUMMUjkRNq2MPP+E8zziFgOBm
A+EFt1tzzTc+098p5Ta+z/aE/K+D4tHtR/NnJpOEEZMrjVf928whOcMxoOAggD9MZyNgnh/d7yau
4oH17J3d81R5Lph429ypgqAdt2EiPWcAOP9qwpEoGSP63IwghEa67D1KbAYdmJgeeutQe73T3W4p
rKfX6cmAII6YfWh4A25J8WB5YwHqpY5fEiuXgjPBahL40nOvGBfKiXxnU+SofaGkI5d7fMfu6JPD
2FRFLGhIWjZnSCFZ+P+w4Oo8RdLPRHdbpLIMCw1C4R8jWR2CQuMWyLmtH3ezt99LAOfZieyz2mPB
f46azYubwzKUCONsodNKxN3a66/VUmBL0MUiWT3SF39+/aX7AI9X5RJ1cIcpnRMRFvOwBDgtdwGD
5qGUklgYQRl9gpcYqGbFSWKVEDKsogSS5qSNWDN84rpDWKtqY+MmH4mdd+pKiXVf4jP0g23vkWsF
9gZKwqmPBfxcxixWa4ReXC0b9Ts1db0n9EORsQV5Y5+Wceon0CFj6XtYFF4hdkWea9N2F+kKa4rT
e01zWd61wP1SSh5K0zl+H45qRC4f7eycRKCrEn89EpJN74GlLBu9Ee0uS1BA78zvviZH0X6m5Kc3
Ci6RFSfJrT4Wpp9v6V1UeVzuHaoHzXBd3yKpwBtgAXjThXGmFuZHmvQ2Hazvfz40QOfS9DNcvRj/
xmPP6vJTA6JV93VNJXO2Qd0pK7m3UPIvhywN42c1vApotxeJPSa/0KvecjooyCwEzbPbla0Sp0Dh
lRjHpbu2bR5j4j8CdDq5B8qOjH+z2In64kNquKES6gcneY6Nxb9x6fKuA6kOAlh2X3hP5dtzDX/i
6D1MUdQ7TRGMvNFtBIsTzlX6d/jZmd+t07SYvvmF86N+ZKSx4nb2T7mJlCBz+Zio3vNv6IGbhMQJ
dxml2E/2EKlRsTdP4HNYq/QuhJ4o89mEUko1nnfW3BQslkLxx0ONv4fUbwHwhgrc4BFv9/NtiIyS
7q2b+LOjDUfzm+oTXpXLTjTvkaUcf3agmSQlTwvO947zmdyDhwzoQUqehkYh/6JD+/9VNwJZmdXY
4S+TrHxW16iWa1MHrBvk5iyMFWzm/g1uDJJixjgVbgoUYEDAyfvDX3izNv5Ts8pdMA6z/gwudLxx
/NEV7bSRScuVFH+OaZoCnSql7w8nE3pGsNxcn2vdX2x2B4sTPPHcEyYs74nl0XPAeG6AgNua1ohr
dCxiPBbfjzOb3dBDpEpnT0VIK4Wn5FZvtaaZVx9uTWeQQCqfuyD3zgLEfsXkJQ8Q8SozuvWPpqAD
dC3w6uZXd/WQvTusdyxJM+f+Lv3GIQKBcd5JJGBP4g0q2PS86QnmPWPVilskMVLh6Lj1ydiFXex8
j8vDEQc9d1XgkkQIaDLqwUyJZQEtrlRA0QCLNnFIVKhwqQBqkwpV/ET1SKOCenZYJS/0TyeF1xjl
W1mwyDdbq42dl0R9C1+0q9R/hJIEGzpjLEh4FBH+0au70H0YqqQ6SIGfe8E6cxs7zS0ZRRpgGlDL
OV/axD4kLCvi21cKxtAhrocGmWjqN+qDSGTQd4/Nhu1a+EVnnMbZCGKvdTiumHosIigQi3mwRclz
P2s9XG3rHp6nS34lJHf2F1M/NEKnYvDfBO3rZR2PEXBai9OJPT0BC0PbMezM897PsLxkFUPIA6vw
lmQk5BqAn84Oz00hkiIi5sXPN8/w84VDEBsaf7562WHhB3PCEzYT21FJ35bRQMmQX3tNk/pThstC
ECI2mcXomBrpAD4bXeElF89+PXhKrmAGM3QdLKD4GjwbmnPZR7jBiIY5JvLtq5zInOu19+LfavId
uXHQwLxOUe0bPs9NfQZX2UUTZheIkmk29x83+a3YkfYvOgT6N2l1GiFLuNkD04KnVp2HdxkZ22ny
86OmeR5pJ5SZohOypOEGoAm8F5O8NgAtxOhOzRpAoTLc8FDCnVDqGyQBM0ReBFuAmxTFXl4WEhZJ
jpTQVwy7PoyeN+QS34MEBcMXnoCgyqsAm1lUbybnRi0CQmIR58UB5gt9kcl8RbeDhC6F35I1+zcn
b4htSNCZLkcg61fi1uG2hFYYePQVW1MdCePJvSnjdA8RucsJmVN93Haq39eFPqUrgdUtKIDNLiJs
vbcoyRvAwjqi/so0QpDI08PdpgJ1QDWJBWyS7qJltKW1QzuW8qR2olgLIRN3JDuLFCLgAaPlmL7r
u+7rNldUHd4fF4+u9gga2OQtI+pOwl6SB23TPH37r6lbPyENnTS1MYP9pAw5zIo/9jtvhZXqFR97
3YOpxlXRup6bBM228waL+CWbO1448IwxXuNLzbR8tMlmdznLl9lXXSjKZyQAubpan6mrSmXr6qRf
1cm/K7DDsEsAhxR+CZTYK5DFkfUklGxQ2l+zGJbS5ECBRCTA3wTR3NGirhEkKhq82Q9GUkYMZiX5
40/G6HM1Fa68glrQHSeuI3hlfhKroiKBYxbtZ1S3SL4+AblOt9Ui7Zgt2HSVO6kh9vX60PFrLWXy
4q83C2HdY20b+6fRC5JNEIEi2XO33MFHjl+KOP85OGy+RfnalqFj982MvgtgTobXF9qxjvgIMiXr
cXZaVNNxTom89/fgmIF7sVU77ChjRUn2plWS4ylcClgpb1ILuBh7mW8cB3BbqHj57XNe7ldv25xK
c5u0mbNVxKKyU49p3htzEhsmCgpCXZrnodBmowksgIPjL6hwHSjflWLV63SINVlGnbPF2190CQnw
Hj9D3C1X0zbxxod3YPPG7+bIHKdOabBc66e3uqmo8jUqQxsoKMFrCj8Q8RVll5ljhHj9IRqg4K4h
Kw6tcyGIAwFhhXnvGopCyDRl0qyfZxbvfYoZobusg83SJFKZPSPRn0lCSft5d3qkkwx3DtzDW5QG
2NoCSTchhtxlbZaUXK5rmTP8IyHfIgK5pW72kR9ZDWPeie3LFwl6FzkwNPqQrmke5aU/t97wNiZy
2FeF5B5yu7I12DXGrj2F+tzSAQdCghcvVae3wsgyu0amRFGKChrPble66T2MoXXiWehtS69m8RZl
PiZ24PjRpJ2aI4R5smXf29fooP8Rk4DX1uaCOpKD+5DZSj9prh3CAr9aarNWnfqsFM2HNeBXpqm9
Kb3taby/3Aq+qrTSdYrT6b6YAKwuXuuEbeqt/Q7thJ4/Ysi0hm0rTWazw1ZHjyaX0XLfUPuDgSX1
P09T6ckiBSUR1wO8QIcnMWg9+mLokcdWpe04LL7ROXwxYhKqsRmChK1TXPwqjgh8wMb+5TbxupB1
LrkrBg4kLoX5eJKOktHokFw8BL0khGmXtoSS7FIcyCWXWN9fFTHgyjx1MomUfxfw42x0KafWV9YC
O0s+svljlfPVSUrGwYYU3VkbeyhH0BBfEbL45kl74Y8JdzrM/3mVxO9Yp9SUG68ZyrCOqoj6pKvj
U+U4Jovie+aL1KLeK9tGYYFPjzULxad2K1L04biFbhrlegxp/o2zlbmGKrnqNywwWuKX+sZ/7NSU
5W1bW5T7sbGi+mAoZaaB0e7GkEPZVWg87GO+Qmy40XYYOuiuV9f7bY0mW/uV7d2Kt6RNAOwCYH4i
b8bPJZ00Xw8ZyJJaGXtOmI3lLLS95Q7dIrkUEsQJokIaBckIkGerrHTxsvaLaafc7yGW5eSrnCTt
ZRHC01mgS+8D0EBMk+UIRcmFtk59BSFzPInSGca9ToL0OXRNlthy9XOQ8nNmgMZyi4zQDRZUlxbS
sFJKG4K74WsY/zO1d0m6+5t7tyvsr0mWmqci972Vb+975sy7f0QJB12YxsV9SCwvGGJ6P6914oqC
DtugDJ/EbPZepzpupkZ7jlXnl3jwXw/XESKKOMiVzaQRU9iBCdM3rBi8ekdBVDd6nFUo5RfW3zGt
RRgvbieUw+VqjteWlwOOXHmEl6mPQUadtR6S5Q0zxkjldcCtnAks1iyGRe0kF2lWsEkeFkXdMApw
PKnh8mwomkH4ii9YyQjLXMt7hJfrgk209gPl5wch/9gCDZqF7TxpEdjHNP54xtq5eFkJgaBR+Kbu
F/9WU6PmZs28XzOMLC/SoOVCb7T/4RseG53HbeCz7/hDvazFS+3IdoF73niBnJdw6THNRRW+wlVJ
OJ18p8hyfY3KjL/XOyk5yYmGiyoRJlkm5Zb2vzAUJsV+vi+brUJpit3aI0hBuhx/usxobMrQqp3V
aMcbdUoKLLzzTQsfNQ/DQZkFmSYicEnYpfa1rMOPFO56tlzCwNc0Zhca3+Q1b2r1C18RY4NyDZSM
A290wAddG3t9FocBrU1YqhVcUOoLzf2RYuCMtBGkIVfaM3gT/YcbrNsoPVLFAoljB2IxXiNG5/6J
/8k5x+CtNC4huh7AsrLzb8QxZqzBP6uXoKMx2Plka/9Vd10YWyw0n4k9JAI6pRSjTnBg2cAAsgKa
rOtRqthCDu9bsdQEdifQ/x1Ld2ZRaOce8cFBLOCxqBozeUnc9D/rK0cA5F1hkZCA74jaUtmv3KiA
vLqx2YCe2zN5p6ww80koqHuqjhE7afaiMOEqfgqH56vdNZBmWLXO4EiHwlZWBjmYv5LeP6m8H0QR
X5snPnFK/Q9eUxiscm5rrCq3ymDD7mEFOYk4IkmPyVl9ibVQYpoiWgzFqlWMtX5vRHbiXP/jV9cR
DOu3FVJFkJ95GpzRK5hZNfQKzt+aZ0GDh7LLfs+IrCO2vVBOQDjNjC9ghCLljebtepzSJ4mQoNCF
4ReeDhex7F60nm3MDulJD+DVmPOdMPXqOvUfa1xL7gZu8AKF4YS9w//IqmGZZz6Ac1Goi/saAd+D
P1lf5N6tF8rbZbV77WwjawKIgspjjbp9+mag/r7gRbodAXaAgzVrqxVOVs1SdhILKdix2XFa4TKf
Rz/UEIxdyJwBxtzRFtrzz6EUZ54DwMy2P1NHU74bkNYJgQ9kCo6NksAjQe5Bf715q6uzFlgKFFSR
f47iZ0inGbBytJ6x1x0zVGGqktlWFTDiR9CLWw3D0n1zLWbee8Gdl8tLefbg/d85p4LCplAoeeaR
ctghHfJc7Za5eRXsdjQKd6zIOiCMxvu4nRo9wW38OpkIBEzCnzNstDCCwkBdc+7bQZfVc+ocqa2w
pVOQmqJxB+N2daejNQ/cHmfdz+rkDHX74FAnlkISpqVhqgHtwdFJH6sXP3KhPQsB0pHhbOuhvH+E
OaBTLWdZHo8WVxsAsKk6bidqFkodHsB3nSH/iuzJpwSKgb31JPGxYC3VHMNrADdvC/q5c/5aiUXo
pjfWTjMtoc3nNyAx8Lh6KlWGtr2S8XAjdX/Zg90d1qSkT1xkyQeYhaFBVLxB4TJEvDtGNx48/6gs
E5kkl1bDUWOLNRkeBG6Lk+JtpsEgLmxXnqG+FP1+8/Wf/jGFejOgicALa63AU9IbAq20Lwnkg0du
ALHzZb6dZifaipwTEeMIvyq+UoqN0/vNtUyQbsDv5R2JItqEWVXHYZxmBy8XVZnYNtW4/1bmrIqe
Zs5hqTqY7Xd5I3EZ5/yAivKPPY4NNmY4NPLT3hhwjNIRpLSSbCy+1y1JYQzXFuoAUqc8HxUMPVxO
dO7SOTO9rJ4r9AFQFp3mBDJnOTd1vU30EFka3NtL/hbEmAwgYFxfCk85zp9lKf80ispsM3Q9VUpj
fGvprCusibr/lSdJXzVteHVA/H4LShg9NLFCpbC+vKMmS2OOBTe65rFhvm8Lhu9sKKG32C0WYASM
6oXKGhOdqgark23s5goy8Lq2L2zbHaYSINRGCKmsx6+lQpgAefGu3QdKDWvSquKZFPlvF4dtrNRJ
/ls5k/1NxMUvKgLeTkoU502xTKMbNihxQUh+CSSSfad0/yz7cKwDApZTrNqbbRsOJDK9F4pQZD/i
eW2d0xAo40/i9GH1UWpf9jbniAoLAAZ2eFYjoXUJ5xn6uAowxEHZZLX+AjXODHEbg1N7CFdJnuOy
6w7l/kNjnIJQjysMffVZFAextynLzGaOcLPj07Ut1qpj4WaCgUhnPqdcIjcRww2yu1q8h8FWTgis
Ih7ahLa5vMLyVMcqRc+I8d3eQMDUDp3HyyjKT0LqUtcmV3lb6/GDkZwqbsNyxTyFXYiFUpu7xgT+
fjPeEpuZSaoJ33T7KBpk37KE2QiR/GZGvFHck9vXG3GTZIeDjl06JiQ7ARECiscv5R2BZSk3QD4i
YDCvTyfjxQEB7YcYqwc21pMixo0YuU7smDQfkEuSBMj44GauIm5AaRAUaoYKJ95i+z/31hzkerOt
tHdxu0CgehO54M3kwlGch0s4lOeRS2X0K25R6VGBk0RG9PCHdtuPy3zz+/bCwG2Gmak6TkWmd/EX
8R+98UYfZaI4weexnCUguyu4VDvtV1fcbypbpPihrNjhEXL7ydQKSpLeuXyEXtjk18AhNaj1pABX
WUYmueKHAM8bnvZUMlM3ch6ck6ZbNMRn2VhGXWqVEjKJDjIILzFqM+oRFofNGGeBtuMjqWs+NC9/
BruBRYcYhmsiyU/8vKnbfs/q2ruuLV/xEwK671O2QHZQKst6/e62wy7FeQ+4EO9Q3EKVnXjjM7fu
ae8BGVJlS1x92cXKiFWL8vKWxSP6AxyYiUptRFZEaH5tQf1Wsp3gVfwR4V3AOcDM2XA0Wf4M1+Fa
17ww4zKLgAFZHODWq7BI1N3uOPWNGr6r58t1EP9LN4zzTzc6e0rBvq1qQOhiQGaVgBw6k37Qv+Ld
IDVLCjFr5Db102+P+dKubKIPnmNigI5rK2S5glhmzmqxAUF0HOzZumF7TBHMDMIxMzYU/C+ZEvLp
jDMaiPzoP6kfVDUEbjbGdmGOFP8eSFOBuFpN/HvQ0mdcEy1ASnrDs5cwI62U5TZ9Gm/XC9WrwFlp
tIwFmZTOJ2AMk4QxcO84MSYRY6SdsehOE0RMpX40YD8hzQW0WqqFq3ZAZntPxwz8qzus3QblUEgB
BvD02/2u7FhIimvC5g7txmzuT7LtOBa6LM8L5+NPpv7za8YrWWQpzh+0WeEOGMYsjMxCR1KIhNm7
uzM88+6p+9UP/zoZLE/mbxTTf3z4UImoSUSs2NAXT9XyeNH5q86h4qh+eA7GwRAxLuk5hg5wdgCp
k935TyeTxL3az9LXjgsuv6R7uvDxIIswYPRcMSUPPWz8Eyg98D5RY0/R+RxzmsTr/pvodrz919GJ
VP+nzhm6twDmvQOyVcebpB2Ax7NcY9Lcn0lhX7Wll2vaS7eApwYD6QQ5hhWS2S0bwTQC5JzYfzBQ
W7AcP5xgP3ASI+nBNc53v0YHLJydNUAk355EtnhJlFIeSHWx7DCCw8lKJaMBR0o9+Xt99M58czJc
fVreRB+Gx/XrqqmmswyyGCYyS3xsyAlzhn3G7ZsLxmIEM8Fz7btj15yrm544Rg/onxP1vhbo2PiJ
r+vkKeXW5WL15mkRu7rSPxb4j5FflbqmYMVSwgt4XZ5d0YJNogfx3iSj0fDbcua507Ti5tmPsaRl
KE9VO667eDT9QA3iKKEKjjvLWcvGEakDmv+2fGD8a1XaNb15FNsWdvu9gKG8Mbb66ytHXZmXDst6
4dySfxLsKfH/fj7IgFU1xhVMb16t21oqrKe026F1Rv2Kmbrcx0ZS+95oYnhBN0xp/P26P/4xtDAx
iENtq+R3M1o8eTb6qJzkPUYj78MBPSRKxDJ9qx6EJ0hSkEOrEM6RyiEwaJHEUZTbNGhB4GIeNPXm
WdHcem8FMIeuSkQ6O0iEWARPaRtjDMTn20DRly2da0WQ4kFNSkHErfllCD7SAf4c9jzYSAxg1fBD
bjWDddx5WzZxfQfquemniTXyHkO7P6B2xyHLLFiYoPZ++Myr+CX11hgYpgRf9d+qF7fe3bG2FSzc
6GgViZgShD+sFQhgzmHMkVSlq4Px2Owg9eLtRC8XBljFUtCPqFAWDPuMO+I4mgZ9mgPbvo0n0ag1
3eUUI2rMtQ/b78sg3PVO37o+c19oy62ON1OVu+JoWreYGTJFH1mfWAYTKVOXq8B+jIxWLIFcEo+e
toOpAOQL2u3FwPj+HjOq29LLSFxS+MmNqb0FQ78MUv43fzpUevoYerpEcI6ReigEd1Px4ANtI5An
qlsyis3RIFxugLIPTKjcvw2mUmiZfmG8uafRzDfvrs1fXDBi41/gL7p1ZM081iHTjRPc81SEZaNO
hmq1y21+bUp2s4ecjO0Kf03PA89qEQQUy1CcV/xcXeRFeqOH53XBU4Uut6rDm5xRCbTxoPB1xnYB
3w1WUMOaYq/s6ijDxAN2PzEAHYVzOy1bSbsB5azvWkWfqxtOT4LjUY4VTBci81Z0tVmz7b5onzFx
ax7KFZs/ptADWuAs3CZdYCsDy145593V8D4G5gJbV7UQ/XIhUmC4CFZU8052UGI2ieQE92Ri9e2g
YG1vj9O/IX4HMsIQDzLsKnH2hz5GL7bs44nirQ5pMWRNunCUeECz50QBDeE0ovMOCOVr3vGIB4BT
lQpaE1aUXJTFYu7Qt+DfGEIAtnkaGhtlw8e2rJ8KZCf/AJymRmiRmM1fnnpMSxTBt+s9ED88AXt6
TSP4LQGot5zmG3w6JRcbwMJTXBU7MxpW+cFLxa3nvgGHvV1ePmlvL50FjrCcySwXPCkDnAWCSoIU
vMa383QuqWNJ/rwNleisa3AlB9i+nxkZsY1L02TiIHWnQWGx2QLh3BupBkUHpy7HgwcEqbbdBpS5
XW0Z0oKFsmawLkY+zeatyatOqvX17AAKi/5TA+jSlb5UyHGUQdVfM4mujIVlB/saLDIL3xfbg/uh
35+juyTK9BgCDsHLdgZ3N6oDgXUyYYrD74OyJjahogS72FqD1ScKGw+uzvnkflyt5bF5Jwjf0nmK
CFqSM+H8yEJL3RHoPsTyOrWbuTJJhT4TdgpMcSNnUfi5HSEjT5p1kcPqSKk1BMf5M9t/u22C/zFs
tBqIfcAi4Xiv7wv7p4bk/fORwfv4xEhmOX0GDsKsQY0P45y8gg00/w0wIyLmJydUD+vl9aaeooTR
+IdBNCISCbm2s4wtdp639n9TMO+pQGqf4i0Nj4klaqrg+4azpM4ptqFiFXBjfC0zsZF/giZecSfa
ev9mwyDeAihGyIGukSdgkC7Tpojkdsdnm3adsLihQ6XyupTinQE34SCq6T105WYAFEZr7sMT5+Nt
psnGh/zuFx94wmSHx8guB+TEp5QM8606uljPWxMJgFNJUo5S7uSbvQBd3Ldg4kxjl3ki0sF6FprJ
uG8yS3drtJB7Uc/8Cb+GkhlAR0LvtJb2RoOOs9pKpbIpbwWySnjh/VSA+MasC7n682ncd4ZFesF5
Dbxm3AUvj3gQobw6tY1ogtC0GwyG6zuiN02u1+bBRbQgUwo2ZPERKSWXQKWzSZ8xm1v9Jf9u3Vl6
uNyAEOzrtkx7Jy/XQnyHf4T6sUlRRYr9DYmJbRWN8RObVGZ1BVWmfV0CDH1IaPCtuSLMn+Q3e9E0
oxMQr4kuzzXf9iNRQm/RAanQI/MGjGoS0MFKE9TnzQUXKP/VBITtjUt72bNhx8JI7ai3lw4KiXMK
ZcRcdWixpGIsBnNkALDdiHlOulISrBBYGYCpiY+0VBVJlbYK4ua6/nqXdGzKaeOHFiYjyunlsDfy
JKqSxKG7okrH2oIVkyWwk5lgiPEbixrZdRARHMQet9wb/Fo29f01Y0ww9nGmilN4f9xv1UiHjZaw
we10JNh7yxylJp2Lhm8eRzOto2Xh7xYXcyY8wo3NGCKDw6olYLfpc5qyDHQn+WInvMmX2YcnRiFz
E+nC+vlERaaPNvYIVRYkQun1i45aW50a5tbNZ8zhxE1NFGRkY9gd7MD0pdmUDyBlP+DU9eRr6qsW
gHquRRut1OP49v3QuObftz1CWWPCQIBxMmLXysclCmGoMlq6qjdV55owxdnzel035xM4vrFXRm4W
rP22yhB8g6rwhiYXAgEYRWF4LoMU7YxHjnXOjT8OOmdPF+FyZPUWvoMXSVY/c6nkQvKpwAKv0LYu
svvc3zr41xA8RPOZkIL7NtfTLVIpQnOkte+8fuX0jlHpT3diObmzxf99vQUmMC1MEhe0eCZdm3At
rQX654hVnt+C3r3w4dnjh+Z139K4XMjm5Xc3+e1wdBJTWxg3+406lfChk/IadB98yfuZSdMlsrKi
rouCTptTtRolf0a2BV6HCYM0frNlKZxg3G+fcr82AfDg4wyPBuxgkwujPfR2LVPPQSFaXhgbHD8Y
fAoVZZLWKtwIvpbC5756OXleJWZWWRn7tp8qWTKzbjZZY3B+KyyDXm9gsJktJdhTFGpoTF4Bk9K7
IoeE1KWKUi+bZUpkJC0f06qpwE3iU8P/We/bGdF73rBRoJbbUhUNANMjl4tNydxj4r7bNKnCT/c4
Apn58U/8t9w7jnxEDVldpStIC+5xnKzlTWepip0Y7JK+BNHYWx0PYGJ2Jtb40IMaUWApyB742NV3
KxU+Qsy6+16PYM0en6nw9V69MF39vyPjSVlbWsKsbFmLcyvmMII9ruCKI+hsETXna8UKUgu5+aLH
f7fKDriyeeCWX3IaJ/IFTPfpbJEhoqrz0UtVNSy2otgR4qJtF131Z41N6PlKnyCKbWTCS1sA0MdA
cUkTYs8zvpdGYt9ioubTuNnlUtWOiLeWQTqTLsPV8Kv6kewA0tUyOyZ5VG8Vy6hObWmuSq5Dp7rI
4RH1MY2DDvk4KtlK5SFiicwyzrWKI1FYyCaLvkwvK9vYRRWoWL/lHmeo5IX1z+7d/vT4zd7hyEzG
WTMlKpmeSu3v52bMOVehwTTfVGupdY2KnRk5bL9oLoEjc45EPRi1XBz2MOQBQmbU4NO2K0jTJJv1
lIxeEVz/rJ2biDv6fQGIAqHrPyQbKNf/1sWWKZjkv7lXoVPAmiJJloAQQdpuNu5NOnqsJPM1dvaT
xt5McEpsGD95tRNNlsyBCvSYlp+Tagr6ANy6F9huNXlITLm4nyWKwTAKW+Q0smoCK99VjEEFpWG+
P/4w6pWyygRPTGqt1/nFEmG1F5g66T2+iHECseHLp0MWvDCiYV/heIIbdltLLqUKFOsw0Oow2gd6
JAe3LKlI7QBtr/CFam88G8t3lZXmmn+bcwJYvzeUcY9Atb1v22TVfZ0W1+5nAx7lZ7Rk0KkueWuc
RCpbvgK3c4NkCJq4V6KgeYb8LceweoVosgJKg2cV/Q3HtVXX1Ds5xslCj2rXT2Br5DaGtK2xjcZx
Z70b+W5MyGvwpmx/KuITt0dp4K9QqZVOHyLmy2wUPlFIKgNsP8kUCHBvD+bO2ZPtvObNCGPsMtVS
f2N+ETSQFtmra/S5J0SPE1WOXp01YrC44859vKzvlZm5gzyZeeKW/PiUb7x/fkeq9035STO9ppVu
EdhzctB3nEf0LIZ3cdSlFbMxe50P6WLFeKUvD+KAf/66eMAPOhPEOFDfKgNUGKPucakIBFdcnmLr
7sKO54iV08AUAB7y9C1HrxMQXAeJaRtSqiXUhsA4k29lJW9mfjcjBh/w5VOikpJQlRKB9iArKzyD
xcitEBEa7MolsyD7Faz8Mdq4nv2DT9aiER+3DxsrkF4P5jNusbB/2nM/X+de/4gw51YrcTAR16Wl
MvScI1ks678MxGBG7YLGjLUZHKmDgTEKQRxoHK5O2ls0qcVahuBS/wP9tEviRiua0wQD+VWpBaRU
5ShDv96N/uNFugqQno3A6osJPnWoSZv1rPbjKLIEwIdBG5BhUKkRLghaTBvzZpiNSOLUCRMxCbI9
rRAEi/EP1Kxk8y+Fz5V5FxgiuY+Pqo1ho+BeBn7VzcoSsjgZhXiBFOyK0/Q3tvLbAzF64HmMHpcA
k4wH72cV0PUUoUHa9v4BzRswQ3AZ0C+tsNgFhcPHVOyqgSbBc0pUga3JEJBV1Ttg9F0XiTva62nB
S0FqlqdS+kCtAV7Qk2ZnAfoQSsssa92VF05tvhPcyMif7mD2N/4qNgMJ9T4QL5QNpVBrdjKps1kb
AuLFWKNnAOKIsj/qlDWGMDM/1dLBXZNhf1GSZq57XyTR13ZWBJsELky6Qn7Ufjh8X4IokYkppP5y
725oDEcsP9V8jZByQHyftNBrhhN8gZP4aS2TYB1IpshHnVhN9jTuuMVd/cXh3QGWIJrIwgcouIcO
G8AeLLaUAtGPt5p6AUbA2DVHJyXjlWYscs0G1OKAmSO2kHMNDpPv3yOpp5Gxg9GU27XZFoKBotWc
R9PXpnWyWqbPYqseU41YwWZBw3/S8X7QvTMyQq+KVYFIwDyBDVArTU+XN2ChbzTQw3TrKYJbQid9
VRbyRQetczaqW29qcsmVOS/OH4bcdL2/eqViwN5pznzEsZ/mowpw87qXCJ8d7Il/S3nUhfQ4x6Yy
mRwzp33FqbdnaR3sIvhD9xxcWCNBqyTnSRhi8UQqitbM7LxtRh7O7RgfmQexGcJ8YkOl8g361GR7
kTTRWgAvwY8FWg89cKP3pNKCsrZ+GZnG6bb7m05VG/UPzomreerypW9voc9v+rtuBwX2NccIPWyR
qNUM7+ZXS8Xg+GHThEbmWxVtKbtRrJACPZTPfpO2XxiUYku8AV7MtlHeCvIzWN4Jcdo70o6QS9Yq
CN6liMeS16UYkNnad5vkQNZji287MSKWGgkiYDK03ftPbAxzpBal3XuVP2Ga26QQgcm2qhG3lRNk
Xwky5REUn91GIQaaTcMdFevyx3tE4FzN9lHRKcNqO7W+VEjqqHkv9iCJmY9KN0eANtwTiPX0VFP+
fnohVIJEYHEkyF5cxEsNqgXMUwhwtDo91MHPlWty5GlUIGACsLb/QiBbNpALEM4sfytNBsFriU14
U8jiebCRL+/nnvfTXvf4G2x2v87LR2aSruew/o/4BM420RnyM4glPFPxBTXOhPYKJHL1Gmn9JKUa
8eJznuwdfdKwkr2I8v8UnCJMJlwelCS0D1rZZE3YTZNA9NHz4YrlaLPCNZDxBzXYY5OQGDwbd7+5
lit/RVSWopQavxcqCgDKFzaSHwiLqUR+U17PVb8Ta2HhKv5jZAYhA6VgOBuU4Ylx0aUk3OxfvtA6
iX75iRR9AzL9008c9JgWBnH+yIq29ssYd7ncdZPYzzcH8cvXsFdvJ88cRQ9hyDiHeWyVxpQbeFLE
LeBaM6M3jP9TIStjlciDNH8Sd4dXVT6VTFuU7l21CvF0L+gXZfG564FLCEAWHzX7a0Mdef97ZWD9
TTkZB+6L0keyo73eBbvfDH3QsAh31eRywhuyFp7yMXR5cYsc/0O1Dz/eSfuq0R4Cw89smXzJEP+p
tF7DT1P9Hay+4H+EngFZe5t09/OAa3tyDYKfjr6EaP3xj1nt6dLjlWONBCD64e4JSBlPGlTNM2Zj
tmZ1nicBGXSwpZqLmt7QR2iAwlDqtZifM1Xkuj0EeXd+YiClg5BUrnwK3DRgqXi6TY4pRKR4FbYj
deB+I8PnpzLojqjy38LW1TWc/WBG63ghq4MdRavS1XQdzOnC0Tpak00U071GdOfyIPRCp85a/7kM
cNi11ZhxWp+Cs86ZjGbyxotW1Va8xc5j7q2K34qLGtJ+SsmtweiWOzQW3BWcMylsv8Hw3ddLs0Wo
zChCtA+4Rm9Tmp6OxHG7f21t6Rh0qf9KlKe9RpJxL5HrhAVxphddDxlf3b2KVPbYKd16mKNDyaSe
w/TLVPjgPOgn8TlE8aNe0EUOU9FJgc049gg1IlTHe1NrNHbh1sq4JnQpCiiYvRAAgKqp0n1It7NQ
iirAaRfBRzCnNs5EBYCBojzIUlAGuHkjI7iKWW7jKDZT44yxztTe9K7fAA9aDgQEtLts1NZeuDxq
wKRUN65eTcgz97Nb9ivVWKaPS0vt0uYOcdAM26C7MLcRIkQ02FqoiyeShCTFZLj02PRVPqK0vPfA
BP3taH6kQP0ZOCWypPrqCclOqt7sD4jAlfJ4kYhgRHVTXHHEH2nk+XHUW3FsnTAfZZGjbh16FXED
5rEGM9Dy/xvEMraZJQ8PAp+koXq0iNdN+3NUd22zYWxLQ1usNGfWVDSX/3t4lNkDIxq1LHBS4f/m
+yYUHuGWraLYZufCBg8ZQdseZ0suuv7VISZgRzlVo2saoJZvP4VpvSwLpUzNMsWhj7tFE0gzJjNr
QOI5hNzx/YRuwfQQ6rOh6DYKi+53AmL/ESE0hB15ZGV5RNvZ4+BUCytoS76qrVKh9K00H840l5bd
1vd0kluRZuuviEK0Cblx2XzzghzOxrub45sG6tjDwKgvpAQANErZEQ1PmoVJ6xbYoUNyIgTo83Ys
ofSU1EsXYfTWn1BXjvMGJ9L8LuSUzTeX5XuQSGu1MqmLkqezZXLk/+f+eYvIuCT04yVavDsfzUJq
p8nRnQZmdEqsq9ILU/wfGb4iAM2l2K5JvkToVLrjkiF2ejZI4OKDNHxQaZE9fUZUfKbthBc9XbX3
/9cwoiKQMKDLeeKwo6nSVdEm4acOg/aqjCYsd0Du9W+uaNv+Qkqi+Gm6178cW2HXgjNPwuFCQ2Pd
BWr529wzzwiaX++E+O5tOnyXak7qWdaFpEA7ghcEDXll+ss1os+Sxb2geUq52mP4rAUcvtPkEaDA
KaAo54RSODbqTmgbW4NK9+e3CVTLHnOFgD+M0lC5YGhTN60Ic6O3LpSZnhHFpSMyh1a59/yFvF5E
8H+6i5pWPzB9a1v/XRm+DhOSHeob8xz6dtdHchaCYtza4NbB515Gtan5at6aUq5R/xDgdg28ZiH3
8siyum26j+g52LtUoA2rysbojxeG8mglia5dfkoQqFSrsvfdyXHx0dsw0IbKWoRsUMR5CSUaZ/Ls
FKvML3wf7P6mftfMHES2o28PpFyERDYM0EG/jcrPyU7AwlmDPulbKznXHV9lWUC6uHSv3Jk4hInS
nA6wKDJn49k/yAS4iJ3v4HZlC3TNg2QMnXZhT+MA8NutQPGw8NfbCg7t8VRUWlXDy5Rf/JAGohWN
xJDY313LLbwokpCFiK5/c4zpLjST0mrXFLfeU2TSLHq0WlVQM73bfQajD2QIeXd02aTqTp+vK69E
ZiZ32yLstjL+nCHkG3XKkSYq2NtZRn9UxzM06c6gGwKhi8XinNIe4kERm9FV/H3RUgnhn6OMb0ld
CD4yMuZZXJ5myZvkc2D0TMhQbpRjeK7cty75WBfJSOEUv1PM89kUyhPlfDGgJ3tWznvJpA1VK0KY
9zobCWQTPPq8WogXzbV7Q/eQlwXSNyy9YZomhISNYmosOV7FeFMy2XaMhQDwR/sNRkwlSFTzoe16
y6+DIIBFFATRzb5FAVwrshyovlTDNFOt7nL+Lg3wCM1HGgZ6KruHHqMGxk/R/mMyLoIpnKA/pgvo
1V/ZIEzv0ulUpGs+RAR4BFEhOsHGJVstV78/+QSuJJ6U7RNuS8jsnOSHzb8fBtZKirQzCjqrjrf9
VTEcVWam/05XiRGIGpgg6nc84XU0Rb0iBRRN2KNO2Ows5BELeaSMlF0EVQwZkGVWRezW23UK6jBw
9GJdJpH8zQCM7GFj4lI+VdbqXla+pX2OiujIqLKsVCL5rC42f0UA1bSNDLfkknWXXzWPgFB3Dnmd
yIuLC4al22aoXAts9qYkgjPxapMy12yuyMOvaLirALJDqLAySgdx+KrIEuVAQ+JxgCRXKAXySuW0
pPEZzrCqsswT67fII4YsQ3p/XkDyZ73t2UyrI9FeXdZ7TkIPJdodgyj4MwAUZLE2Wblwla4Ab/L9
PmMN47rEw3t95vQPpK9I+aVOZqwbcQfO/LbBBAzUlAFgoHeU44MADHm92dh0PPXXIXSAfvU/yDse
4ay+2+dnOE6a9JV3qioFee/Nw4Hi4rk/pvc+GOESy3PR7C10Muc2Np39DZv4yCBVTAn4JhxvE0n5
+Ga0R+rBR32qywDFvX2uBbvVzWb5jto9cuc7She+N6uoOlbBONB1Nt2Q/Vdf/GxTUmsG4vsRQRv7
Sv4zvd+HhtsLKJpvlYFkTdyr1THv45eGPeNR6u/M7esF9XmkgHIBCWLNbh7mbwqTgR7XQKjKXQMn
C5wHNjX6MkCqT51o+vQ8sCu4w8kjLJ1cp183cFNUq3CZfZ2Is3rvxvChS9trJS3x1Ph/bS1yqQyL
wr4uXYF2tw/ZLB8+dBqR/RkdsWmcy2vXnkISRcyhI0JD1Zn7Hnu7x5iuIBt2XSBVGoQ4g/0EwZl0
qgdfuRrxRuIAoczIbnc81Bh2fOSHQVXYc9FujT35MszB3o7xdxWfj6mwzdfmQogmvhWg1obQb6a2
ScMpHNaW0J2QyIo/X4pWpP+bN4bVto79gBFENIX1n3fcTNUiwIcH5T3QReS59mCFwWIbLz6NaUIX
Qy6xi1S8GUUdf1UJLgzZKWnKOKfli38fvllir8iFl3k6NAkfr9I1bpmifBATIS6doj+nk/01fpHP
K1x5EzY+DL8GOrw15LgFQzK9FB39DhWdZauJAdt39Ode1MFBUHn1VOMx3XDaTkPBjwZV+g1NKQdW
TGe9GAbups8R7ykmiuT/Y/iDC04XEaqz25n4py2sJOvqOjQBAj95vtGtTzWO53cQ2Vz3NusGijgc
Dl7qPc2ddxJ5+yDQG1PjK+VLAuco2TIigkPwXNVo5yv62w5Do/xSdP/w6+qBYFuWvIXaCpLW1wrQ
W3Bj71ocNNrIu1IT8q8n6wPFs7RHJak3ABEwBSOsxZqU2AsWnAZCvlICaeAJAcm5HkQttGkxfhYc
R2hoGXQHmGnSkkYfKmzq0Br8CcPSS2pHh16v/LwBbY1MOXRpkCapR2eOLyPzOJ+ONblRfLiLQfMv
gnzDfMmM7vfOm2DhgrSUa4H0She28Q2Vn/jsW+vp4y2mc2RxFKT7BHJSofV30keaUO8sEEKln0Ei
TYknhF+p4bT/xOkcdjVTtgWM55uWOvGSfAUZVKct5q86QS0y/eorQDGarkRDdd1+92aQTDNZdK2Q
VTO3pMcRT1bQzFEazUco06mEWS4u6qIHd9umlBaOhglbrdjxv8lelM9XgNLJszVKwpL3QYRiRRTu
2e8M/O74YQTKD+8E6S9vXJRN0Z4GFsmazSu7B6DI92Z+BvzthMFxlZXU7hV0k2CojrOfa91XImov
Y+PcDE+Z2PaK/uv8/Aeoz2FfkeunEiEs7zcmqdfp3fAPOVSlUE7ux65SljqDvmGsXO/1GfUJEwRr
R5TDjrF3iV3W8azP5dCpRz7BhMbu6yHNK7THE9fzqiinVkZxIVN+TUms9J30doTHLh6OtNuscreW
O6ooMEsj0tNm/D2hDCXLK9ytHC0F/pB0o0B54vf6EFQDWeSOW1EYg54ec+qIxYdmnG1n30pVgMVL
Uc8WWhnJ3WzgvY50GumLK/Gttbmsyvd9FM+aICJPrm1cY6XlplBtAlGtZAjQrAlr6cNCDwq83scu
F3+INLFMv7c8uozqCwqk4vaOOSeJoOPIG/vd08VZbEROvuZj0PCb1umfbOAg0CwMH6pBACOQ2K5V
+ThfRUTlJXDwS9Q1AGvHyB/GHmeoqENtO1EhlV8e7QGDTGo7s65ahiMFjJuRNdKndB5zSfakwWDz
eIUBtaGs8b7sZPeMpk92gigM7Sy+e4JvKs1rriVR+1I0IlhKizQzbZHHq3q0PE5j8I9IeptjVjui
lY2WxgZSjRDsq3y5iNxiD1YVm996T9VXjZhRVql0uzRq4Kqf5/4aqPMwIYz1fYx2M7GvqCf7uWsf
kuuVDvdh7BoqngUN1Tt1GRCdy6zQd9B4qMn7AQbYD1R5pSz6LC5RvC/kQQKYJGCuXc56QHj9gDGS
P3UrKfGyRLVC1VlKjUlcBtBlubpq+u9+77TVuuGhLKowbOM9SE6a6VDxEBYJfqQacMY2bJSMpWbg
XkIgA4Eia8NRT6EMpuippsqbwjIyWydhCOxsCJp1bOltp/dwExgiLVPeiq52dSsxdIkgXdjB1SYh
LAB9OwZP237ncyws2mslw9AVAVAS1Cb/MimCHLBUTPBEYygoTSytlHynabNRak2X4aOOTE1Lzy46
rD9tJnB65a9NkxIHGOFgz2TLaO7TISb6fSVsc8ZX08vx5FszhVlCaTLTUDzshVhmqTf5pVUpVbbT
thyqTt2HpxJEVy+FbzapsxpqajUCLrjFk2XakTO56WBwqLEM/88O3nNbZIm/ayrJZCcIpoLQznOz
VO/ArWP0Q3U+z8Ihr2eSm06qxyYAi+anjglap7dtploeCR18VzCwb4oEUHdhpbudIyoJxwFlPGBJ
FFKKCUVYNWk+plMdX+z6W1ZzENauesvk3pJtE2zMhxBRq4Pc5TMHoN4z33h7YRKZVGXqQ8XZ2NO+
Z3js0rf9WPOFkgkioBOrXQwiFYHfH58fsrNmJIrDkodJJ/A2/RNYYKom/6TxXzkGmYjsXU2iojtt
eSe6vE8RmatWeEMcv+aOoI5AzQ2AsKICsMuMPIlajwgBeX2oeFZuva7t3+Y8XTnfGF7pIJVtDwTS
uVSWNbvyXdSh42qFN5uZE3EgJGUzegrFya93YFa8zYIPFn31dNVSrK71L+dM5z2fn5ir79b1ZpYg
3ibr1L6PqzrskEtfA/owd11wcv8cXU8Pchzl50+YROsoT98imMz9p8OfL4oOXVRb/oKiHDM8S1AW
DJeOFLMGUrFqNLS2pvSqkjYtseN/uo4ycnRf6S/CvGIKKnAdKvQzyzzfdD9agUOk7ilh5MQu471m
I3tqak8BLAI1AUTBBf/A6ay0D0JkOAwIs0X2cLAvE3vll7fZXSN3/L5JDNdhYW2wPxFIdpcG2IhZ
8nehFJG7UXuzeMP1ckxsje4W97hObvFVT2YhFlucPjcYArRI/RmJaAJP9srj1fPs8N3VioUta5XE
X/h3HtrfEa2pxRUYtK8AVjkCo78U7v/yylTeIM+FhnjJpuWTJlUBAqLKO9QpfAWmDz40uq12fKZC
/5rqe2lQOStdm+QKOPOMeYcnpN5Eev/VYb40LixSmI9lsjiIaokctFW/7A6dvlpxK2x1Ssk/titZ
wkKwAmNBQ2BHL7UHJCXNKyK9ev21N8IxXnHR4h5CHiXLpumCvCPFXturVapEIDNCpDVSnt0CaVKF
LVPAlOU3JPDp2VxZT7ATffJovMBl1GxP38y5gykXj/bqIetorhP6vAtowJs+dCFq5bcD2+sg0nm8
UGyWzJDUe3PvSrwjb9dCfaQBbC/AobatG/kROdDGkkKbzlSpvzWf2fqO5vd4gaYc08W0h6jXhoNO
lWLi9mOariGEe9Hu7dzd/t6WCGXv0Vxnos8oJrMK6n+w5i6WyhNdfDg0uvspx1j2jY2FQSXimgyK
9fNOIBWHYxAEvc0AqatBuJu+rk8U4us/D0sgpIM/GbYiZQebtHfvgUQ/qDsCcQOO3CfrwbGHZ+OR
EAoATZbgj9qTlmwWKGWUbbG6v8TWMtXJrjB4+s9Ighdb3gNC1VY9C1gKt2RGoAGd8CH23vWw5lWm
CWt0Nf7HjUf++Xghdt+gdNl1umdbaCaf2IbhQ2YnQMjYXXcokQ8bxjNOB5bx70RqYI18PDbQd3zn
E3W7fi4/SHhnbKOzy87YMFkoEwJAonD6RJlsrP46jCT35+RxbGllB7r7ssVnQYz4ZsUmOqa/5hBd
DEAYJAUHHOItcOtSw5WNau2qvf/2QmUl1WeT446CMRwBinhI6BCeTC7IRT1hODajWiK6PK3yfpvW
cEgZhPngFQ0rvoMypnfHphf6JbCCg5x64oy7eD6jM0+1vMzN/ywIUmR3mwO69af72dgzPCCL8yCv
41ir/3qS9RVVGQDPnA73fEO7SdwL7SExJRpmkzxgcPejhe7m0K255Dknu6n8NMRainpcfR62Urki
Kya1hKjGWu+ETp3uoKz/RzRDPnvbduUtyL6O0geWT2HQ4u52cjb3LiBbUO8ybQNkxV0SWzrFI49P
6fz017p9EfxSHNpy+FGR/UkfP4ICUc/3g50KZ8fn0EjrwL/8f7ETjh1aGdvcVGJmd15gl/GxGOpU
mB+8xnQT1n0H1VQH/lQiJRH2Y9Jf8l9k17I0gB4fVzgnXiidytcRygzlYMK8+1ZwAAN/sZH8tkhs
b0x3iB6Pqb3Kg7zeqO/NJinYg5gSS9qxBUlij3oMHdsu7SAfnTK0/AuGMhYEPtxHoV2h960Dd+Xm
8vNh/3sxDRUaFVDNZbQbWEj383m4bcOn2cJVJc75IXrUMIBOwe0x7SK1WsvdF+aYtI+texqGndEv
ecgHoVoUH89vto2jaMqE/YVdMIsDb7XOVQiV1y1DsKFYzPQyL/CicLJi917pPkDL+fLFhrkMWbLG
4zAnSeRUHLEYV+XnM4+2Hz6UJz2bi0dVu8/bbbxt29ejeqY06Swzp69cT3qrItq7kdD8viSewCKQ
BWetSrlgGfhXO9oducOaoFQPX3jMFn5hcJ/Et1SJ30OP3G5qAnjswIb4ECixTIJy3F5Db19ZBIDB
3nJCtxlC9r+MO4Xco0Z8a89+ml1GkEG+nJXgoPvjGRkyrG4rtS0xef8yjknfSbdAlq/k8+S36Ve3
POTXzyrvp0tT97U0bepxLIbQ2m/Nhyz0Jc+9QIpO/mXLz9oyIPUQ6h3zXMQ6atfyH9To1MXt0jdL
jqH8TvKLi8r7fM98bYh6Ee2k+uReQSHhN4OTiDA2dL41R1io+LNmhqb/EDUkTYnoTBfla6qhpY49
iVdpcPxEB0FypGFr1H4oi13O7hyoPDDMW5rBb2b0x1Qni93LgwP4mHlCsuIkR9Vlvv9XtN0e4nxb
mUx2UtJUuzCWQRUGZH5BnevniEfiUNdYkoJ7Z+CjTt/KMEhZcxIHTvZP5G/hrM6dIDV//OtGNXrA
sX/dRnv84vYydUQitEwz1Opwor9jh85B1XMwKMSKZbyL913ZCVIegtOR38P7wYkeQBtiuF1lBYdK
Ph1K1Y2y0+2tM4AChnkft2ay4/2CfxP6ZRkUB79K2dzF4rSyWAXA2FICukfhXgTXarlUdzy9nLjd
RMywsV4az/uMrZ9HFUyzrQuwMIFKZxX2yTCzq2MnUAhAr5JCJ75hGiMLf7fLhaetcgzZJoaAx8ND
LITdbk7nzONVoC1c+UoXZb/YnRfG2G4R13h5NEwHNBHFLzLta69VW8JdZf2qDNFmx56ABpxjiFUu
W+Ia2z9PP5crrfaeBB8ku59L8c5KE7uwIdOGMmaX99oqd/i4PB0zSmquIJwdCBTjpHRuFa985bQ5
pZk8O4miEVDYUZ5VP5jl3R+F/THLF1KSRfVsqn+lKqHk5n1VfdZsf1WvqWcMx7Ke2qal3EZ2DL37
Cn/ihx91P1vdByv6VvH40xSrUyLvGSjUOYpuM6gC0jkH+l/nFI5gRIPYqwqSGkliuSEYxzDvzUBR
ipzWdcfIjfc77Uzbu4zfqJqIdmFaCgX2ToLxXCePVKmY8UUM9Tm3ISuLhsSZupHYeFzEYEQKY4Np
CCuyS9V/UESfHOsyOeTYvP1XRLew4EtNjWv6k0z3PhZelsqe/qsJTqefqSZMosMHFmWl5ArHx/18
U0dkl0/Vy08+oaNL1kKz2bjKxyrZ91N8xAQwRqVHQ24EfdbhVo2saTTjmZSHGe+skuDGsPbQ+MZN
uLwChJKblKK63i90wkgMLsm7N3YU5Iv9MblJlw57iP3FBXV/9ZkEuPi/aEW5Q+eImbolaJockc21
UyjBL2mVWDQBKXCZPBummcR1E0B8vM5ZqsZecZ3Kr78pP2TJFKjoOKYYulynjmyzSE6sVDsUZ6G6
wfeyVfKvoalpA5qRCfTn1DuvhfhnGMaLw6DKQKeKB95IvWpAGSuGFfVeDxfrwhg3Ev1clJZOsFdy
Q9gYN+U/KnvypG17aQ1vF3xGpg/dBMvF1xXgbIldlHhk66cUrG4HzANXR5WHqOikdFV6htklBeQf
PJ5gpzZKJKKtS8hKiWrWjjRgAVWlOgJuH7KGBPuIz/szmGgXIecvl8eBX9oE4bzp2K1QudOOay0q
wFbBCaGLKYa94eecuaEU+Qm6mlcf2ISFudx1cS7rqTaJSffdGKQjMcJx6Mcn2IvlBygj+emt2DKK
Gjll8f7kbkIjDEggOo+rjfd0KRJlaD4yq9KKjBo8VKuabqrAzOR/jPFJaUnPpEy53S1vjLCFZtlZ
bmrlAoEnBmX6fbiXjzVIqD0KYtLtCr+xxqUsLsFAxeiBGYEbfo2bv8DPyVWA2ZFDvrUeGviWG8NN
mor1lfgGkL1Di/CHD+lD8cB8Zu8ukpzqOtud+bYpgb3sjYjjRwcL5yZHiTy7rjznTqiKOcWv2upO
4jh5Dd62zSzUg7zzfKpmi+hHy33Lu7+/5iX5pz3cJKsTUgTLiATvA9b2jwtUMPyTuwt8TZv8ZYh2
LePvgs046Kt+omGUOCf9aWZ28oacGrUonHeW5KUMJKiCsBSgUMfCtbGqROunroybG3AWpmm4hUE9
llcIfiAjsdtcB/WiXPzlrw6c0CzliqD7My8woEk+T8XHWOfCKkxHRIEGaM+P/elyH/QV1zIDfPPH
XnWMMkKScq+hpg9zjUkDQxFnqXlbBAbkJdXbFVAtLcOifT5Qh+8RgFUCgfWSxTz/dxuudZLPHihA
wnPsebsbGAsRWEojxT8TeKrIvYgsiUB0QubaGKQxswKUX6/V3YwzIcGawthwbMU7qbRbkU6dkDGR
kw8yZS6TEkuTesF82US+KtspOntV3NyzUDnWv1Kk/mgjVYu26xwSmuPtM3ar4+802CEHatJREHwu
wC+wt5bGy+shoRmm6upU4PDpYu7k1kNbkjjouF5rT6RK76kOqcGW/aTHI5nov95ze7ErbOK9F1JM
aDkFFRSb8R/gjusl4wTfaKIsJByGtvy2gvCj2mMp1K6/fyta8bPRw+1US6Y/FJoh4UynZFNPBBbp
jZ8lIrRA9pV85hNTL37l+ETwyYt0/f/SDUn9xknIEqRgKdp9A2BMJJVw34xnguzbRKXWMU+s3iUJ
cxh9PyFhQGVxoevOX7x9KA1iBNHrJn/Y6HVMm8QnaozuiGg8Dz4J1DIpsMiZr89OCnM7NSWz6t0b
RmPkOEqiE+B133gr6VW6FAL9thCb1YlfCwPGXBaKOw2TfD03IaO6mE90OPQrrVuwDDMyFCRWqG1J
yeMZmDCpBWrO8D6ygF55G1Cc1ZHXj4fgn3/UrkNjSBeIIvNVOY53CL7zZCh4dXJknTbSkQ8a9BgD
qCngNjLngyVyvh5pHukCeoTGOEEGrBKIS1KOxD6P4iJK3xDwUM2cu9Av5EsUIyP9Reu5o8rNDfqE
K1GihGqbT6gx7emW2nsH/F/Ooh95NY45ClU/sb5Kj9p9hbNlZ0A/UCH3uUzNDc4l6xWnE8+ejw1Q
IWt948iZc1ZfhLC4ZY2aETivYqNm9hhkAtfUbSajPSwEkazO5JCIzffpc+BsnfWOtl02djoWpFbh
ozIeat+1TuyCIk7HJwcmedQiQLzhK9BrjoN4GthF9V7Pc8dccDbvwyfngQZh2bUUa+ZGZjajkDJf
LYnbdE2iKeXJwl//3rKpaoDDm3oDrwz/p9gMIsIAxnHFmRdedCF8irsl1zcySJQ3NLtBOzd29pGm
a1w8z60jzmw60VSlxITH6qH2N9+4OzXOLvrSY0lyxEQlLN3h7Ohu6HexmmlwVcMWykaKBwQnFQhS
bO0h+G/bKamJpKRMgu5O9L39hZRS3jixJBNjhoIqyHx456Q26c1eni1+Cm8/tf33wE98V6oD829C
3pqu63RY/Kn9ee5KG3BaXvuG1iJELrU4uSWipY6uf3/qWOx27LBecxQQT8God++voUNssRRIHS8Q
TktaZY6Vr+dCo5mNYJ2FIhJDvodkbXH9EnZvAu6ncKPyI9d052KLzBNe9tuwHmbon2Z5jg3QAArk
F60iCgmde8DF0Lxu6lJ8V0XSo8JXvVkGidZN89Ssx0aaVHRvwSZa9RLxeeAwl3wuRkTicf4qGC/k
ivMkBYCD7NXWNb2AzEZsiTcruBVFt6sO7wkkcfUmSTMmxHTTlnynJkF3QqH/cg06VmU2cIgTIuca
44jaGFi73I/+euaJZXcBbo/xQKcYpYDplhsAUqsLAPKnZMOSVeQnlDSjN5xyG6BzTKf48ogluGv0
0NzxCccrlKBD1ZzmLxVr9n1WDX9Pg6mLPS7wRZl1qaAeWyGz+lPGTUnp2JnlD7YYXy3OhcIeK6e4
Ke+IlfU9qhfbLuKCsmpVg9iUbENH6rcstbDfpaMCFBQteNj9+pynjATGoAqbJlPXwKOI7MfDgJTa
fZ8euDEdF8oNcLRVG0/XdRIBQ6O8BX+Kr/OvZ8kIHFocin9ttRd6Nf65t219DwFPHKm15YN+wO5a
c0PT30SZHSd4+/eQILgkZAEMRAtK3ARoEV2Cz/DBPBh69LnIqp+AKp/zhCZew1FGA/9lPle8M/HG
ORqhmQs6JA9UJNXQBg3gqo4aIW2PVz3Er+YcV+xeVJ89zEQfGjzOg7KzZziBeVLxFgv0xLcTwaK5
gI2ikEtacn0dqZ1bQX+9AZN4PkcKoDF2cfxC2Kex0p1zQ1CG2mTiKn5hrsEV+s1eM4qd42RKiivt
Rk2ctYdzbObb56qUOJfQbhYfpMIKHptRDyJUEPwxOH/K/nfHLpeXnv5uDJ9nKdmKLV7eDAiVf4xh
kHCLjBT9DLAEPfcmI7T+8492gVw44y4pqI1/CKNx3kycL2FloHAQct9kFNsTbWI4nS+MrmWNETHf
pKjM2W7q7hVN/K7CO5+Yab7LAK6bLqBJ7IqnXdg9izcDknUT5hvCi9G8QPJJ7ULdcZUaR85Y4R/D
ccC0cPQGM22dRL1ogVOrfbahNW4sTBZXm3wwHjbWC0g/HPBUS101/VIvnDzAiRHQQbQRyguk+Rj0
rpi7+ML62FLtRZOc6rDoSbGWn9NxcRGXXnN59MN5IuzkHp0qKRcn1sM4zPWNYAJAPb8vE6GBgDTy
lGG3boUK2J+3L3/28Ao1cutdVyJLdpq4tldi72W3JF2H7r3uLShBa7bK1gZI3N++/OtnxmvrcNsu
jkznhVS0nnPSy4k+9Rh/ExIlOWz4+0aW1+Hge59kBOikQqlKRIPzva2fupytosHzjQ88QH8P6rxZ
MNIG9DNsIoAxfyQCrlXdy3ZUQiABJEaQNpdglPqO7qdIINYb4crGoKCNRa+pINgi5jG6iChsabDQ
C0Bu4NCsjbHXht09DAyMTFLWNnSOnUr5mUGW39WjmY4rXlfq5vTJiH61693lsqqhT9qhTvM4OHfR
dGNxbON5leepi5yVxRPWY474RvlbcMyKwAlX6sq/gvMKWDhVKI6ULbcAtACRPTPzAB9B80N67VRA
rK7i5Gq7vRX2QT8+hAXih/KkoAVUuLRBTWVPkOijb+qcuNLGlhOgdTp+LQGw8QJzKIKQ6yk9m3Yx
WIfpQZzPo4pb8UA/zd9uYEy2dp09LK525CFBzpBEsFOdaJX0Gc2QVw3rj6S4viyUiF8lzxGWXO7J
LMIF/Ts7sEyJdQkZB+4yJmZkZS905hg+N/7QHQcQnOVO9GPWMxxofKhKN/maXI4H9tRuTQln4r4q
CfwKIEs65e5toksaOaGxla91py/pccTsFjSbHiRAkml/8g29hWziT165Sv9m1BtBl7sb0taizk2X
kIGW5UG2OjuSENOUi4B6moUzPFmbcXxFml+zWe2Upha26slIBFX9LMvc0+N3PGUYDFAnKSA+nhYT
q2QSb76vaiigImg6p6gMi3dtNWwEguUdn+uKSz2eMAvNjLqoJSZXumhctqLzaJwwZ2l8g/wQSONg
DCir9BD/PCDcm3Q+FPTuM2UxwmAL+fJ0cI4iX6uYtKzD1IJJSlPQ0GLPaOp4laAGQzHFZvjEtPvK
Uyeu2XulCVNUZFRaKBCuuSknlrtaXwqBQlVswIb3P5XQmuNp10S7/BruPmoU7CaUIhfNsJYHyQqp
XOlpZO3kZ+ktyx77zrigoywPGRDYFCUM9qX469rHn1pvOSA3KvZ26w87Zkf1jAOGHLc/l+tahewQ
Fr+/LyJ+iAe+h5yEPeEj3sc/n88GYe0hpGL0coPrkCbh8QTIg3vAXwStKqwilsvU190CP2Zq8O5v
gWlLUUQfK+U9REkWOkwE1hfJ4FJUu8S4KpPUG9bima9iProdnFHVCzDjWBu5nTKGkf3f9Pp2D00M
0sGaiF/qDgKLcLwEHZaVuGiXor94yvUlM0jwlUiIL6WYNyPA/NI70LNSeNp8U/COB005I8zHae0O
xAFhrlv85I2apUXqO1uHWjkuAyZcYVCPb5XAFtVCqHesK9GgS0ynJa7IKuqNVUXkt5c+eFr0P0rg
j1Ovdvyy788mAxmAiZ6tozVDbt7NGhVessyPOYu02mLVvKRN/h3eEDbkP8vohK81Yj6MrFwRgajj
2vtRqu6cxpBNbmHAGX6aBxbkbWravGbBCfyZsRw+l4bcGJHs+bVPRxd6cDju98fBSuXpCr3O7yN7
DftxfxakysHvSIucTJXQ+nsRFga/PS2pz0eWeDPsZt1MBSK7gIjIHIN7FAuvcbFbhGe3zAcT5Uki
X0QSQOlXyzga8C3F2Aw0u3p3e/N/mD2VrjqNNn5of4nUr3F0BxPR273iE3FbBq4WZje3KqpkAccE
wEwiqBpQwCgztvhToCtUB5f829Ges1kRVQrlBuqqHFPIFBQrhpCR8tU8Y+Fi3zrnO96KMhKoGsxy
vmcfouhgi8P2VWyt4PIXtjPccnzHOp4oWWpALk2hjXJHk5JOO64jD4jos7Dd9trdGCaPpgyMPgm4
rFCaXc64rx3/8GmjrTfcWyG5k+l0T1xkJb7LjAIv6/tQUU5JBJGdwuiHi1lYpPmMVCWbrqnPfiX4
i9d38L2uvQa2Ohc+XdIGmdwGDo9BjuEMLFXY60UQT4vbOX6oecFjSFs6QBELe1d1AmL+BdTy9InT
OhEJ3odvPwPmMXpDyZ9CgKMUV41wkh37Ak77tbm6hGZtw86o2K8qiTlf6VZtyaPNKEKZ9m5PAU34
WwHUt46IFaGOgaemuY2o3Vl7JAKKfsj5D2dTpbFdPcklBlFP0CHhfs/vsTBSQ3QLRO18Nbubxo9s
VYhXGwXvLGFU4remxzFr03GNJ4T58rtVRSbnda1dy34mnbWK3Z4Y2CPTxwAnWGnyeNLGlGOX8WUh
ZRBeIrjQQTIvf67XD/CHaE4HXQ0x/RVLeyi6xO7SNVaikdagYRo97mIGzVqFizO+/t/BLbN/JdZt
sm0HIGPeUfO5mhlyFi1jMoH9lbL+9i0iMwODhAAC+47OhhI9pVbDgaeQFgnYAttvSPX0Z24QGUeh
lRNhPoBZBPEEUBsBqlMZHkNGgjAbi61P4Sq2ty1HdSXF1vUY2J99N1D3UII5g9Xiqf/loW/YUDtr
iNaQaT/qfnaQBPrd0w/jzBQGiPoNB/MSk0B65ZQNklebpXdt31WnqrjfTz6P5i/pz6UImgn/a/Un
/ZkVLsuXN3EUXonuf84TqPtUXgYKJ3AfNc76KXpGZyHmqUUY27uGTGPa/1OPNrsAkKg2nTWApZBP
pOXGfd4SliscAStrtFwcfp/E1JzLGyQymisui5rVcKp/meHwnhG1l72VqVDYt4V9+FX/cIKF9Hxm
WnoWRPK2q+O1dvp8eV+pf/fgQrvvV5hotcFAuFOIgcoolg8SzWin6g0lOyLagO9dqG/ylQevqAj/
sttYAuv8u1BkgbeAM0CMED03TQ38B+z6nDI6Yq/x9sQGCqb7W5Bx5ZypmnIzFWxMtjGVApsHFtUQ
M0eCkQSk7Vw1FSfmR5dc+rC92ra2KVRcb3f9BfNoM4pUd6eGyevod2po9HXHLhvgOsVHYlkNtBGj
5bDyOzYrGOTpMkXnSfcXP3U+aJG6itQ3t5WwpxpDRgEFj+xFt3BFKwQkNgkhRale+mCKwKc2Mfkb
iyvbza1CvZqIElFGdKPO3/8C8Qy68v3Z21cwom4zprJshpkLDU3fWTNsbqaMzEo5j+H+M0TNS3Bk
whSMpXcll0RGN3+qXsfeiKySz116Fc1bYWtWGUp6pQ+Ee0/nmr6ilzLv+l3BTpMB/76QbHqA04wJ
mRfRQbs0wzDy+jNISna/vKJLL0Lyr0ZSGXpaYj/5+nmSoJSXQB//6aHCItcgP+b4vQV9hnQW83lR
YY7AXafh3etMgdeeN8XvMRKabjVtQvnJgx9H1lGhraUub1xGWw7pyxFa9jUs+hoqGS1Up2jjy1IW
2DMDTHI1xVCLySRE25KV9WCU0sufBp6jQIntjOqBLf/xbxzfq8zEkbjvJqbK8nk68Rh67ya/7RFv
T5pamTWUoQ1NkchddEJlPeVjfmIEaE1Ht915AsXY9snGuwI5/GMLlDTRfbKx0v/ZNclA7abOAkK7
2SBl0sdl6Ay6/ksR+ki4HJDaL3FGCJG0o21y32syMV7GMCd0vQ7UlrvN4HUBztAivGenLKv5AUFJ
oH1Zx7eF4VC33MPyq17FqHiK52YjaMJz6qnteGnR9YS0GfTSlh07GIUpBVF7Ruxua6pbxyX/2q5c
WFR1JPZWCiMegMC+G3+1jO8d47Z9GXpupZ49yhLqwaXzld038NtVaBc7oVbTvG6ReEUuWGS9MzSU
HQh3KriyWcMAV/iJZs9noHSDJ3uv/rTN+VkrhLzXxuE+8jjf/w+6vcRUCU3zGi4ON470FTgtvMPL
Mj9tRVYL9/nKQ0zMR+5x9AYj2Z7kx/lHmtohl+Y5qTT8GtvqkHRW5eUW9LtmkGdF0Hi8s5V1JSJm
Z0gC+ZEaeaAWiHIaqx6gvWAEaCuJ8Vl8ys1goteP1batk99fqlemxegkp1PZVluJBc7XHuMVVSyn
wqUyUG0+pkYnYdH+3+pQerDhExGQiItQAJ8MHr9lCCuLLh4WacKEJBtp11z4Jnw1ywcTlaKnI3Wy
nnTkv0wdLyJdiiDEGL+CmiU/TBFbWayUdSQUeiWvqaabEfHoML9U/JoaQsk2lbQPXNhbaVI01SGr
QDhSS8uRsG/eNP+a0tTPgFFK4JEIcsq4fvA8SNfIQfUOCFm+kzzOR+2bLbl2RjiWNQun3P3naX7M
t9uJqdSRsEMvkYmX+7H1iJVt9lGfWzjXus+XHBTfZREs92xaD/OY7/GfYu1oMnshfSG3zT4mH7D1
CuEO2x3gbPENXDe098zF/5vGiIuRHdpFHwC7x4y17LWeOlHaWDpKZ8US1Dtfec6E7oi5wV7WZSYm
8C2gL5Np7esbcLifCAG+EP4ezQeX1PY+k16J2F3nemMfPPx9wGx4REFtrd74m5lqu0JcBSxgFYsw
aIJBKFkkWGYJXYrMuJXiNpmDbGDfBMAqjq5B0T8otHCTuyz3vnnAFsSOHopUwGu7efgrfHN1YwGQ
t0W+0LVbS80uzzgUOe/lEzzpUtdVYek0wZEorStC6MTgCuDyHuuMYCOc1LN2JsM/Yi4U+cc8sMex
8Q05H5uPMEP7P1RY6Xf532y5cpo9AaTKzW/dEA+aeA/V9qlVrZkOoBgqAK40XTMeRb5HGGTvxv+7
Khd0qGs/m7SLxMaDjNFd1uxfEnfF/jKMpMLeCeTsbzmAguDRfEgEJEmJSRLj3KbK6kFu3c9fHIED
CTdzB6UdTNwazJFKPKH+uChjpzs+mI6xuEZHMvjiXrQ3aLnTeDXqBO8hKTK4QT3q7yutlGxdyE/Z
ubHBx+ZOmMyyocVkgBE9UplO5Sd8lLzcqrBItRbgH/qMru7R7wk3pce2j+fXx9LxgBopwM2zQnvT
OL5WNc8vqcne26YyMi/Y/36oZvTCFeIa9/R6/9cPoRrKnNt59nuW34TgO/ata8bcbheV1AH7wYO0
GzY63bzYWCvAzNJOgMi+trRdHW7DG+5PpzXLDpLmhJHhyqxVCUElawhI8YjfasSnxLrLHIeNiHzM
43aQrfMi8edttUCUV+5Vy0q5sPGPCIEA+qskV8udZ2CPqT8JCJjQmVy7KNKH4V3BC6yJv7hgIDgd
N3yoV8YOMSOJXJla0lpTTrh2O7fg1G9hxfdmqn8Ij5Qy32/4SFu57P1mgNx01sy2Wks5uLekWMAc
p3ioHFZLEpLGoqYMcYSlcJciP4H/Uk5p+0tSe0jrIncfcd1mDRrFn0KqTWnrIrRo3oOZdQzRjM/2
0edP3Iawy+x9NDbl+D4/qzFjcm1koCQ5FsErw+ME3fBJwSrBBrJ6EUOf4IyResYGF0LDzqbOcZaV
56RS+YuKJCGAlgZT7OTpS9V4KU8jMpa8w+jzOQBlG18M4CNy8jQcBrZDhqoINfvgEmAR7i3xEkeQ
11nBSocPSLweELf+Sf6h4LTTfcOHgNWnYg1FTG3h0cjtVDGMNB+IqkSzJ4hJp4u28QXqJn4QSYBx
UXsBzP5td6+GDNcqUbKz/yYrHARQ7On35DIEoaSQUO4TkYemg3vrhGKZwPJ75HDVnSM8pXuFb8HM
0PGA3it0gRKj3KRpnBphEa081yewl6iZaLLiFIy/n+vunUo6i4/pW1MWuxdzyjSXSPar+gNQ6XbO
t2uRUofV/+VYOksKgKfoXIIkAZUbs5yuUJE4liCrbJV74Kc0pRf/JOh+YkvJOoepb5CXCPuVJEgR
T/KfOP+UHo3GGPTGayklwSggose6YVP7ysGqIOo+JV6Fg9Y1vpgVcLpOm4ab+r50OaGX67cNsxVJ
SPHizcHwCSEURdehzZgaVgeNfSmIHOXJu+pzFXGkPq0fgN6+7+j7TDLRr+02mGkuAoOLDyAEqj2P
vB3tu9hMqzX8C9CVG4VxHwLiNrudGGUZaQ6DIYB0GFrgAi8ryy/HpTKQtu+5eYdUdE6M8NkurRQi
6UPdDxTI2+IhIacwnesQMwhr4znaqLtL91TLlOAMMHkZN1l5Kws9lq+l4hduG8Nw673YOUpJXuKE
+tLJB7v/wpYQjMKTRz77q0/u2Ho7aXXclJB0FfeJqqCUlzVg7nr52MQs9tTddTXQBvapKZK+gx3Y
JtVIgRUVuy2xMpFU8g61nBA/RsZuf2UW6KG1oYZRYjSjfCDqEHFoqYx+XG4vCAY3cFZd8ClV3hNo
8BcZw7gaSHGTcb3AVFaoGJnNDsBVCN6C0kKI5Axpk9xGvXYgvs/KO7sal+gOlrVMEe4meogrG9To
sCGPXs3L7SAQ7jZy4KFyi645RGKT9o7GG2Pjc6wid+iSOp2mRXElb5KKej9Hn16nCYuHVmSOV7hN
mSO7n86BEBqGC1rSrlx+x4mADIXtwEwNXriRzjsZVfOsxMnTiwZbKHtbYt/Z5D/AfZn87vFuXUyO
nOzdLD6FC/34HrdeHAMG8mKw4gTJDyI8GkSU3RPpczxJrzlkirAMS3rtwHoT+rdH3+AccX44UYPV
H4zwMfTg9iDekPxRNCLXWH53b2bwSbEkSdtmDwEXQ98s8fJA4hw5VLafrG8+CoK4G+kpSL99uc10
R3iW6MWAZUvZa94aixcRwfDiprqad6wcUFjznJXgsrrusZX0koPuMiuEBmw7s7p0mOmGcL4IjCH9
3VfnH8o9v5Ixvb/rcVRBEKh5RpI49tBIL7UQryws8ol6G3cVgPSo1LnvOmt0BKXxIKM5K8S6BWTC
lXgLJPR3NhHA0ai/jln262p2yAuZ/Hy5sZs4Nzg997RT/3b1snGO5zzAXft38TMFjd6gx4fB5FSq
XPipI6T/RV8P/jQWsFi2YCPRDf3a59QXvJFmsIozqXsyPcXwK5ZINvWvSay/27vYm4yXYdiiON/Y
0WrCl89xJnH/aCW+EU+Va3qB3p0g8SpFi8xKCnzUNTPWXLiL7MEE2rqynfszZ/RV36bLZYOnS2Se
gcvxuZRB1LAaYNAOa5+cR48srbvyQ9LJqRY2OSVWCvqHhLKoVX3HeITpif2tjj7ImyMKM01+skOE
/TNQ6HbUqdpcmqPzSavcECzRsz7TRnDEeNbIsCb0bRQvLCxJbq42nrvtAGeQ8y5SC8WExP0ekdM0
kMY2SyvxjNkXtKeXpdqr+fHUpA5hPIrwqhWJnENQ7aUfC3ml1LAIHjGhwwzM1h3e/nJwA6XMv5pa
q6s6iOJVbSs7cDJoXayBRpRRe+HZ+p4rC9QENmjuJnAr+VMWhA9ZksM5D0ch1X8rXur+CoU8POUB
O3s0W1G5dIOOgwrE9hY1RucQAfXYv6Uv6tLk3NdKPwMCtVJYvIEpjqWtusGz+GmL4z4hDAPHyNOs
Mt/mLo/WHV0rMh+0QQ7NKvyv9Dvz22lKS4fxMS/oS0eEUSqutYkL7w/0qTaP05eIt6TGcT3CXF3O
H690laSL7nSUjgjEBRWhisXbCUlF8TS08L67EoNC9d0jw+ArLpopzdix6jRGUUH6vQifTaibsrHa
c+hCJTrdG5cmU0/ny1QOKbBL14Rw5di31T/H7gzPYQluAdXoO0x/lGAjbhxCr61mLOSu7hkr1+J3
rwBqy3Alqakf3c/Cu5DkT6OBDyiuFhZgjVqFAqJWZwypAHIsBX4G/pLDwJPolX00mLUw+9be61eS
izDv0WTcf8bXCmk0I9vtJlbbSpe6VQ4UTQe4EzD5j7GWPiGpCDrsUTe1OKXVrkw32clQxYNmtKgz
brA8KwHZCiOop3CgN+ffRxX+SSBDq0FjcTzTUFxtrywjx/hnUoOreikdsfBRT1B9yz0N4G9LRmb3
sCUqJGdPYgT4b6vhQHH73fE6H3YvupsXcHNRXoTmaN0tXMvO6A035QdxGRb+9V6nfOl3YtcM4MOP
uIOm+lB0t4FJSFs2sY1vziYRmr0Zc7fWGCO29EYxV0o4V2J++TeD+Bv40lVn2lZl8g7WePOj/DSz
2Td7ct8iIZNseDw3NIwum2sUHHLvWiWYmirShsZLkC++zljgICWmeZPUckO6UF+V574ZIuoDgs8m
+FOl9NXhwrB0ocb5qZo0g+bZqw+3mNSWEilgO0Eg7xQUSrtREzoF4J+ljGpypZJVJayr/C6c+sIp
lFyqWQzWsTufT0w3FRx7VbEf9lbjUG1mIA+0BcUsx5zKaPhP3ey3g9pijweZtF+FXxY8b0bSkEgk
2R+h3xgu7ZroTivXwMGtpsimzyX/IwiOa1cibLbhGYfOZt9sSTHIHYRy10YJ1XriLlyoASey0qF0
kMZM8gpTY5GmwpYTOIMMi6ZjnI0WPQNwc0qO2dJmtwGu8UYgQKFFgeCxpg6ar4SlMlB9VKvZlCy9
po14LC00Rms4CekOaSYePpUDVMnblwuDqBiLW5opMhknqDToN+k7sjwCpLkzPLde1eNCoX6eQ/3u
84gWZsqpMxogX99NSb/sQPf5jHhCuHbeFO0BrZXvLajoMyMWwR7fvoqbeNclDLV8/L9jXkrRqXlK
4rGvDhZnwQtCsMaHFm5H8X+4GKJWBKSVRcexqwDd+cJ0vT5OJFP1OL70IXglSLCdbZteJ7FAP8Lg
kN+JCw+VP47UC1151BAHsDmoNgXLw6qmRASzr51um84X8trcNcdSovhjj79b9PS3qfI3iS/nhsql
A3nZ/sQ0siTWwCxb3sDW0zvOZWK43UdVXUnyALueeVKWsi2ni9nhtIIjbwhm4RG4b4u0hcDjUyRg
fIzqQDo96dRkJ5kJ5Ipq2Hi02xHcFRbut9cOCPO2EXYgBIxcddmsjf8UzsuJyr14h7ulvjFQZDCG
l+9YSNMbaTdSYejMPRcl19LRFiD3LHBJ66bequyWCD9FYrTutQjRIn+BgZU/wvrsZpYTeh5Nnsaj
OzUFrDxWWfjZUqiVGWmCDgMffrmI+tLJM+V85OGXS/kV/RBogX513B9dwFIelprlgMILcYGHZ9rd
+v2+g3e3lvbWc+cu77PMnGvjun/5AWvGVoURBKtqvAp4kFhSgMI/fzF4O880M/F45PDmHxI1fY+X
zrWMBlgDLg4yPzI/AlvSz/IQNly6szgWeEdbvoxwaucRxiVf6D90tA8mLsJ2oCLFZdqvdPDlRvIZ
YlAtvUIyGC2UX8tCwlh8/Ya34+TN+alTE0CSkAocByzNsqiOt5yhTG/hETXUG4ahH8G/aZGUcxS5
/+E8Qylzs1tgqkFBmQOHJCASVWaCTgtGXGcsQ6fy+NKmxg8qwDCiQEAG+Ljlo4hCx+MXEpqCaQzl
1Wnj+XRCfsWD7Lkg0aCfYcCtaXjR+1N8Uqtn0iEzJ4MRPZKnC9PZNlpmijScU6VyaA+ZLE85Q+Zm
Wh32OuBtSJqh34QQpeHgt+LhKUiu98BLnhnhEnJigxRtgruaUkeAwLBNFt5PCtbEoNWXy61bCQxO
Rk8gYnaJIJ5JPjeF88yGs57Nh/2wLOI31Crzrz1X5ELWJTPux7ZLnDHgR12aIu1l3kY6LBDBkQ6z
9/t5ZMQ5vX1DAhnR/magHk2GqTdV7F/zohX5Yr1YuxVeqzNZ0J67PvvICLr5iv3n2QZoNUjWG0KK
ae7szcboJ3Txa6hYtKPVHsgQ1GnoPmYUm5ByXiTTB+h2Pmk9086cK2AxBcJHbYqjazjZHpIarEEw
uCJG7RsdvXhj5cYTsLxycMlFVa46a4G+LP2d0ohOkx0Ziw73E7DAe0P3HOqdIo3wpcakcPZBJvwZ
pofOlroGJa+A5bPAp8zyAJ5VDfNNGrs5rOuFt0OKYNpsKzR09MVEOAeM+VvUQGDYubZlEqW4Nkmm
j+jlVj3rwILw/VDJ2Jt2BeVU0QsahQqWrNqG7SQ3J24uQI9FA8NQqB8BprbmOToJRqRJ+gsBWtcA
PtbJyr3tsU7K3fDF1eJN6iqGDhw3zsVj/EwQlFJEVgCse2x6Ne+RTBot5O24Sh8LxDZVvthr3ols
+S4eewRikVK8xlncEIi0PdiG0ZqPi6piNJ8HCm/FrJckI2b0oJIVDrldKLY1MsENWahIMNhI+4Pw
meOZ32Zpi5Rw/K4zk/5efqvK5S9uQMSf8AQkdZGkee1txlu8kfeXPu4D5tB0bNRW37RCuQdXsnEy
xCQi6DB6JUoxM1CLoFyZJcyeSQgVSH8a3JWLePKIHqiqCNkAElKPgJuvPRp5lhaMgA5++WaAhhR9
bopY7jdJVCYDqwSnQb6+mZcPdOSGfSo8dPLMTO0GbcuCbmFFKlw/8y2r+8UMTavdY5+bV8tClNv9
SOPx+E6BScfwjG9L7alNBtO7b3t0nPV9b9bD0DZaPM3BSw571D5wEJohMz+R4qRXjPUc7ZXDNXTb
4Sz36mC5AAOgqruY/Sxd8i/yNYphXxNZkndOjC3El4BiAjchWrFl9mHaBvUSXlgqDeeZ2B/Jwcka
7lbvjzILh5FtDwBshDUr9tf7Afk3d0xvRgGgEHlMAMPyXbulGDCcxaTjD9HGhnjJr41Tx5mQQvJ4
4zXEqqoBcdbM8cLz3SwMzXbXV81p0/vbYWZ/BwxyZb3neVNLydOFX/A+93NBYzDX8mo4yF+8cDHK
K1La+E1bFVfZ11/Lu6TIlMyc6+grLPbBKiC+TVM98uXPiG7fj86E2rGkgPPTOsOOjqPBZrpIH9M/
xsvhs+Tn+FKbBcUa+4a5g2OJCCXwoJqBWwlnxt9sYZEfVYitIV+eltNrdaV2d9HUj9crJn/IijPc
kXazTEK0lXajIe24FNUxUEIFsWoFTFxzAwpn6quaSVBibDuz8N+jfrARsENYGFWbWGrjV2HAD55j
a5oagjh/2LA+ZJ15i1rRKOd0b5noUwVmjSWw9cM4Sq32Q8KKSOOjuHnuQVNr67VrwEFBq36SqiMH
Nl32K33v36sR+p3Oui7N8aoy4+1/8Uzz/FqdqEPJlRwWGaGUfCn2UPdpI24EzBpc3D35CCbjPOwT
WiuPm42U+ktVPpBMS1N5c4JRnnZgabctPGw0qmD5R8AupFmWt6GEobCjqyqowMuwgxye7m65H3h5
Zh31pO5ZSd5GAeQ3pEiggPciddvDRjk0KckhcjZmRQa4e0E8Z6CYZPSwOAPvUMwMPIRKcK85p40q
ekTGAmd6OjfssR+2+HG/aO+oPhMM71XqWkPnrmv2du1uE0bq3HXar4BBJwxWdp/UMLLQJWGMr5fC
mLF8Zsbu9nAkwNNN4O2a69sFAxfjd7SuQrB48rU2jJHBdPG+aVoDBlkyTJBJDdITYg27utZ0OlE6
kM2CBPFPrhVtjVlo8gqUQAp1+UN6TPgJ+EePGYNytfkT51/u09C7+6XtsSZtEMdFTOjzEOi4Z4NS
p82eeswZkxSXujopwFK77l168TQoiA4Cgb4CCnc/jcvOQ6YLirKJh9oSpraKGa1d9Ya/hpaPlHUz
oqxAtFobyPLtsNDFIS047mSCQUFyvqOsGxPcFZyQTKiufX7XtCBJBlrumRqGYAWcK+6DvMHUV+Qd
f8Zwce2JvfhqoMLz3HKcwwXL1CayJkigWje5d3hiIElS7Lxfdvq6lFloFxJOVhvJvzX7dTq2WkJT
KtaitEPslc0tbUShacXJPFl61munJWkbdyBV9eKU5J6tiBKtRyFnIT1yTFaj4YYqLILaFXxKNdAJ
IJafOGVTATCm1unkPeAai0HgK6Y7151LJplteJmQ+PHPrsITJNO+W4kvny3PQemWx8syTrE7FCNL
NxZj94EnRPD2fPIo2o3OiqGusVd2+mzU2X3/DlldMmYUmU+vADCit6bQW3q86Vw4TTVba7WfsaTA
fMdD+KTgl7ihlEfkUVSt8P96CeDL8ZGXZUYDN1Q2TqraaV+eximGa4bcBcRAUpQu1bA6fYlBgXP1
10XaPeNcgy4xgo/YmDSLBVO1KJ4KG4rp3oc+kxD67qYKANOQuntNFta6HOIpXqwuS2GWG49hUdg5
fthxyHtkyJLcDW5Ghi7LTen+MAQYyvzOJlv1FJ+iXjxqkmbkZSYh54gvEfX4+20iIOWbEq8tEZvl
sYzvGW68cSte1ZMBvMU/SOe/2wIicd0Dd8eqrNAJ08aV2mYb45yHtHIYmGwA/3sux4YhzBSmIjZO
pCYOkcF17pnYKgKgIRMXL+VeOJSQE19EfilCf2vvdW4uEdkg1PUNkUCqxut6d5/9XbqdDTrzvWRZ
aCjwWdb3llJzS99NUVMpTjprxERstv9L8+xQHyL0UvX48pAq0Ix1PURRWrqzi3clhcW2zNufx+/G
qEMFqHvuaXDF8YXWa1/L3gegbIuS5yd/N2G+gvDnZTgKDKOlzO5AW+phdytobsvDzAJ82sNoTVbu
mlFUqVylAykiiVB0j1YRYIyUcQm8Sc2P3euncuRjne5eVrZ9nvyD9UNFg8ImliOgT8F+bYxceKjW
jgoSYb/AS0iP6tiHd2jxIvqa4+CmeW7TK3MMDRiK8tTwQMkSn9l7Y8w9wnZ6UmR7OyfbQzOr1NVk
em1FGOqLOTOCKvP1UgaNO1J4pKRPwS5h1wZX7pakuKl6ePNLkqqmwY6VUo9Semr8tGaR5TDKeMFx
EatI6hF+1Y9I2/JZUSMVbq8b/EhpUqJeqNYbHlAcxbG6yQnkQFwDvdCUXBiNCecOvfOSfD3PqhMA
AXDrCQ5IQv7XG/OKR7GEX+Uvuz9fxhAK9SofgSp2G6JvLQUODIagQNnTV841GA4wAudkjns0u/SU
uag+N3hj6dkSs592iElETG4deVrgt03naqvhnP9hYfZ0vwEd2ZJHeixlHqahf4GvRHaCNWFlatiQ
oT0FoJimIN5R7hZrKdMQS4AiHFWgUL4pTG8+IpuyCAxosfGol1Fpq/rbrIhQPG+Io0l+g6LQi084
68uJM+vY6xxkN5XpJnDtf1gPsNkV4wx8EzCRAG8mlcoQqidao25Ftw11gScCBECYPVd+8CC/hsJz
b/mvSjNiipRdN17pPHcMLFycsOw3f1WaSM6Gs1wvRmzxxJuYarW/6aLw48m7oyKTUDsJUZPSdZTt
Vw4ievQB+Rarr89QfnoW8tRdAlSPTqBnODtYZfF2SkaLJTsj4B60ySTzWjzRuP+OwFKMMJn1MUID
3a1p8O/2WYIihu5qHuxM6HJq64ytXV90IlCZkZEffB3SqV667sYojzVuWetz8avBPmolISPpfqHd
5JllFA+BX1/dkXb0RgRpRv4wtOr8uwihjiTCfncEBxFRkmwzDvJX1ISR+vsKTjDubcyfOy5VKGes
k/zpREq3G+TAWznIgH7TRD+wVXwi2RHUrjoi7Vi5hSZor7FYIW6HN0ZeiYCtmQtzPr8gGrOikTis
IBw9kYH5yjWcHuZ+isR2AE2zXZbovXO2jf/6CJmi7J349hgHQA6M+Ofum4ex5muXvqCljUAt8opP
9/aI2Ha8lOt+9s8wID/aSVRZ8puKaa12SSgIF+0hnTYWQycMOoBJOEKog1nDTBA+whjQuvU5nObQ
ZVVuWh710R8RiiTc9b0P6WBJkQInBao4pQ2ji27Ygp3Ey5Hdg8NUWpNuT+warBnAwkg9J8DwoSzS
cuqNMrqiG4v5j4Nm4vk7LnYGAwe3rrR6p4u9HlYIxpDWmpnbb0Hg76cmz/IhOUVVsHes0rztxyDl
Qm1yYdczRhO0G87Uq+W2ReQCgx1C3ZJleCXWiE+VQa3qZC0phgvL65w9j0SkjZqJBSiS+fES4WY1
tTgv702Ob72jDCGRKFE6JTSROVxu5NxlyHrpHJ/6loijtADznKpAlUJtAbXoBcb50gTHQVN1+Td0
bUNAO5nYfC2BzSg5RjfoyyOeIwy4L1JpZu3WBnm2LoyeU1VmGd2kZvATAbSzTygjQmQ/ktlyGlB2
vLKA8YPRw9eQ5ibKLKwTLbbS5omm5e+llVEhbxe9N8CCkC1ZKJcaPtceWb182pvHwZeAhaYiDFPF
qcEoPWQy/XY9Oxo4tmTAhkVtxKOFty2ruwpeDp1mfyNqDQSNFo7UZRx4ilxZO2mXzTtgmbVai7+M
Av9gbdyP4iFQ5I6XlcQfGfzzaE8kxH/zMASKS89vgYftbBxga9jWo1Y+DJ0YSjleIvSHq38nXiOP
Mv8dZBmdYMGN2zXlf65Iq36ZmOeBUzKeG64MDSeKoYJtnL2zQES5doVhvb4OybRQbDFRTtfoJ+8U
bEpp7oKUmR+fPHtJGniItXHmF/9WVjrJjboJiMJG/pR02ovgVK4KFbz+woTmqPyDhcHBtI0r5R5o
O5hIPrzNmKDUFyV1uqD/P/kze9C/dfNNDOdZmZXSb0bucjbSUo1qrDBPFl27PDed+6GCi02vipAm
NgS1rp9wgIAN/dlOauBkBwb1Co0zOD7Ff7AKBUI2Abjp17KdOEUUKBxc+HgiCxRLM6beIZLr4Pzs
6NL+yJx/Vqu7DDhenppbz9E2muHFJeTBJ0ftv/9rpJN9sN+VR5xQUybrONgczHXpiHKOJbtp+MHq
hhwuD2fGbE9bL9W1rZMvgz5MpalgJ3+INpnmsssRx24ZeIjRw8U8QZgC8I37xSxGUAXHmG7ah+1A
ozJ//JIjkPrtPzPmfI7XLM6JWSBFrJMwYvo1wkqhOByKbcgo0rmtWcSZ067bdVPdeNVf1QfhOHmy
ysT2Z50gvGmVijZoSvu/OvY/HXdvKhgrD77IjuOzLc9y1rgLf4FPpCZA9IuY8gvzIubMrwO3FDaE
+WIFwEzFkmiR0CyZaQp7xmeTCL9HjRgBCFLW4WU6DUS5XoSiHZHyY5bjhbwDidA+ZrYYOawJ0ues
9l2Cz2SttBFfMMQq0egx/gSr43IPP2LTv+MoLSo11pnJHV/KOCE2bI6EIEMFEOFuisDlAIvypfdS
NeU7BuaYltzCnTQ12TSHyBd5mOa8AyLBxUnZTiaxaiIXxmsAFU92yH9qTFGRh8SnZOJkX8TGWIAT
N3pxo3sqqcO5KiTyXAyGt4Ij9KNYh74RcagHgDvdn0aVndDLV89Lt3lnYUaoim5wgwKTP2gZV4BN
BTf7/2CZcwY19afBhvZHwZxuibPF3+JoGfbElmaDtz6f6Z4V+Z0S5naSqyqbZR0X5NqWDMaH4RJh
tyejM2TpK//j43wXNLQi5LXO9bnkA/unTdUy9LctXf1wLHJnBHnV4Qt9hQkJdvP4eMECLOmgvt6n
iLHx9jEUyUaBvReFFzwgmvqA9jZxpFctahtdZBpE5vOxoK71FdSVqXufz4nG5n78D0fcKP8E/Pcu
IvU6ZCVH7qWUnWU6b0j9WsIqnf3veytxW0sfxG7vraYATijpfMJgp8kcbnnzSh3Iza5hkT+75NNF
WZW4E5e6xwISkQYTzd9GvaRms1KuAoET5QhloPPKyajCMJcFhMiwQTnkIKFRxqVRq+UFcbTByZas
e6OOH2A8GbdozlJ2k6xTbj4EBHhrOLG/huAX5F90gTinX5ohXIoonJTE4KY9JXzVESophq8+xloT
2cZ5PLfQPGKGbo7OUg3j4SOd5xYMpHlFqB9xCa6XPonFMyaFk/65uSLmfdG3icjzQDspvO15Ip+o
t/zADqGnZR7hRIPscaV2vj3lnxbw7re9ZXxv9ASGg8XCao4slCDTNhjHVXcUm0Ut8m0OmKKA0t1K
7x4NajQUW1mi+hhzc8OS48vZbupJFHS5qnH9k52agxLqRe9z44NJfpiVUZN2g5SXIAALUMKXpv0L
3dD70mGZj/WbETGhBWcM1hlQnOdB0yUYUPX4YHu1qZi8TOsmMveEKTgMDH5hzo2WeexuyO4dh+g5
sY85b35lqpJnPD+vK+QUckX/+XHNPadIxDXmLLEyWm4nTu8fT39MyU85T3fcj4M9AM28VQTZH72+
PTtZ07ESokvrU1w+bahrwlosf+Vcutsw83OhCyyU6YhOJ3TUMnURf3VTxgPyLiENZegCa/cFdUJO
PZ9swxzkd3AU880Wf3qnkIx1uZ2Y50LF/86oO4S/qjLpHQsCcC6XzISj8BfW0ytMIrF4kfkRTTMt
UySYMUUhFw2qp8LH+0Au/75/dLLUeOD3B0DYnoSVvTvJziy0JxQdP+NGksQ1NhyJbHvh2VLJvUbp
XojwfvgJKMgklZBSYMg2vD3vX1nBed28bZtcakLj2CU2+Ut+3DGnBdXyYmoKbUQpOnFcxGuzo2vg
Ez2mwvonFwZ6FfCddKWO/HZ1vv2627xl4zGPouhT2dV3zg81BTBzITBQ6CNGZ1meJEvWRzoudnxR
9CUYGDDBO7Eglcrf7pAWndajsS3f8pheJleRITDn9euZ6ZM2qAw75gVi+WmeHyvsXLCtu8MyHxpb
iajesHoi7czQqAXUpjciBT2+sJ/pym5sIQyZ2U12HFQZVxlPxIM4C+8EL8d8HH3FhGm0kcforeU2
IX5Ie3zM93ixV8yb3VoQUHRlHQEtAU1mETrDg988C44QGNy+qck+Zc2362FyRizMVDjLAR6wesG2
nIc34eT0e+2V5meRKmNnVYKl8ZsMCY9DKQE4tVnS+yNSW4030f+G3n7uD9H/HJ8CkAXUCtrFA5zB
Qp4Q3zmUULrRN37/63U1VJyk5891a5ema3Ur83RrWmtBeUA+/SOO0lkPVayCnLZ6V9ktSovYphKd
wRtdzFvomsEvXN4i8pDXqCONRXs8GvQnU0dD/26/3ekQvJ0vGQUju5FLX9kEdEasS7L4snfFTvhw
ZwzkpoVIfwv1HX/l7Celq5brldgW+k304o3219r74M8kMsFOjevXQyl3veh9W2rs//ltVkV9NvjS
X8amh+ACCQTijihHGDZt0OpdxIUgLBxpA5kf2CkqFa6O+/1AVfk69vuOj1GzscPeh9Nlf8BoG7zb
R6oFZbO0prAg6LGQmUUFW0NeIFOZ91OgvK/bRC/ccHjfjR2G9QgXlIrAy0xSlFCX/DdtAu7w7FEo
t+jSaQ8bNPX+eIS1YV1w2Aheh0EMmeBU7pHUw/RaQ4hKz04Q7/l57nVCs/QlyqUvo7Hlbjm0z/8U
olou9I2BO6sgOUrDgdMmeB+tNTCkFQxqyre19zSLyRpXzupeGmTRQJZtAAZFqWurxwCxj+xG6Mvy
O+1KJNh4m93fBGfaF0U2XtXEKGpmQPmzIWyhAUDzfBRRlhOlBnpnzT54WfKL8p/Hc3zSaH3qxWsK
DPoEJbhGpzZIjv6icZJb3ZPL52G4zTju59qkOkkuc5HXChzfBM4qSdVtyV3FHtsp8kUpyhK/h0ks
YGZ3SktsFwq6mN5DMl4amNPEUtZSo93o2nOoVS8zJCFg5JpsIHlIUYM+Fp2pKh5AIkQcdigSdflt
kBGNRT4R9FXoHh9RPQmzH4dz7ezpyI5ujHMyE9Elto6lNZU3wjF25bKKFRrvC/+GN4FNtvq50THD
ufvU1cbgpcEigIH/KoB25dV91EKomRa8RvQczRZvBxDZDNIeZvV4R1Qo/RWKiqJCpT71R8Fg2SW5
cks//CcOBseyxbRMP86SP2JXkC3/TE8GD1Hd1fdmpuyzzves/HL3AZXLSQ4S7mLrhPazXByj+3xl
CQhUWL6VDdNG+H568d2VyTVVfdDOIGcr2454Yz2xlw4KM7yAaKdHjRl7Kz+/ewqsHfwn2dy5ad/5
sD6sh84VgNvRb1+SpIAfd2kqZY1Rza4RvzKrgUgZLSOUuzjX5gXTbnuI+QgBUFv5JKyx/qcXsE4/
iWLD9KlmjIaK2j4pDGgf+q1VJ/9M630NrdUfDd5/uvi+gk/KnkahvDFuR87ydZsDEkwjFTfK8Es4
fTiunUDvdKvtT3aTD8wVtDcTI0ugKy7bni0EeCEvKbOlTefv8CFqIUzzJle7XaAh/7Jg1itTAdit
jjBD+Qf8HRqK6LbDYmY4n2Br666d9vpk6r9o0CiIuVf6/G3H4qEXm4VKY+9iDF+yiEK62ynVAmAT
c/M067lGwsYXL6CGOajvWPLh8rVDbLKWKQe2yPyPTN86b/mQNf+H69PXt+LdyhPFE0AzCvJUROxV
XUPYxqCJfEIEddpJznDNdbRbY/itXxuMlVrMqyG76RYTuroZW/Z33moZvrjqWFTiTFDf0mtRiYxK
GkDTPSIAuORTV+Jal69j7hRB7bMTqv8TB0hKvy/Om5rcYE6cfZHsBTqmL6JTBWhDaq+u5Mi6tF6j
yxd+6yyD+OW3uSkghe1lWdA49J3ZFeyO66KKdtlVdBQeGH+GiDTOz2Z2RfBhvhOjKXFcxOpMxdOB
us653HtnxJJER3BFhDjtc0B0/k2DoTcD6FkWeEJToURy169H/eX1VWYssNgcPCqIW14BkUiBfAaL
kLdsYDPHTqVzHnGjPw72RWPQFzncdNbUMqzCLCW2vH+KXL1CvgBjHMbGynvcV6sbo8/NKMzdbxFn
9P0bot+NbELzkuqxnkd3iAcCT0OjgNvcKHm9ksCpWMiUY3Wl+vkAJnZCd7C0id7TyMi1DOkDGZru
J7r6SdicNqeuDctz4zJgcsz1VbX3UMOKGg0LlG+yvuby+WNiIBE7W+Kp1B0GByFuBjSSU17GsJYC
2byMraenYszgBxEUxq/Yh9nNFlSCnZGv4vZppaGipx2Z+gq06o+FT4NsaLzJl4GKu88DaejzjEd/
MTNddnJcY2nSeX8TkTYZg4JQ/9hOamx01LEolJUci3xXOBKx31YfVhYEzZrCtnBewa1gaqW6lKDC
4SB0WIY0hoYHicRWdFdOotVReo1k3bIqpzny+DnkJoWC5irSE7WqVSg9HXFSz0n96bz6rghkUPKj
rSU/91TdQaefKYN0wl9xt+/rctSQONFSvP+E1xXhr0+THsLdTnETat4OJ1PbAJNqjRM2f4Ec5TYC
ryyVhDyx4+a85NaBeHknsn8gJtbQLHhxjM4o5UX/M2KU/kmDgUT0qwlHyJuOd6hLpk2BTbrVKBCF
cf0bdSAVGuU5hyd4NkvfdocxYpXuK97WuwUFbdIWvSzLUW1Dlc5cwOfAIdoyrHf6krqzMVr0IBk7
gK88kTQqr1c7EA1LpTN+LVh4jI0IeZjTYBFerMjU8/xC8zf1GUjtAD7ERVa4xNxrjJx37bcKK0S8
tTIgqalDufgC5oLDiowbuvNcJ5pgobwwcdLhjRaebfg4fEak2bl/od6hYAdatsDzVHbHD0bTkPAU
ew5Xb9q4dTUHnO+6cVSPEiCjIesJpITqCQujIF8QQLLPY1mNuIuwzQjhtlCFZdP5Gr+f8IwPCPKL
4wg71gatKRVUMhVR7awLMu+mUGcjXRWyPWQpNANnQprytcg3G0zLQgjpxkq1dhsFua6zXgVeinSG
spRvmuv3ZHF1KgkU3oKVKhYCO64ICcf1sySjquWhyHcK3tnJJmFIClpnivW9K/PRdEXYzlEi6xMM
9QHuMaf2PQ+l9wNj+dBkUVOr6kPhmWLuI3/T98uPoIgOTVJ446Pv+1vJq6AzcarG8crJQir/5ENm
HTqElYejuoEpyka9PPRDKoEQibxfB0LsWkB3Ufv5V3070Rh9vf88iZdz9AkxSJUrHITj1qsB7TB5
Q6N7WbbyVrJEEVJiKqgkTNaUSMbRGfwFqTQ4HH4SmSlTg4vDfb5N5+zgNrA+L0tXrgngXtYVcQZv
eDxl6gRcDxQ0j22ITrNiM3/aF3wDdX0ZNo/opWgoZOKbQHOj8TyKXABageBNW/En4CGCTrfPZ7om
SNbRMCGn40HT3PMC9bo6FWb2dRM0G9gyLpbdTQZ93A1usl6Kn8J5f9KdVj9+ERYebqBYPkahNzTi
l+J1OZEyO9vlIPshOLwNf1QWrzVdjAMbWqiu7o7ussn9qPAtn6PmfCkQJHC+bH5jRiT37nH8kyQX
01Z+D/I2106AXyHY9efMQXiV2T9L3Q50PzLtv3AhhhPpSQ8Zxs7bHwMsehVVhs2lrQZGnYMjW3Pa
oLJbSNsnt79CSn9dXCwPs4Lf1h/WDXmAtPwWR9CEc1Tbph1s15lS+O/wrjfyHk99eKbY1JnnQ20X
CahRJtw/hRpOfoNjUXNAC5xuZoe5Wfk7Ja2+HMiTqWm8lwKCiqEc8YZD8hD7hBuwIbvmgJ3B8k1Y
oR0nLjK1BtKOScxT4yNNaHnL1ihkxoljvez8TvWBOc1YNYHK5liNDkXaFQY03A0viLooKeUoWyTw
zuIbrt+AeBdarEkkA4PuuHzldZFEI/hl5r0mA+j73h6Tj1W8XI/eNxmdjYQIgLkixgdbJCZdlrgb
QUdXoUBu8bnQ0HjQ2rHACLwrfMr9FwS6uoD7Y0YVCvUAqtIl1fMbflwZVz+6+vngNXBlZllml6N7
VqFVZ4EPhBlE3MduRqh/gga3n+UK5vdH0HglZgyJGvruOeEJhcxMMg+lj9zyQK4jkvU6LADr3DzY
S8QbP8P/LL+2VxqpUQ49dVkfutjaecfv1xrq+pF3OIfE/R22p5hd23gMQAhQT28oDUjJ0UAMEB6n
2gTvbaGt5Cl3su1Lv/RE2ihKyit1xtumklEbmz8Gl6J6lCW6lLX1oxwJnSZTKLKcE4IdO2csnvZC
EXPZosOdGZj3cAzIYPbgmHq7jrDcr64spQC9I4cDYMUURxFElLA4ip1pu1X17BJbCwZaiAm+E7s4
YA2OXIG2le3wm7h8czuWzRpjPw8LG4vdrC27n7PjktulHif+eMNmukJyCeaBKCuMJkT3nvCmuH86
YkztSVfb/6BBnLgscJLn5GpPeTdsvIKF458BE73ozkzMnnOEXBZabszMO/m1prvRUWAl4nLhfEQ4
6PG1GyApyeR4MCMJ+PrAG3rSqlv1NAF8iPIcR6KX3FwUhOz6pAHkv07KCYboTv2U5mb1hE6J0AfD
Id9fStSG5LBH5pdSH8fafBjXbZ4kgEmIQ+rlUHP/fklvRuDuXixE/mDLnjvlx+7IyHPvVjLTSCkN
kX+8E5jw9ruadFLkV9ly/C2UEi46W/lQlVcNXopTqhEuYZfqdRCpFPBk28I2X6GToeT8RRS/TW4O
jn+a2o9hzh9pqO0r//Y9dM+jviqE5e1SxQwyb6yFY6z83ttUyScOQVTM5GRDbKyNziq7FJKYSJ1h
2W0eQeff4qBX2uipnjLg81gY0p/HTAnCSQK44va8EsiLav3i4EN6TuA9J2lcEgiTuN2sUtVP/grW
qlre/Tl5IKtdtWj627DdaLKXO2VXfRS60oQ+9CuWoT0xPvexGdP81KKVIAdhn7AInzfjfhVX/2ch
o8OMI+QHR89Nl58oNAeDAievGw+GCax3ehaiMFDxLjwX/jpVfkjDuzvauNe29GIKY6DZOkzsrkzy
tm3Yaw6kocvr65Thmv/UTbg8CO4lmNRYpzUbQTA0iNRmvB7qQdSSm1cOzFg+jnzBcSmzvbVjrf5T
M4KFmXPX67mLaqozHyUKu6H50FfejyzKZkUEXmCiDWUlWQU/8cd6Kugj1FGEw8m/xnIJSW+gFb5L
EPPMK6wv6xb9IFno+Q/SQa/z/TX1VD9fV7ad4DxsbKYwNM4RkfWSCr7XqftjaMIAhFD2sKDJCWfi
l6GcXZ9HGGssnnUs7cMRAUO2a5CE5HpC4oAA5nyoYHe44iK2swftXojZ5MlguGjKU2Lwck3zX1ss
fSupGNuWQCLenP8Nm1PJlnWUoxoQXzQ3udJnE0MyDZ4wtEaQ4KaLRBjCG48zkBO0y46jf0ktiRwG
FlRaedySAR3kbOwo2vLwBc6eWOgdcaRWsQ4F8hmOXtZIks+xibgY5mDaEvaGxY/76PRQTzsCPANq
wCGRcln520wPpQugEjCaKNhnPrUUB/Lv/LAtmBAVsS+ACfOHajLiC7al/Bb2/JaTn4HLDHamGO7l
qreY56bkgP7jzNzYEby0cT4rpQpUWyvTLKECQMMFH9SeHjUOqEKdCP/WEsnQW6phUU2iepp8/lQV
z662G6f/KcZryd2Sz/i+0HTC7jKwmHrmImERpiZpbxN3WZihQj/Kyj8EEFIo0tNxs9W7h/RD7wKE
H1WD2Q/6M4okRTOWMPhbZqrjB5sqVjOjGo2tjqw+lgMDRkidVRdo6jDvajVrD62xcMdIPRTaxAwx
4SrEBRRxybLklEyTjK7vlNSv+t6Bf2kEdpq/KrdSwEqiWYO3nYebL9469jWjJ6Iujt3YxX7kS28N
ZzVXHMFkEGQR6xT+v9hMKA2qQymdFz/FbN0ip254xmUeYYUT+isfgAB9QImA11UBzucSXUvIwbzE
K+bBZBL3BIgN2c4r5eJJDam6UZTH/VcKxqO0ePCZUabwfSmo6tSzBh8Apz3PTK4CmnIVbxDpJivi
iawXgkE6DgmJnFxIy93V1Sy4jgun8pymfyq1CyamUKtWiQDHmGn6QI+UAjr76YI7sT3TB2ApzSEf
z3M1vv/BWlsmS+Y7K2Pd9lmmVR1cr+g5JgRcZAHDA+sSUKUQ0yN2wtRKTHUZUjJz63gX0TVxmI6W
r5a+ual8ffhFpzjFQAKi/e+k/eXSOEof8Y7x+wCTptVMXDxqpt0ktKRrHbxFvz4BSLO3fQkIBIi8
ND9756wZ1lD+H4so9fNOV/73Qtc8GezLmVvABcoilU/D4M0ApiJ6pxdK6DW+cTZokNAXpfKpTgHo
rEEAEfu2OzCYpD3hRXvjKv6WXSfLfB91RzPnzwnqSZNK8AWquzEUnR6icXQ/kYeKHCchXOBOlAk6
cSi8m0IB05CDVb1e6PIJ/yDwVSnrRBiMSfpyMn4RoA6NSubNrj/Ju0yYHLpKtcRVUEQi/j0LriyR
3M3EXFv6zAhxVHhqmx2CrJszEYLJmUrH9PEYZG2ZcJOKsLkhPLvwKpGkEpfc5aJlv+9ftl02TMqx
sEPawnkzl/DcD5JtWoZjW5pzbJQR/etpIwPzIO5eyYP2xMjumLoxrJAO1r1T+SREEzbdzwDk9BZ2
GUThErwWHPd2jEU3l+xjzjATUaN/wKhG+xTtULOgP9rz6yzUScg7SUZXGSBO+vL/mvjIdFE7WO/B
50OGkewUFb2hoIC1hyEz/nX19GO82IObLwsfGS2ezTFpyqn1hFrpDDl8LSexo8JHnttcim3LQ0zT
Cva6g6n2vSLdh4F9eb1MiBWMXaSfpRvchaE5aJ/y0B7w9nZiDOaI1qcUGBXTKlR+E0QV4IZc1ymX
w5HmxCTwfWZHlsnYFd5Z7SsmuLSbBCtA08PDEFCcteeS84vVc1hBi2A51ZHIKL9nFOySZHfZ9PE0
ReWIOncCxFzLPwq6enG4IyV/1ydRWNVko7/0Rs0VTg8vM8qkqRvECoiLjCG+A1ErXEOpPsq+t85I
V9eiWP3oPF+INidkyL/zZ4/MuO1pXWDlYeH+Z3ecyoBjw4AUZLyHajdSq2usMW03WYlPvslQMoPK
J8Ung55mCStQ5rPEIjIyWlETxBXnJ3ZDrcwXS9JCiPxQFMwAl18YpHJHbzChIirkbBM2loGGSjDl
YoEgULCQiugGB8nhmQfA5l9Inv4odMW6W+bK8UinGNp4FVA4aOAbiYTWnSszu9jaG2fAS1KMLJPJ
gPZpIlWeJ+FczFaC7YMHmtHfqrbEManfHVp1B+WgM7tJBSc9oGydWDZ8STDed49d0sIJzH7+50/r
frKFFKb/9++9tBlo189VbddJohzIKeYCM6UhpQ8P5ANghuNtm1cMT9kIOAEGDsMBtlAQAcAR/sDn
q7TCC7JQ/UGUTNPs9KwpVLXejXzX9o5EJodj2pXEknZd7G4eJSuj+r9tqRpOo0lm7ZktA3Stp2Bo
T73yQShm+a6X2ZxK7yxGdr5JmVkQRaqrTMDH82oeohK+U5zNlXQSRmyzNqf+0ObZ+6IHNr+nyp0f
b2Q1U6nClw3zPWHo+UwxUSwlCsK3ejWKxBiLvgI/d10kz5phd/wMO72Q+a0/WLOU05D0Ne+rEtgD
71QxAZOYa3HGJ/7/36ipyKzN82MOydE2wChpfbT44mNNTWK997IOlPTmjyGTNg8tv9iK8YmTtFYV
TLfkJKwROy1oI29IRC3XKyUaKhS/OIphsFI4MdguIxESeZzQnc+eudXD70vOGHLdGiSkWO7fvXln
sMBn0ZtfV8xBrRItf7tJaDKDI6sLh8/DipQXRMTodZZmyFMISXN/pIHBroZhBYexH07+HC6FX6Li
UfmAoX13VapVAWuUMX567JUXcOIC5hNF255A11ZyrlwojL73Dqc5qHHNSZVLQd6o8PpfbZsGVhwz
FQ7wQdDhT3R/o9Mt3EYWUdpk7t/dSZGCWwIvBgsxjTS7L2Se0FW2etERZrBit62ul83abMN4Ykc8
SOnZTnsFc+Db0RDSPkkDeu49/gmAt/jllw+oUFNMYSyS7HeeCYV5otE1rLIrRHDkgKc4mES4VbGh
CLUZeDo6LthB6VbYU7tOHqLdsiuHOURG+G4jH+29iH7JPuhO7bj60tpFer8EOKB0xeyfMdKG+zmu
85hQNhzPiSpM8XgX5e63h7J2Pto7O7bhObTyKtzSroctbv/yQ9cvBK1nBftgsk8NF+xPlP+Ny7JQ
Gwm0i93sksbHYj1fYswZhgRCPRDc2q8BHlkdcLTc7o/k5U9397vx72AlHO37UHSfjB/JVkcXKDx3
IOySJ7PXj/1taYct/J0OZ5cucoupWPnYS6jqPbcDe82pIzeqwnw0dPLAiYA+u9LfaCR9QVWkvTnL
e5wj4HiUX+lcDKDbQgiQMZzZRxzdyyv0AhMPapokXQIs5yogSBf+gHFXTJLMLUqUqd6rMIPbgMdK
7tBevklCsvri2V7OQZqbTjU87DweezgtIXGm3iHoli4+IDj6efmn781oRIxjW8uF4DoCTyjZ1q5x
hPQdKm6bU5DMW7wDm21ZIqSg5i272AWJgQtk4Hhkwfy5GtETUasFN2ON7KUNQM6rcI5D52rzMFsm
8XzvB6C3NkWjpLSsKN64oZo4Jvx2AlhrTGII8R6vBsF8Dk3eqYZFDAJfeoA3D2GzWsgGCxDfLo/d
GyPDKxYqr5FB89nuEzeV03Zad1wW1xCwOvpjHKeOfqf4EXKyP2cxbfPUob0qJ0c5J+eeuRAx4i7c
qzkNZdT0dh0FCtVmzG1eChas1Te9WmdpmHCjjePdbQK2iuMxmuRzx795WF2P9iuj3DfYEp2BvixA
7uGTWxfGfXi6c4VIDkTsYbUn2FHuOqS7ij54m+EhcU/UTexUnhQ4DkwbHDxYaVcV5uAw+W1QrwQB
H3vbh2TtyjNrxmakA/OxvVXXPVm1l5/MS/PWJvoqCBJveCqNZ4GjJ8a/r2I9ZgFK7Wj25b7Tq/Mp
r3YA6IxroHoEVjfBcduB9ofIXmGf0leMf1nv0+dmzqNa4HOz9VSmH5HnlbXk+Kf/XfEnGhMd2/s3
QXRgbLm6NWn8EpWhbGNabaNkOE1qBGDMLRtacquWoLXjL1h8aFlB6ewqRPdTA2065HcILElC5I00
mcm+0NfsWiXB3HlSrRC82Sh5YprATicc4Txqnxb2cCrp775KNTkmxK7ilNp8GjT315zW/pmVFs1R
dSpPAF89r1dXqMfNWq8UBY8BLovA9qa30/iUC0FuIYpZL1YzIHvb0TgLsPE5yKqUXOT6g/ijj5RH
QNe2S+KkGQgPZEMgO62Onj+E0srhleWCpGhK9uK9UfhxTg7Nsxv3izimd2iF9xcVbM4PsJYOdBsp
Y4trrCqHzngvZTrr0LfRR8zxyf7mJte48UmL5CFWWGdb2I4vIdppVXzHlfHBMKfYkjod9Je9uIdG
M2FWt6ZTJ17q0aEmRcSPxDgdim80/3uEHP81/t9wH+OSLOqY5r/hIADJGQOs6uXWB3G8z36gLmVa
PHU9b9vIFvyCRetCpRHblntFXF5oRD/3tiSVgOmATrejBPTDcS5MGifeTtKBcyDLQAd7y+boC2/2
ZWziqw0zQnv5qbtZUJew707V9B1rtdR4dJbSN3khrP8Aem8Ww2X73oUhzMtJt5cYciCmrhcTwD8f
lntNPla21DC6yL0veV+kxQQAj9SIECP5mOWHg1ymKUp4xN3V28tvHvTMSaI46j/alJ9G1uqb2VWo
1lSD3dItQLCSuPMB5miZJMuO2Y2by8cg18Q8DR65DfPD76c1K4Eh0TscnjKI73czHX326K+Nw8Wd
eqFxbB5kw+vkAQEfKpQHJeeOGi2/5pez4ZsaPEiGEDxglYfMJvwmOMi16ODxLQIUCs8BT6fl/bR0
dZ9mqNKe815bEcDR5a/4UDd2JkwhEyAjbR3wJ3WseTgrfX3khmCFGKIFWGFWk1X3YEU1cX8LAVJg
Qk5CZdLwdDcvhhOLoPWQEM318IRiwGKOC/lPhLCdYsSrtkwhAPSsRCZI8GRDdTklVnHI/jk210N2
upanHY+7n8Gk0qWk+WPDsifunAqZeg9SeaymVXPteqRbu5PxDscQuzG/MncJ478VntvnVuzrP0zD
fSe94EvOXGYGSu3qaT00HmvhydqFm5E8X6jwxdMPvkNmctnRrI84myIaqz8gxG56WDErq8a2Ay37
pHAx+u0yreOqMneg0Adcdivr5c2qM44NpsZmg0E6KOReyWlWguLe3ZdIhGDX17gEQpi1oDyhCCDc
mQbN9D8jn4d5tkpJ21fjtvZhOlruZhac+GRi7D+Oz9/fobkCsHjkyZmCD+mqOvFwgZ+olXF7jbH3
VzodOrgIom/aSC5hjZbTUVue5a1B8qJXwAmxvdhghCC2gA6iW366Hl7rCKEPKyZlAEKUVDy8MVVR
eHE2dO+QxdgyBLbCvQgcEcRFMEnK8PxtZM9DECZdaczG9PvgUHfBFa8ITJdxr8VY2cOE4+JdrkAd
2xTUwfz25s5NHCHeJxC7nfhFa90inxWiAhmBdbwwQLCEN7cA4x7honkZSBttOTQNh6dqsUDLqwjk
fz/LXeR2kKqoLHAi2Wn9VJ2Kl93EJ/HJAk41BNq7mIUI7VuH+6EEfH28NFUzJOLhTER+JcEEAF6+
afOY/Je9+h7Dkg9GD5YX+lkQ5AXHfuQNVe3Uy1cKmrE+3fGPRxSayOFzLM7b+x2dyM/juqPqJSuQ
hBKvba3QK8jLpj6ajF+eiwjLZ04HLSIsN+0gWw6ttJr99Sr4xKtFdf926bcPVSeHgpxRksMhOLwA
FoTNzTWLIL1xXNdjMJ6CuC+sNYHOXLEVYtPckTuxKUK9HBkDIB+y78SlAKBCddA2HdX1ewdm7F95
Fr1NuBeZ4uf+QlqdroPU7ed7Fzq+7dIsWs3LkDV4PKJCuxjhjxn5TpDra1YwjW67OaVHFEpcGpnv
au4JmRFxG06jn6jk0FJQS9eqbIt+AZy9jF0qnHL4mOYC4WfAdfEQrp3QdxJMSOwxCZyhUgPCxwVg
fA4vN3aL6d3PzHCEsu/K2hWrt0V3fIv91PN8jsnjdIxtuI40ZtDUfEC1/XClGX24WqMEKW6LKyjH
6tldZKjnabj3MnRWt9pZnfLW4qTR9YD0SZ+bdwqC0xMqhqa+kZe4iz1NHtvGC3pecGpOShZpeMIK
sf6zwrCktC1HQoxVgSLHj8KK2PjeOgxnrXnOYGihsUvceHY63DWTy0sNe43tAHa8yvN9pD06O98j
t6qPXAf88CzsGQpaZi+tfZK8fGfFn4iDSF8cD2lDmmiVL4qRAs8zkzOSGGjQyDD6SqusfUad2oWS
KXq9v+G7k1r/smNgfZebhKntFVUxGMPC3UvrjeViVzJeSddv4mXoXLykBR/LwDfCgoDsdr8M0NCe
M2WefMQjXnFKnqtJ5W0EbvtkivMY63HHfZkQa8lIRgJ75l+VziJaLOW+n4Uo+Ncz6k9VpF+3f0lg
h36/nE4nuYBZRfAbxgMCPq23attDTTuTnP9dcZkyE7UORpvTYlll+eCC4cAd4Joq5DJBzoooaLns
swyMWeFKCYwlXLmb9pveKnqZ7UJSpCJeF60C75hm3rFAZcGf12yCMnkKW1iftwbj241SKgPv/3mJ
INB03ap6nIzVmxfC98GgT8zs1zL05jZ96KZU4cHXtzYWXc6onQylyWWH7B67wrg47H+SbWhDSgvs
ZfparUT9VDS7U9kOs9jBkosZFPhAx0jzVLZWCLQQyWXL8u1Mkgy3TLdwT6FE1tBdZIl3DhEvZ5bD
X3wp0czyVC2pb1u+UBwdpK1mTcbmNTQyGgp2zsb/9vNlQpc3hUsoZH6oi7zSlexl8ClbeCu2G7mw
AmUImmXS55KBCzpQsWQl9e2nJ9seEQWA9LzTUAar2LcEbu5BSot3c+6DJJ8w1rFeFADF0avrgs4q
z+5MdQyRMuD9s2EXTFRqiOd/Dvy1BOKzZMP1C3I0gbm0II0HxYV46BsMhG8OS2IpzdH9iQJhdj9H
BqYzKvzrMk3ReytOt1X29mHmV2chmy7tAiHAty1voAZSBBIeuAJ5Ng1++CVo3K8e2H/4P07CTEeR
KHrw2HPp2lLvNkzIuAIocBWz7KmIOAp9JaSyV2ju8uS5R+fmlaDgtVM2b82/bCr0ymWXWflyDYUW
xZDw0zZp+yG4NmYpBEAcd+biF1w/4MytpYG+FEy8s4BEbIXlylJJ3YWeH9bawUnPUaLi9tsJp110
rI7kS6m+AvSxuOm5v1Gzdx+IDpOGWKwxavnqfXkkp/ww+LR7jYIx+kHiMBSir+FCw2160wrnQ6Jm
kB0RcUKQTl/VpdqGJRBz3dOqPi2vQo7uF9EeYO2QJrpPgmoqBUw8L3z8FeuITyGK4ZgIlHnUWTcN
CrCqmjBccy4wdJQqd+JgKA/nBCLhEqfqkWkuQ6Se7P5THhnPuQ4ICGvB0/TVRG76ar0XIdJzrCid
3IZcQSmvnH7Gh31YmKrv0wVD9nXSEaFya04Pfj1Lcxaabo2rrvWORhwotF/ZEYINhFnYG1Q+OgDB
Ns3xaF14wH/Gv3l8JkCIX76UQzGynFk3HpZgOQFJeqVkU+CUfo3xjOYahzoMuO9JBjrAmJtEjExz
cpoanp/7fMr1mpYRe7ELlueCGzgTKZlifGEhI7stbTWjLBgOV0iOdp98I6EpLZxetCLLH9NOs0uW
0zjYMEOsUVitPcjeTB7hwc5Q+rZfND6EZc677aTbQky/XvnHmvLhIfHFJIonpAigaEikZbBlQzP8
hEjUiNmNtOa9amN0C+oM3L7nw2NDqVgzjNjxTVfzcOxRTI50vk4Q6muvSGyjfrkrBehk1ax8edMb
Xn2kJAnyCuNn3WNlC6xRLKvUwOaE5JfVSUEoNvk/YUhIrLulNHMAap8kMDuQVJTxPyLadidAaWuR
vu3FHJkOIeP3IrK6RKyb2pT2FJtWHVvps2Gyt7AB0FOjWjII9+X4VUNkVkDM+f29lvoEAMhfmuHU
GsUnl5IBaj/xrgTqYBas75AXcx5EKOf7f1nQ3/RyJ9R89FrpU1j+zrfvzlUY2nWRQ6a364hlnOlc
zQMFc9JVEzABps71oGbfOTW5JjA2du5Ugngjd7OlkwdSKZag3kyOq4V40jBJmtZSFjzbP525+7uo
/YRGDO3TFTB012++09Bqx9IjPQW9hNSJrVFK3Hdf8mEgDi8oDaLdnH+UryNyz0XTZ7t2o9L8xsSM
aXC6Ac5f1BWUB7ngP4z0y4LNIsByH0MIAkkHFaDYOQ0dVz4ma3lzwhdU3cRAebpXfkDEGqSz/7Cm
83Tycrlr49e3ShC0nElCpKaveMsIMJAfOb8ARwsen0Du9iKEHugp4xH8QI5pxwm1aa8EaUvVRM2C
UE9i6t9jPZhdUBA9E0h3k2K6ze1ljHzu+tVKEO2cSW4Scloucwf/lY+2Y0/2ccm5BgZn9f5ubvPc
/OXviRMfPbkBkLHDRh8GW6JEvyZzYnIz5TqnXxIY5HQi/dwdOVsyOW89w/fiAv3FVA4sjpCloQ/f
goGoNFgO4LXgew6BZJ7ZZ/583ozCQGYhwQTEGXv2hvEKXGJoJz4Abfyp4NEqMj5AbIMSprc2htBS
mTZ3NQJcyC2SJh1zVdkUc0dG9s0rGHLXD3j2OKvx8iUCqOF8mXIsLKiXs6pJFhCOu6G6rZwCk5Kr
yPHomPp14OvOxlNCVUyhQ6ndd9Mxk5RyyjYTRLn5Gi7ICL6CJoQTt2+jybc9RnsfENcAh+0TYkDv
HD6vTyDQ18v7ccuROnwFrr0/WZHRtWffP/ZWuR+satZ8egKMkqHrMAh2umVAeHOm0LORNCWcjQ6x
I7Xd2h4C5jFxe3T9ob6xhlyrmQ1R1UoPvhLWrDeA5AY0bTuuEcj51/VXSphWHnqVOFtqOQ1UbSKR
7XdibEFrCMkCKQ8B+skmpYVyJ/K4fB52xNSLKyN2pEXtnoRIKlqRYWftdPxM9z4Xn6FAUwFEVxR2
laO2YDOC8aeHjPrhMucYskak1ii8itulKG9iVNI+FOQYRfeHaW1/n6UVodwGq8ZGXvBjFDH4HMJh
RkhMxd45xufkuc6z6yqhh0GzxTomStOtplmz4+nrZkm/k+DDeUJnb0IzjoR5MRLgVb4avBZm4Fi2
XeDidO0CsF2vM5KHkm2ngwiNGHLcn6onUv1j5CTaYcYdPIbB44CXSdUv1Nb/P/dI9rxjCx/B/r81
zFuj9h5o3EexMHyEUQjpGKanmMOuwBVdwTAMSIpLhGmPLRoFvxrSgsj7gRJ614kBQJMWG28PnOoj
s4lWBLUVn9Ric+aSoU0N4HGE9KSWlitPPGldI6I6slTddVWqVmqWqIWbLvtsbThm5tnIw3kZ7NcX
TLUCMQOVW/09oRpckMeNtPq70wPfLvBIOZnzYiXEOPAK1ghu+d5vvtsUABJSnMZP0+bPsLkmnhf8
Zjzo3GidRe0NPJsxeCNl3PRAxFSEdC2taGnnpMUv/J9GubfVPXwsxC4jzrtqT4hTYkX4keOHenSJ
b9V5uhk9ncoXNUIYICf3+Ve7VV9S8/79inpZVes+OKhNh0D/+c1qcLc+yT7n+yBBAdGgwmq+5mku
kgkvn9vqgABcXSz8Eb73euJSVRNP6hBrcghNLNoOwnwIZ3EcATAJHA8NYsjyPTAgFLETwtBePJSt
sm6LN4etD9nsexzqAjOmKd6++V036RctsNrDcWO+1ldWDM5Ow8RM8Sf7h4nANrRBKOuGhSQkffrq
lheiLLOnjgX88OUW1Vk0gTiSA68oZ+vzunKP5dV8xbR6/NwpdNmEcrah4pfTT0i0eBjSm+PYFVEr
cJl3umkq7HfqwqhnidPBuCcF/NKpjqOvBgnuJdT1/5Lxb+iquQtIac70zCVyflIEFZg+DMuQZW3N
+7xvLnf7lF+sgyR0t3y1zCI2qD0wGSmr123mnvtzTNephfTCWHE0SOGGL8pH4LIwnaXqqUHTSrZm
yPcnc1EpTlN47CvVMNee4ao3ZhyZJh6g3zkwmvCFt5eD8In3yDJsAUbLxSE5nYCXYmQSvjyGSDr2
u5OZ3v4nXp68JoN6m1i9uGZtqT8W3kXdYUSxV8V6AStnOsqDJjf3gfO2k5DX1tWnIuyisnt7qm/I
1enL5fbbx8pyTd5HYxlOhOLy8tlMoBQnuNj2R/A+D8CG//QMK+tx2vz4gAv+L2SvMet6nXr1yQjE
T/nv5YCDNfZqpLJEHqA1/2XgtSGGySN2ALRjWQA7eomOlWEPa5INQbKASanWA6xzHs+OTJ9Au4Dz
m180ClKVniP//C0H2/WjBpeCSNv6nuXk9tFMpKE3grOYYrcJfbVgFcDO+wOweu0w3dLIRsK5iZ5U
C/KCea2VE8WnyzaI1jphCv0/8newo13YUGS+zUljmtJO0Q4UtQ+tFIt9O86kAFjNCLwUCXNplB6S
F/cHNMMlwA1inimY/jMoZugpVRFJL0YorxX801NdciDaPe0W8FTxOa9YqXGqtte2BScQdfsEbbiv
FEJLv+M20LX5X/3uS/8oQnHT7yzj1y32wsdvwuJl2KRG0//WA2gucmlv8/cKtZWEnVvhm5+AUUiF
tI82os3gVEKSAmdSGuaNyE3kLVZanz3S+sYnxlrbyQ9mXlajHA39J5V7yoqaUtAoeZ7NMzmrHXmx
QpOsm6zZS35xqhdK5VoQWCjS+eAXPxIFKn+o21xPg1d3LcdQ61wUkQxIXxjJXh7hyFafOFe8lxoe
2Nmbf9tzP1pGiJ8uYkvegNBXopdVLe7zROtHLUXOgH1djcbY+75U2Pf8omlhLhFMY4ex5qhlkd3X
aJ1A2n0d+Cc3zW6UX08vkOd9u4D32sqdESwP2Z392XatTeUhE547QQKefMNQxPxtkWLGdO6T0nc9
DVBnuVxvLftBellfa01HhKUrzGzZzIBRbVGxTtpR+dDqo2Tiwj0/UyNxVjBk9czxu87VByxn4scG
uLov7S4xI90f+qwyRwafCgG3NvmjnFjp7EtLFAVn+w9qQtZdvX22COo+y/WJI8Dfkimk+DT6aVuA
jH97BGSVws5Coe6qcrcIXzhNMHzK/AZUISry60S0s3ewv8ba4yhjr919hpeMBs8aD+fPVzBPIk+8
Qbtw7v20SLsJMvmt8VnFzjf265abbrJlgeyqPPlmTwRIaZlLCAxf9tu1ZBKSs/a0ymXfOVd8fpaR
AIpInvZcSUJgCRWBQP4wlZMYrbnXIFSWi3WIPmp/q6+zwt263OvcS00+esW0BcsDTqDynp7pduAV
HlqJF6g/rgx/RpGQWB1c6elcEcg8e3k8125sFeucVwIL6RteawCOIsCRWQkt9ED/vXz7TN/GIrcs
lBJIuc0jAG2ONY81rLVF8XQWU142s9yoLJu9MlXMfUV3wqnJK00dIO64vNOf5MjlFoMG1OkxohB9
0BgeYD+4hmQvu9vaSvNwRMSo3tyvaYON5Jg7AxNKjpbotbdfCWo1SqHgGMHyfj2kQPpIKPTvIvXU
PwfFPEiF4gbADN8CZMiA2LkCPgt9rN6O3KdiXqRwIASHe8YoB/fwLpsF95DpNdPpBx60CbBJXl5d
beBamAfgoWr3R+F/gLfU2kykkdi/2d0jm1qJbXGu7F8EyVPr3IX8ziE7hRftlT2Ob0wqrvM4Pq9d
s7OCRd8H3xX5ctuRZqrmmWrzpz1WZUuUtkmQcOlnEP+TvDva2e54uhKhow0WD+4mG2vWafsM7kDg
y2FOF6E3G/kI56HuqzAOB0NKxM+wiXkezjvxwCRzr9QGnakgQI9Z4Kuh7mY6rWh/H/3whxUyTVPW
rMlittQIiUVfBGqK3d6NR64iDv3YUi6xWUiixixxsIsMgAujZwUfeK7YimYneImtaDR7KDyeBYAy
eE3SFvz0RK+RRa2QUO77xF3XE85bw/yvymdwsGdKLPXjaQeuXisEwxMjz2rlujUgiLoAghP4wzTw
F686mXByhR4L9dyEDZXOpQZDR+pkrlKjKuipSPLymYVGz6mT3XspaSv+2CaEOidpP+ggXPCXRHfF
9togt4LRS2ZBYNAwrKM+Tpyp7Zcir+TYxyuBn0PWeIOzXmK1If9YpR04tAIMth7FvgXuxktZEFTy
DYW7D9FpjdcqHBqHC8FGmPvGkHOhYUZlm8J4WNoXkF+6HdutJauu3c+KGf8vTDXkyIOp5N7LqOhJ
TE8s4Iym5uWOdfDQ4BEw5JMvrZLPRVw7hy4HGGC3LzDgZPRxnIRaF/CyWukOCm4FBE7dhFaoBaHw
WQ2tj/XGIhf7n9guvDp23mDjOvK9md86qX6wTnBjbOZocCOn4JpUE1fPphbf8TP2U8/5jmneMG/3
wCgZTxU8mdxZJugeSf0U9+oyr2ujOQVjtWmASPgPjF2WZye7zuj5iTxyei5Es9SSVKFdxd3Ojiox
lIE+UZt3RSIIlJ9TzGX/1IdYnwCKhJ3iYUeOcehpbx0OOr4idQ9d2YonwuVELLmO4tOH9YA+16AI
FU7f0cFyiQn4YfuTc7M1EO1T0L/ri09y8BK6xoYAweeduHSL27fJxz+gU5X4yBBDpvSlSVfxiEdt
s0TeNlKMNiZA8+xEQHGSZRQaZ91mHuh3kd1uSzITh4q7QZMYmmS5JaweH1NJ5tpfD9XGRyrZtixL
h0K9JRhjRgwtED6HJOU8JWL9lIL9SRN8W/u2zR50Te5IJowHCjANk//YaniqQKNkX7NKjIX3DdGD
7wdFhuDB4907JYB4nHIemeFknr2tYKj2XU6RM8QklCat5Bo3gpFhRPBlkjEwzlHdgcgyXtOl2vy0
hmi0iKTf5VeKKZIoIfh4DiYsprYi7W4w3zQTz7UOEGHexb8YOjf3lX4bmYwhZIdaYSIz/XIvbOrv
1GenPp4ka9kN+6sjlmj3ZmPQHPDpMCW7b29qklPFAdIu2QTLAReA5y3TTANDopbD/V1nCjv3+siw
m5WllbXGwt8yuHNr4gzTIJyhLa5OReToVgMsxjvz+0AmysXmhEH+PMDIRhUB+hkGH8E851UxHvcN
ePhi2tNJkak3AoWdGjYlrB7HAEL6cwGkaG14uzechIzu1b46GlQaDtDTR+FihBp5c4RdlyohY091
2TwVCuafUjdBlCCYZ4wnmPn9qVWeMeLn45rxjwPMLDI7C4MlQqcO7e6Mh7p6oilsHCkmYyy7Nb2N
FJdQHYIof1GkT2+9eu1nwwVTRD/7Bk9L56CJX1kGyLGpIgsAFa7i2dDL0tzxfbjMOyIw3C8ezoey
MbCqrI3nNY+9pgZdxRsKRab3v6ZEe+p70dkRJN+XnFXl4NFLMsc3gHW1Q3zI3c5lgNbH0BqAUuCm
mmU8CDnwO94H66ELrkfdaBqUTDC36oIFkowPFfylxjtreF9kLclyxxidgh2drrgZ50Xo56u7S7mA
1r2X7eQ0ccW7zZ0XNyckhM9TTdCNiJqqxst7oEdEhr2sQ7oAQfj8CrqyhXuL3gUjQL9H5Bpj7lVH
O/3U1i+cT9ACJ1Ttmhzo6j2wCWBZ1OEDkyjpyIKP1Sm1g4cMV1mxmcipemjoxlGMtnYqldmSUtQL
ja7nzuN5fHAqMkQATWns5r+P9Dkr68Zq7bqcctq5K28EZ3TE+y6L0vS0pv862NTD861wGh7w6f12
DyGj8hZvA7ygQezb2VsBVagPPULoh+u/Kv9Icq93V27ZirOEUv+V95n8om9WTC7jPZ9s/bsmK6Hm
8KA141R1mpx4c86hk1YYE+BD54RW3Ikb28yKlqi7hVPSHGqBzQ2r8oXnIc7SEGh/tgmExYZOTcAH
Q/qH9Wamnd75CSHvuguB+GcT80NDtCq10MSt4mfwOBM1L+KeCvPh005z+jOXqIlPOGszBk/nzz3N
MBnEoyKRYJ01xgWqyrvNg4tWafTzCn9/HnaP9JXGFZRJ/lzPkBtT2IwR1fYF8iocV5AAhMBmW/sO
+ya0iFekFhN1ySm+9c30dtbxVg2F7QI5ePM6n/t3pUbNQhSh1YabfUM6hk/IRK0x5bXdCu0OF+/X
QRVnmAbzY9qTFDyhl9sK4mvW0dhMnivv6rMj4VkOTJqdRHhgynLjhAuBTlp4SEdFO/LOvrJ1m9LJ
mgiAV39M7S9bT3kR9xUvSvPAPRDxFzI0I1G8S0XtGj04JSj/LhmtAvQQ4YuAnDLmxcN+twVWFeZK
oDmB6EIjPJa1BnLBmNVt7iiufgw3edZkMD0Ohw9vvw7noztL1HvW1deIs3p/ra/Zhu5XMquYXeOq
jHnOS4Sx5vN+QaRCd6HYhSWSnhCSUuxklbKnXwmN8zNQvHlM4n3DeQXocpsMnpw/pwVFcGmHyWJe
2+Se4JoqD+ZurXhFi/qYH+cYHr3U7RSJ4EdCDD1b5J0V6r4idndjRm/nU9V8QVhUwUK9Y3cVf3Js
SabakytfX46zWW1iXFdXNhJfM+REuHidXVDgz68ZYegByaMIlqqWOSLYnxBLYlVlslJYUb4/yVw9
J7Ln/jAjT5/Mv45kQJ/vXW/wMBJpAfWF5T9ehEQVdUCNl7U6DxprwsTNtYZnPf7U3CQMPCbFS2uJ
gr0+Hby+neRD3dLYxVYnzrFtqftKdKJSQiy5e2Y9pz93Cv/UDYjuIIlf4RcEw6VeuMiUrvLkdEzA
ekao/hYYh61KmarOgPinm0riJ/ycZc8QC2mnyZadC4WzZEWSnhv2U5cBxNMjwW+ylegDsj+rQyht
8iB3ifSjqzNlWA/RcRNrM3sFuW0DLLzKFTx/XhrIb/byLLWE0bVKM5dv78zCAlaqz9sftSuKI6Hl
iBR1GiL8EERH8xXo7CvhUzky5Sx6BpbPuMW8HmriIWe03OAyGAVYkASvi48t1cUUMkbcxuAG7lQI
l5/UhNhgrx6Ak0v9NciYx/AyMLSRfTM8AqhMHzP00V+RVpwVN9SMSIN4gX1GSX+3UU5avD7yVHy5
hauJu8F1VQG5OFwxz4VK+sypDiEJTvpzDSwQjMwFWJyXGo5sSh+SmC5j4MBWauPPTv3hwAzavlrv
OdMoshCYInKJGEaZ7W/+oUnCjHt5OR4BfcCvkfn/FqZpCQo66f8MKZu2AsHyTvUgOnMHGzOF+7Rv
DlVlGNPgBWjYIerr0MF0l0PVgwRpXoewV4SP97TiwA66RDt3hwV41EZjWcTiNEDe/Bv49tYyWlCj
RbeWJtIsEYpiJ6q7OnFv833lFbKqwJArmzKtnqfG04DbtxUW6YNN3xrb/mJrH0Da20cixWC+JF+u
a93MJ6dk/yC6M0+10T4UXrzLNh2pQVmOOGRnLVmR/P5Zr9Jpt+LrY1f/OV3oDUysksZjQkKM/Bma
QTvRfD3Ej7QSnhpC+k/yefPe37P3PCw8vyntlnKvUFi/26LQLXdQw+g2msMa8db55JWHgtembkS/
OcOJf5OQT0KY1I8ZMuKSNpjdL0ON8W9rv3KmJngfd3sdYmejvswjPQV8IXEjGFfGDkHUv3/cZICf
AD9UHWeiBw2Z4u+6N8ryOt78c1Sab9I6rxpXKCkGgmMUbZ1TA56k0bHjOJVM8tudCl+fa847CI6W
w6CSODvQ5LhwMm2XH/DAvTV1KLaypFwSO3Lk/0TQvJdONMthIdQ3MRPc6vKXcY9dS2qJmQxylTZW
UXvs+Xcn+Dp9uKqngRp+XPPD5Nwutwvb9Ub2wWapxhpsSADmaX5z6lBgMejGTy9wFVmIVFgu1eA8
mnK3V7ehIkKgD0I+mg1FQZmF8l4s9BrCuydmXpacJmnvp1y5c0+aX9CTyr3yZfphzOxZDTAdccga
Vm969sJGqHB7EQ3VAEQNJEuer7FXSnYrPrKnsT0YfZd8hSwYdZ3zjtoAp2elg+IGHoDtTELuFrXA
+NWWGGjNg91kMieTnhKct0hdAd8hCzNLhfa/FoSIMptnHMfwMaStrspCNs2576rHIwiDQAK8FDSP
Sz1m3ga9YJyHbZClH5oFLkKZt07pvpZEc0xjJT1m/2podHK3fognShruXK+sjY3nKwtQb8kjFm8V
epnrG7UFmnH7RNc6gZGvDEQS3C9kCMOSN34a7GsqOmKV5DmOmtexROuXxPLncRM19p/ul9eH+ZZQ
nqMMDOic/50wDN8DDpHJHrqWhq1nKfvrMcHXla8u7A87XwwRXnHDk3uwp8zB+6BIXwBYsICEmPqb
zc3PS3aQQVgAhaGeM4LTRSDgEp5NSGjq8um+vU1T8j0/4FnZHcaA0JizP/RmvUtDiEkB1cWjosYQ
zkAMEFHSvwhihjKExXspwt6GK4+qhIHud+rJtCuGciG1HqrsP5wuT63LvFCCphg5lGQjDFQTBNoK
JaOyDI0/caTEPK7fIVw/lwjWN71CMMm4gkjkUixEjb+uNiOv3EJTwV8YQBL8pwAwTmHIc5p1lk1/
pxAqat9ipqBMDN8ydMArJbVKZ+UoN3C1dpo1E5N8b85fS2niq/xDubsHNREa5dBwML4fxbawEQSZ
6cJUP8gdHB4l2dLKBlCqWIoTuxAnmX4CtjvYPop2w5FNhA3825w6af4qjYGZO0MqZEi3oEvkIg4B
NZId5+9EEf0UuukuXVtnlsGhsZppfl7pFugicPBTyEZAVHCkKC/4FAbUhx35L+PCPMYAcIwiwMA7
KNaBM/uElW0yr6yOlB8RW78xY0BbKmhzYyd8KN3A/GUoquyLvo62WNwvwgwmxmL5rpZq1F9pzynm
EKQuclKGLGgTSxwSgfnNq+lW4f/9x/T3TNenNgODFiWDQpPQAiFH6I5Nr2ZQw7h/YaQFREpYwPfw
BBioOv7fgEh/RNpwY4LBQxrkcdJSi3BGYayVzYmLk42WULeHkdsh98gln6nwa7yklvsdr4FtTh3Z
Drqc36qreA9XhS2rlETIB3e6iIXFaYBAracYVUzYOAfIo9cDHNtkq/K6EF6ukSiA8FruVsh3rPYT
vNZ4Ai9bJNeO9r5ncNyfZqG7rgAf+r2sraTyCkG/yZy3MIVLmC+Q3vT/PO6rFB8vAt5nslCC9HZw
UPSSYRmGc0hCv6SiEApEYd5uEws1vRj6qSTe+v/VPqMCjmVPHfs9K0Nvm6Fs9rye2OI0hsIJ2U6f
STd1+6ZrU6vrKevZP3ioC1iRYtxnnj3Z0U6coWshgVyxvWC/7uZD0nsiXmtRp+6Pvm+52xVlKpfz
4u513oV7iGnOZV9JWCiSVp8pntpCArbf+SvL9ZBHtGWEESgQOIpg1R5PyMSerl+5aFs9cHysHSiy
JmBUPlsFiBbi/Pnb8B9F4bD0ksQG92VmAiSweMB80yuxSE+xZ3u4DjC/Og271CWc8I8QkPB/sbB/
CuTVMg8fI+yNR/bFZuGONRGou679tWzaA8yFWrJZvv317biHRgTluWzu3lhbaLTOLlbDRlW6tjnA
ksFc/fAB81cjitYiGjmiLsAsTTeSupFfR3NTQeGOWFusKt0f0fT5C2WdTHG4TWuMFNKnD8hRNTSL
KzqSR32rJQ+Z9DzGz6GAMdXBnBM5BEJSqB2SqSvgykHP70GXsGK/x1GbxYEV+aV+Oc2Xye3ASLBd
gTyOZbAuZz9/K9u/GrGRMIwOhnNKsOuqYIRl7+D1KvmYy12S1P7RY4BWGo7Bd1pdpBgVoJ6gQNhP
oSzjmYpAKY2chf8dsD1yc135uDWG5As19wCMah7r8HPE7Lj/OlBZSICNYZELGyrB1z1mctp1S4hn
7FBd3N65IuEYnYvOgIsYjOu+f2cLnSBzCT/bf3ds1iMJVgc1MWc+Mm2xOd3Xik7b2x9+PEadB2Zq
4R+uU0YW9VKdHHSsjaofzVUWDnY+RP/CM8R6Y1FXphTIIYPCxikzA5m0M2EFN39D/TQPi3/g6vXy
8n5rAhfuNTgy5wLL78PEptK7RTeiuyXPHNA7doxWn6Mu6yNKAnTKubQobqPmqRoz6oWFhO1FDg6T
vpBu6aiE9yKp+rx3F5CiE0TajMDADOHfy5qQkM7kTPVnjiOsEZLFg/qhQRQ3sEmAXEhR09Zwjrfn
NOd0a8f590uVd2aCN1SzAOIVtZtn0fPekN+Pc/91sS0JV4HXeKD1IVxzmS/cXMrPeE4EsnG8589k
5hxyUpJ1d9Oo+F707X1mo8/It8qjtfQgvVX9Tv17YfyTpcmg4MxTHYQZdOkKgv88koFzYltOI1go
3URbW9XFYj0Y8UL0ckGcHfuls4fGazeFItKpZW17WTR3QomyM4Sxm5ADzinC7lTaLXkHPKQfIRbG
ZzQcrafaLwqyLWwFCs4wEQ3HkPzP8OqZgMM+eEL4Sj39AunboQE1jlSNdJh23K+SpMHYqwGddZ7O
+w7qzAj24MahBreLnUPodUU+6Q+PZq7PoGDSw3Au41z6bcA/DqfHY6t85Ti4ozvpmS4ynQwZ3ajP
UqAsuv5sas9CP9ggKRlPRetVVy207EISekhpC0PN4/Ek8D4ty5zTj/PWO62vHrwA01wAf23917qA
zEF9J10oQ1nbpMsxlvK5MZ9M5ISqMZopdG+dGtQfKq0HiNp3CAvNcyJ4FeqvRIyHz9NK1B5qe1gA
CcKC/Fy0/9QLhnQjnOgn36ciiIQTISm8pv1UPCUs+FYZMwfBpxfy/34+vgu0KWppQtc/mKEz1Bds
pLhKWjFikE+cNv/6cCQI1mENEoGiwpkFBDP9brPnAFU38fuIKRxVTa17+Ce5YzSh+IGJkwSlFead
mz974AorBWV/rFDzd1huLnpv3m5hgqkRTcD50U3+LeNdX7h6BfgahSs/nXGA1RCdrC55jk3HCY6P
MFgwGqcfqwanVvo8gt+6hafTsF2Zmbu1KbRtDybX4NAvHJA8X4kge+/YrxD+GwvGfmffHW80rf6h
1TMVoR7EgaXSyLb2Jj0r3QCVwgLWzFl6RzNOUR7+QePShkCf4fk4s+HnsehPGZdSB8P3YMr72F8S
zCpb2nawYZ1w1bToLt/x/RwTGW8eud2bHpws9ceRdKjYm+3ZNfVNeJLnyxx+kf/TveVeu2HgD7Dr
9s8ajsJRHxTXPlRO6n3EvMaLSACA28gSu2sA+yix6oXxX/rC4tTFaPLFuUzX3V2d9c7nsYsthLPw
I83E1ITBaUmOWH6yzSk1z1QqBnsh5fAMB3X5sICsrBOs9ULC4St/uxE0Bc4Cp8++Fb6ANIsjnRWy
dad/WrwXC+v4A/Vvn67MVEDvmeCjItAkknbaZYNK+FM1pZqLmKyWINb3ZRiRxGfEXX3np8jKZ20o
09SWN0Ujsrwc1NezUPr1NLKtT99GM4Wqp8YDqWHvvbfQ+CW6j1UvdgJ7RC8Ihkdd6T69TPMOCSVj
ERAAmk2yWtH/A5BU49puDITgpyTRm9ZInBBgsyGW8RutcSSHfMYMkZoN62JEwYiY8CPXvJs3Z+Ln
1G+XxCd302aOYYWH0SBc4u/Y86KPygD0Ex5TXtc06LAeHiM0MCLq9bmFNPEohFlAXLTFnu1CsFEQ
y3DOJPxfMrX61Uuao85W8P8iEUPN2PJ6waFV4kZxCMqPUP3X+Grr7rRwqtJu0x7rAsW7bek2MZJX
nNep7iRWaVUjxFS3xF0+cPGz+aOeKDIxGtFfw4PcUj00kHiGuvqX2RD/wX76eEA8tObDsg16vOuH
uo6jsOGorg0CzhbFyCHiJC0YgLveV5YPJWFuXpORzmRethkknpj48a4bg4x8u80V3LiyIM/16IGu
JvhGsixqmsbBdF2DJVf2ld7QvlZCuX2sB/v4blEq83FVhJ+UB0J2tkk3jn2w79mS8J3UeqCGRKp5
SxdsmBKMY/TDQD9OiFmZfcCQ+waI0NmdnHt+RCWND5/hET6Nv5incLK2BIIgHfSHNUND8s8BOHHU
gBgjdB0hMpI9LQuYsr5JfgNxRkW322HCZfxRkQoHdsSe2QyjBm/kM6XElNvF2yWOQd95X/07vC7S
DOhXD4BgRkbyPSaA0d6hVyG1GkIHXfVVHuY4MJhjjyjwZqVRzcQK+1LGwlmZCKDLfYHcJMwAS3dD
VGui9Qxgxj2lsBZ9Oc9DHDvS5fQnkU/4Rh3FcZWMlJ1TBKuk8x+l+jEYuFmWwqXKP+ArBW23jOs0
+phV72Saj2uEDcuWJ0Cpo3E54i8jnVGzf9BXRdL1uqKD+4ZQf3dl+VIihXWckNhy9gh7Yu7ghEbx
TASWbeIGvPpQp9YWK7/wmMG3MPMIqvGcj/10DWVLxhn33yZsUJptG5GpNxE9eHUn5M8+yHbvC9bJ
qwFbOj8eluv1AuBA2QKx/kzGNI4TwL7U6he+RowQlOGLlbl6ZwFF8FSUyZmlIfmsH60i9V4Pj7E5
R9JniPxn/FHgMOAUu+l8MY4EK1dYwXISFmnZ2dmx2l1sfaS/Bk6xJ+ZfKIu9UMHsN4qgGz3IRA49
20AX2S3BHcy6LsZUtXEhWM2R7MNV71oVCRc4q4e5lZKaZgmrNuM/v7BcuA43R9Zztmi3o1o58TDs
6vfT9wELF40/tqKWyO6bgE6LBRSPAmfRLzneXucO4KEsfBBv3hGR6/qdFXi5CFmr4PuVx0aXj4ah
l2CkTh4gQ4Jn+B4MAyQD3YMBTQbyr6YsBQqs2mGZ0MxOcADq7VOS0VDKmwLwWuzWobzYa4pQjLoP
X6zNL/ReVkM2hS2R3gfk9vYyDYHAjt961KizRI1MC8yQ0lRBaWEaLQPNf+7+9/uY+AgjrJ6Zg3U7
++FiZM+TqtB+8dodt8NB122qqKJQZjL0If13qdKgVN6nOJ7e3OdE6CozrCBZxtpH4DpGXF1HrQKG
zPL7iUwoqZbxpe/Tm1RMDtbFDGaVASAqE/MmMlg750v99QqsWWov6szcAOSfxB0Dg9kjKHNDN60O
xc812BO80i1XObF8tYXaFdEwskzk01H1JgGVRL0jQ3CQ5cKoxStQQ7GVHsKcNk0ccOqijQHXOCnR
QIEF/9r+ErRK1kRb7Rsd4sDyOht/U4RbtnBK3AjaxqFI+Sn9yaOf96ov6L5JS3DKv0q866ZtSEUY
DBizebD4NFqgJPMHapRHXz9itSozmkG7vMTlR5Sc1VPGj2HtPFOe/w3QLfYSWiFkMYf8+IJ883K3
Qpf/GP1lzC2eLTmO3kSsDig0q6zzKhfLdQAHd2M48bRzZLHHHswTShOtRljxsW+5hYNeJjAS8JgX
CSWSZQ+2Y5Yj4xxWZZ7P+v/LxyrIYXutOQuWKwhG/egdWcUfb1Tt0PhXKKeHzKLcWS2oP9SS68QH
7Rj+Yt8v+vJcXSvlBIJQgtflwfSV74hoE/JFe8CmXX3M3VLj5jsZCzmgdexaIm7l5BKDiMoMwz6y
MCD3P2pt6Iz3CQKQBqxHenkWCRz71l1U/KzlUnM5z6lhaZnD79lDDCgusNCTVTJTv5QMsEQYHvb1
yhRwp4jA3qq7K8qTQnUmVDIfDO7a2igRqX7P+POhQpHmcjP2zcdQww1Zfgb7JjqpsKyp0c+rJPrk
gy9I9bGv6380BvZAV6u9E/jYHjpN1BbC37gWM2p1qVWJCITb+wqTKqj1mEsdfBb5hJz/vOdu5j5l
cBBBduQaTdC2HqTHbug0QYNyci4NP7V/xVsXUj0ovTie88GBThFp+rwza/HpFkFIrNmX0h2WIK3q
/57DApcJamrk6BH4pDbI7o1qJpOn7lcNA+LvolEgejzqYkK4AzjL567RktYzcLnGlN3X6caExoZN
3vLyejmM307nYwIZhWJkqMJHVh8MspDehTlPcniu3MDg8B6OWWqmwq1lFcpChIE6dsvJdKDqL2xj
w0fhR5ScbtLCCovaDXHaV6uZw3fjFhgRCvOicfcsGan4qBblBvJx0HPRyOinup7mkSTdwm+aMjeg
nPoKfC4lPsnjjwi6uLH4MxKC3aGEcV0EFTOsFNqCTMUDQkEn/rVZTVU87QcL0E+TeXb7O8ytQ92e
TsoIIzOsPaSy2xmiqGpLoyoz74M2/csf+sDBJpqSamRzeutwzO59Ee9J76xDl0BzEguiJF/F1wGz
4YD+ovM77K2MEvFU+lenKpQKEny93UqBP0IJyH8uYBg+DcluwmxhlbsP/jX5QmIpzSHQtyb4J+fM
Bc0eLh2Kqu/uANtpkWZqsTIWBsMUYvmNHMqnzcTqrHXYQ/fNb6+gqf2qWXLlaPaFEYMqPva0Eg9S
DcdcCTQkBCv7A7xNVXlZ7x8EhYZ1WGlC6x7jtOoML2o9JkjhnJPlqzx+3NNR30DudRhEPQBFK991
Uebj64DktJC3aXh88/cOqRF0PYNTzEa5HAXqJcPfAqzV4KuVD52z+f4aNfbnHv9CA2LLHwJ8jwc9
4G6iva9+9KYs1e6tjBwZ8zsQ0LEPr0+Cky477mie6QBboDlDpkT36gUu2wU3uoe9u0tmbPMQXycZ
7SJGyIwTb93IqhBDV7TmJuerqT/6R4MiRx1t95nR4ExgDFDPYfXUvuG8kDhL3jAqgw5cgny7SFpv
elmYalmbmwTPCTz5Slx3adcn6bBrcI938f0JKEfa5ERF9fVrENCqnAO6r2cD5SSNyjfm8vzbeFri
JzstscpiPhVw5m5Ph27rABB/QiciNtrmWF7GWfF3CA411el5xQElKExqs6CUOFWZkYQY9Prwd/+g
F3H41DTEFTtid74F8h4ACYawGQn9M2o/Nngn4Hlq6y0vSwogPdFpy+tpVQtYiUyz1N1fwELv+qbX
0UqYYvj83UXN7J8yjlcH/R6Cb8/cyFOkRWckTrRFLB0exm+JFCf5xmatvU2xcRTaxIiD1K+/sh0e
Ck+Admu+LTrL5bO/yU/QCiUqIZmAtiJdRqox3yZwch0U68qPlCI4GkwlrUnSTNGp0kbSydzN/M9w
ThWYTq4HZOaHw9QVLqCzGVIpRJ4GGvKDP70EoXQjv3z2stukVc0gXuNdx1l1gIi/jiTZf77yub3V
m3YJE8jNgXBuJI727lVGi36jCW4cprDOHgfJUwWWSNdnA+qxI4PR9AhkgY/4UJzjv7hsLoL8/7Y/
k6bV1mJzqfRA3tHN3s6We7vrnmhJQHVBhj9nrC0pn+6/xZ1bE3QG4Rag/vUHb3othVV2jLZFwFK9
EHThUXHBSDhAeXYfqZCs4tmT2daoi1AKz4EVwWEWpnuuWqgf4sBQk/udFn9ZzTSBVsOpFJ9YvPDH
SAxxI5eTmvsWmjtCqZgVEGhQtA3Q2lrNk3VZ61joIrzLd/mlqh6KSH5TYebhklBhZUc/JblTax6h
tF5+pNYfEpxPreDrmwrZ5eAcvh4op1eNnOVmvELs0Kn8rCgwEm5jmCT6w4o3Fmor1qVD3mEbse3c
4IAeon9oXcnEkycN8Kjf26jYECRIYhbj8hKH7gICDnyBr7iBNCstZ33TUuHL9j4jcY+9Bscdbtzg
wHUqPdisC/ifPJITDEUXKgfSX7D3TUd6AJXN6xix8Yey0gFqds7wT0NgDnmcEmD1w44uafgcVq3R
xAabVYFr8PHpwyg8sXCNW8d0tZQdJVznQpgq0eYuur5RpJIIuH8pOWVq2FJSXJPBOz7obWY6IBf8
iUp4UFcdL3g7wV392RlxO2z7ELRR8DpASVeS66UfQgKRdEyf9ELz8HsD88SvosG+3/DjYa4ocx3u
kHSV+Hl9MQptNK4Y7Dpm3JLLNkKCpMRo7bQmY0Uu4QBz2nRXxVdgPDfZKtevgreDYHHNRt5ppq7b
jHwj/GAlNYcK0S0Sj7EjVRqab5pjxy/8yretJVurN38r8/CKiNoKCsIjTT9FEjFCZuGHG8/k/Qtk
rT79LDviXtR7BrKjPMssZ7BIS9hq+QXIS56Uqy23hW5mrVn68ROoHFrTtQNgbPMVQB/vIkxIxoX1
mu47Wa9t9QLZDuQFKQJkT3WsQ1ijfQ0otEKwfUONHMt4i4bgJIdH3G6oaixS2woNtNveDhGJaFAm
IrMgtv9nGl23+yycPE6ygpJbQbUz9E2Ql8FtqM31kI4qctJ7dBFUQ9SLBzlwni2PtUBuPd6ayXag
Q4Fj5Wv9/IAovB/bLZb3Qi77S1B2wJjoPZW3iNCSLgZ0ws3pa0ggna7/DhYSSNrLiv/XNkxkkjd8
AyJsvPBSOZNT7+21LGen7Fryeob8x+H+fmGyBaTV7hqMmUwglByMeOFXhgvaFWeyasFHqR91r/Qe
LjYsO0R1C8vbUNKe3d8WZS64S0X4RagUVo7Dv3TaUbfePUE0V+zBkFt/TfTw2T5GlHq5XRzw8GUB
IYbD3gRgg8jn0pYpfLmXH/piU/dXsl1pkHIVPnWWmAbLc6ZLfvLvbgFN16dvV9Mh4wfF3ivI3xPs
M4Kj+Qh/Qfq18meWHyinGWb5ZiiRQ+PqKQ9cecdXZOHTqNQ1RliDXLRgwog8Hp+apArsAmMqHTB3
RVcI+WB0DJEyOP4+CJIMnWK0bd/TohnXEyPI2ZxktgHKoX12XlbHGi1c6xdCSr9e3QCdWDRBDiMr
0iuIDxGbq15rFKcHj/cvs6g2ycTWF8ijPFFsaKnXzJ3uqzk2klMRF/vQoQR4nQ3JmeR75kXCy9pi
2F0VkIAaW19kMgDVuseyQGixAy0ZY/82z38Zc0qEOAO+BIS4cx1qp7OyTovliKcU16RNc45ogNbC
jhNqpdYENpU+THnmlw6Uthvfz1rCf9YB5FCFL7kbpVhpq7ITUqXENVdQTIjwe8r1lTscM/dd0edX
ROM8NDc1N/TbPA21IS0jyEyuu0kDyuCcIP8VVMhfQ5RQxifMr6fyYSD9mGFWaQA3ni/ps8Mmy/8V
Ec3DpIzBceGPd7gBPxi4kxEqNGznFDn0Z8w38hbAX6AaGjUHlcI9GGBa4qmAWQSanRWaIz1zuwPw
VJ+Ezo52E70uisG6s/+drmgfq0JimgTA57cseGBiwC0jzf294yTe0kT3QIOYJNd9uHZtY/7xPfbX
k0GCoFef7l1fjkboPfphbHpLBNiSzChblQMocPOwdeRZ9i4vFyILo9TtnEt6AqsBJhlZYlijaH3m
rqb1OQKzNYejF6dXW4DegPP8ikIezpdE6E458Tcz5YywKM2YdpdTc6lr6XcVW8dgM+KCWptJ+i2L
fFkiGF9MHJA0LWAgxTgvIf+tlWyYLZub53atmX3hGE+chX+TqkVsrdX/z2C+SLtWM9TC8i76L1QP
rpRx4R3OvWITm2TXzFecp0agtniO1ieUPep2+1I4lojexcoE2LiY0SQPCJhNPbVCzOeUHcG0ata4
a7A6IQFGaZGFH7av7hcsyPYwyPrKxWmjE3i3UzH0NJRyGaC660pPG5DJ4PqtopEN/8tDlySKEwyZ
xqaUBO8ghTERQtMNO8KEtlLum+lgIykEjiaEqZpoktKxaZSoVnGyNNcVMFAT7vZWLWerRQ7D64Ur
yrV8u09p8ULO70qMh9dV5eoYk/oDMb6YK7kNSSlS9xMERl/FF4pZvVzJa8dLDqmTmQHr6eYV8UWb
873A8dPAf5ZSHMXb3WOU0ZhZW/2He72UEnYJMR8rlsPp2SHPAwqgm+GeyPQkP/ElL9vbGn02MKP+
VADDpE77aRNSETAUlc2vtoNU420rGm1jDfEIdS3T1mxW4WVv1DZ0mClhWWcVLeOHlhBw9+GdyaBz
+vyU65VkmdriPmsGIIZhNgj71qCHqNOvr4BT+E6LPE9P0XqozoU0zg75uY9UkhzQfgjqkLgmLi5x
AmTw2LsdriFY6A8BaYp/8Slui1A3S3+mmZVVjR1CjIcRKs9IzNS29fvls2pQ7YxkE1zRKTGoeD29
8sWCvznGLf7ChnnsSI+blaHtT3sc2uhHoIVApEU3VrT70niQPJNjv3Y4xZmwdtuDR9fHeXJM72ib
L8DPueFN7I8aeu3FC7n6i2HLtwlrl9MUBxR19uWTxk9ktkdncXuBzb38CqDsrKg4pqzq6BFUqdxQ
Vtp0T4DzxrPU3TAcQC8auGe/8s4eqThZeUpfHrV9A7ruyEtaE6Hity0v+u7VtvmgoSrZeyMnn9V3
XK46M25AdviqHge4SCJDoMawGStjr/ovS7eBEXpSr3480vxFTDBQpKMKd9Ze3AQVa0YgTWdtQ/nh
LrFxKF/W3I18WB/VWMs31HFAhmoZ6CkiyU+Zsf7Ehb9qIFAAZLpL4A2zhatIRO4jZgYuLxCGhZsJ
mmrh6XIB+IpwiLjTLbZ0bF0T3btU+oc5ic9ZtsG/q2rplUI+3GQa42pG1W0sPRgsVBj8ea8Oa05I
q7oXt8bnBebkrFLcYHpS/WzRXuKrimhcbmaDFXWfThnKkslPLsLGBH7cdlwyz5Wf21zEOvCuc8uZ
kILQlWv89eT29PMwSp5KsQOHRAtjtsPr+n3emofQ5VU1YKU48wtoJ+/niTZrA9Lp2r6aU7BQS+a/
zsYYydzVXxYoV3PnvEESG2wUm/WAIcKbtqV5dWwcmjzM6JeRODzQXNG8aDOXZDJmPpKF1Gp3Knfe
xQEML0kG/xUMSberRK/f9SvqZESPU2LROcEdupC+nma53IdWSpO70MG4zkJ3RpJpphTg3Nk6Z5OX
Q69oOaJxxSjjREp5NukTdmw7GKyeVhifmVxWbAJ6ics8kL7dqfxlHymrFXdoZ7qJ6avM8Pt+XiZh
VCQpjNlNqIXebRoqLdQgsP4tUrxCYGZgHdIhvpKeIbIJQtzyRFYcgNiyFVRI0liNuR23MYJoBeDX
aafBER4D48tILzs+7gXYZgNn1SIL8SK9BMxPozqrFYLWRxz6l3hx9mHLYgPOz2eRQ37JBfbm3F+R
T+AflnRAtK9D6zVx+YeUnxosC4heTPjaY9TVieIa2wCkk6NpA9u1xPtpX8jVHDuqNI3F0aTFAWNk
zxR3TqhE471SrqI0Quv8+tqfLM6mDTiaD47YjQFr2cWheaNnwKlqMlf49DF0mmrrfRceqUPNSO+s
KV0H/tM0UEUXOwKNUo5oGUJeiJhN/OnP1eTdS90Fu3K9MiZC7k+p6vhjSAm4IfBtfnrz3mv/Y9e7
kEHaxBVQaJH99jM630Aenu+HHJx45OwHGscMTvOLdMsXVh357c9cut/QZXtR303GPEpxHEBJH3ML
iZfGYRewLoM92ynWLEHlY3/Ie+DvGnpdIebkckuJGZSjzPtnVLnhZqx8niMP/uJDdSUoqh1uLfud
dlyzn7svO7EMBvhaXTykCdFyownH0HWzPrORcDImFOabV/9XSUfqEy/zoRSN+VednmMVl2WQl4TD
JR8uGCINuzaxuljUZe4LWV8ABB0i6TI9SKrRuuTnqyCVRPeCIkJE6oB2LZEw8+g1nt584P8fvUUQ
O5HCF23aQok2P1a1xOD8Wqvt+esUikBK5MHc/ujMBiY9zcKrfXJerhWufql15vSQ5LF0uht1X5kb
tSCTg5CWECNpziI5yLF92lsMLWzmva3aflqD7fUeIQak4uUT5CYVjeDpk1txe10cKQExlUH54KIl
YjNIAujqqcAAq5oDpvFBoIk77/S/UdWOlocnMdSLJukuVSJO/tRu7aOLb8xk5Q5J2Pu60+sZZrL2
bfQ0fWuDmLZuv/I2gDhfTVGbbJfiknRM7aZxz+yLj5TxG+5cbQb7OZO1IAROjICwpYffLpy15+iy
jfqxU8pybRnBsNudVTjGoaHYtg80PYLshFaC4jiGyY/ItDlF5yGOzLLuC+rRYugtuyX59XhGqSYI
ZrwH+7H2GMtoFpFkzGk8sRcZLQT7+YltSWp8QK/FJwkBIxkqxptaHZlp8jUYkQTKFYp5OV8UAFUn
iTPt1opAffjRkIwa7onFiVrmnDjcKtkSxXnR9LxLF+LOJiCXOoqzt2aybO3anEOg+bKnyuoEGLUC
wNY6KIZncuYgnWrsrkICYem+KDOubld5sbGDkL9InrRXVNf3SWEgjhqyTkMxoe8jzJmoA2TWDrIZ
F/7x8dyKgn53hGhmaraJF5xx/rlm5+Rw+LUls50+otM80luPcitBlTVkD/EOaBm8uWDpQWBESHHl
LCcG5Ye38HQ6Mw0Pw2piauJjDocIO9TBHZ9H5TqBwLjwLXi64ti5fFLHHEsA+Oi2Xqimedya2cEc
s2Ocd9bsND+Eo9mv3h9IIe1otUu5meVpahWY/5xY2EX5MH58lxa7gl1+rx4Tq8cDIEAb4yt33kyL
+wzWnQWsRAicwcsZSTHOR0dC548WaWo9hShhy7ve0Tiz2Y6j54eqhS4x46Y7mAZbtcrOs05PDGfC
7ZPUAHj62fKxbFWVFdCRHBg2XJ+sjgPuZgZX2Q53QYbmR36LL3iw1qlbajaheLKk+tKrkzIPlAVI
bSuDc98yKQz+5o6XSsuihjzqALafbs3tYRA6SRiHYMXbhLoTLVilZneYZRrIEw+bx86ojN6FJdQ3
G9FMR3OnHVbYPjPBKnhShkJfNrGvBK4U8KgQMA+T8dB0XdFRDgOuegO26+Wh/bxX5j0p7ZUzWjqJ
hI3v7HV/WShkQO9mBfW1XuCRq/x4hP9DgW7hzzqcw17+nnl4sz6MdKh4DFhjfjW12wnVOzCOYLcz
7gBSUcewa+Ebj9IzCGro8YGeqeS3A7bZpjrUX6hwrP6bLEb/qQZ0U2yH4JmQsId/vHdk58dZbuJ8
llaPx064ixRK4B+qJO2QH6Fvci3aDuj3Ac4Y66yVCMF+zYqdwrO83wDkrvM7fWgg/EtjmZ6TH3pw
7Nvd8FDuyV5cyEYKXAgo9rhQZJNyUoLApZDK6Wvz71Ryamq1xjOVSHT5wi202Is2utLHs8NRtfMU
fXTmgBpRI3NxHijezcliWp6CJeOie9H1CIiAVp2+SQkcmWIQzkNmAG0Ty+XnyZuWO0yVuPOgkOca
dxsAk7f3BCnYMxlf7fuN1m1SkrcIV/v7SQZAoim7b7NrssReyhzCoViLUGry05B2AeGTx9jCAfro
dzsUooeNfPqA2cubs6MCYjNgZkjcZxmrHecUTHT6wmbiIWY9HqLtzw6re/57hnyvGh6XBlPiDw9R
RKidsinvcJSf60Jk5MS/QntwmG1oj9h/wkiK9OyAOViZHjg/juqTC8xmQa5eeYAUYe5OqBEcDaMU
vhwWnr+9xBmAUrz+q77UiL5DGP0f+ZcvCQzCapBu3f7D88jyMMJvE3P8lzvY5LLGE2UCxdHdsRGk
hvf7mpHyFqdy9uApr9zP4tAUBdqd0nO4pC4OUpnVlX6VNjBMIr/iTmHCWVpvMGDrFUjLf4uUF6O+
UGaRAsMYXK4OvnKpEW2XZa9MUGLNDaWxdtsgc5U54DcZ5EmbNz8+CwqIz7R5YeWyLm7kXDSMQOOi
pyX14pokGwCt3Jea4FLJNtiFhpV0xeVWFWIZDgDOodT0wEF4A3FPFoJvJMRau+SAqpNVken8aqTL
lc4p6Ouggc9WECcY0OqQavBmnSu4qs0bAmReO4SIewnbKkyazPZIBD4eBpqnMCOycx5aj0WjhnMP
aMAT2isHy/Juj2nfqgBkAEZODAFDx422GqfrqBIxGlzjkdLjg+Qf20nWEDnLiQLKZMU8MC4kt9WV
nlmti4jo7UFfFTQr4EuKmBER+Lo1FUK3Ns8PNkF919sBa2Dfq34YTuSglsF4PBArPAIHjyb7O4YG
Bt7UhC+haOBi3bV19u8wIl+ePdVGZY1eoyFmBWb77sdJ/5TYWKRc3mKg7qfrL0LZjcLPMSZo3Q77
CnmO7KKsdTq7O00LZwM1+q+xUyDnqw7IBcVZkfDowpD2eXdh+XTTkmrLzVfZLSVPKUidMeQ0ZxtA
yQsT0sk5wc3V2ke+/zprWz6yGERF37ASPF0a9LGIF1tdzDjTqu9IrGtK2/10/wK8hgpBM62Oagyt
YyXS7wOl/d4CNO2zLieU3ZLaTUoRK7UndLHplR7LW7kW/pH+iGmhaMagcbJ4wurzClSet9uh+UNU
N7/u3wKySZylJnqO5vFuYaG9pz2lFW2/58Dzu7a8CoR8YbA6d8LA3s7jcP+meGBw4yUisrlWipXk
K2hhsbh7wkZHWTga8+yeDtiEkDXMoRkuSkKD8SGuAuZt0uNX37Ek07HHVj6MPTm7gsoF/nARLfNE
rhDVDmosSbuoxp7WtWgOxN8c5V0pXRTFYPP4riTVdtrNxbeLRXvx16QO6fQxV5Q44iPSA+VcPL1h
7dNOmmrIOcRu2bPJvEigPGkbPtaK+oZO6+97L16BLESU665PjFt0m/+LuWy0FxWIRXVIPPt1JLhb
Ymj89ESEjUkwk2t60Joq6+EKbP0wFci7lk7MsXZ4pv1DTkG4KsbE5sKgLuNTLPirIZ8XGpPjAqqZ
S7FGf4l+GTIBFl1Vpe0I1lNYwHb4JCGiz6W8hkfX27GvHxMAUKn4uEOruKPDLjXKvPWBiEsfch7v
+uP6Q6OAcmfiVOisIebqfa7Ou26rlUnf71thma3jcJQI2j4kB+2eMRbtC41w/VbEZWtCc0mh/lcG
fTMNINmw4gpLwFuLPoh4Yari1yCki2AXYBocIG/er8yMxMkBS0LmZh8vdVSL4X4vlI410DLAcDu0
WiOnBgFcnSSElOFX3yssKsmcUspJAPTKY8HYFQP9xLTg/Nrs3na8ygeMqXWZ+gSlHA8JDxoVtFRN
U2zjW0Ca/zPIfwKQ7v50Twcv2Lz2EnvJqW7VYILYH+qTc+xLXajOkH57q2cnyfDDEARp2/A84LIr
80yvGy8PCmRoepLrROsHwA0ILqg7kbH8KaXEYIzaFB9E8hQYIIhj13dQRabiY9pZdQlQIZgDHNwC
g5PsMN1IXU3QDbr2LO3jcj6FIiz8lQpLyr7xEMnEbQnfrk6ZGCmg9er5hosNPEjTKeVvPDeU1d5i
AWgsZe/qfNzdrJDCch7crIiZnBkmOVKWRkFiqvOOwBrCN9W7AcBWnP/86usxzjUgIG2+gL9Qm72C
9+zMVzZcuTswDVX3hgR+Tsw8HfftewrDsPZsUezRiN35pvpAJktzNWaIB5J65y8WPd2kO5S/ddg+
SbP4Rz3sFGHmuU8IiYlmXT6+dEO3t9XkDLVmz/vUpcMlpWmc8uO8eHRgaug0CTZdpszOu6XFTUlb
kTsGDSdb1ZPc4tHZOfTixkMxown99mjE9Kfug/XyHxLvZ6wei4NzNUbFshVRQA8XGJZNWyLVva37
F9wiXit+FJPW4lKEj4ZuR3nVuR86RGTJvROBqPILhcUyMfmKg0cC7J+F1I88DYsC406zO4cPY7Gl
CjHgInrOXxUbr73p8sJkQRRnaVt7GVuOJrPd0H2ZlMwUYfsJJe3Kdi0n8AKtNmYleRHV8JrSiuoN
9/9XLaHdC6eemjVZceKt/AJ7780eLhwl5RajPs9oaRSo0+dNJbp0Xd+57rGM3gUQpJ+xNZ285Uux
cid8HmSfvxUKtp1rx8DNDEZlQrVXIZBj8x7A7oaLixGS9tWztMh/LswXbWQfwZA4w7WTjM7KbsTq
Sf9776CnwU3eD2RslafHnFrdW+lE6miO4TOtdlchnKN2ekkfxtLL/N//iX6YoCUAXlLT5rGWGyty
SA7H/XtF31HRvuljPQE6T4Nk1u+Bamqmk1XGlAslioHQ94n+QRlhS4pc/f9SAxmAx6ttdHGhd2PH
kQeYEj9Pb92R5BMqOOtkvXCXsY+nGGa71Ss05kkgIulzBKU3/nmdJEZIq7DaCiF/2qfTjGCtchic
uFIYZaaPhk53OnwcPjv9rK4Ghk9SXFZwo/UeGZSVEdpJRnlZ4c67N/pSAiUIoDBjW8wGs97gbMbA
EreRQdtefbFf683upw/hju5aMT5He1uBv/GxDVnVE1ExPQqKADkd/ZqWZC8gbCWId92daS65ed+J
Rksf4hTv54Y7upWWz4QBM7PaaRR1IQGkGL50NruxF/fCbweaS4B7dinEp5b5KFBr6NYVOZlx8Fxj
CxSQwCkplw4+NWyJdTBK8uVSQbaxURyiBFv91qbv8qt+w1H/ctkDnmtAYmUK3HErhc/81n2OvIbw
W8Zz+ZxMeU0wAF3vUj6Hqj0FCvawT2xFaTGKnZ0djF49QyijP540wn7IaHtl8SUuhksOTyiTpib4
ZEVBi/3y4tvFzT4fxBmtzJ2olo41b2ygc+A7GTQFXiZMx6qipmOr+pamLE9AYgPyv5n7p+1yS0hi
rYS6SU6U9/Gb4cdFZgDuVTQq9DWE+bqL/8P8q8b5SPAcHuOIYOD4qgkmV19n1o/H+yOlPeEyVsEV
ODx9APqNKuUCUF24pA7wnbr0NOb67lDHduBem729S/Wpy+1P3HloqPZydJzJQ+RtajSWuXG2OAmy
shMhr/AXllReWCLON5Uxa6tLhWIZELznNS9NsKFE9PMm+NXusxxrhTdo/jCYc2gjAQjsdN3eGXON
Wi3RbW7WJsYTyKQBxHRzNf33BIGv/p8Aueoqsym8MF3FjfWfx808Y81pvyFpjjAhVe9d52RKkXeK
ahRzTwdY0WwY8Tf7pty7yTya67DiO6dF4UJCmFHxBtL7ZuObhaqmRnmJvwru/EMEaHbYnr3RPjaI
PNOu2Voo9t43MZJeFfLQOPo2aDpSo4bdX6jebBqHXkeC6UzB08rEIFcR5YCwBrLwaOMUnE1/r5ys
e02WTulfIvUJ2WkdPevK0tRhFkY8zzzkpfmcAZ+2EpW5hea7+Zn5zDBvVes6zwNuYrBv81b6kHw9
eMXXxXT1kHVbQ/CO/Up0uE6V6z/qdJmYuwJJaI8/h7WyG+fvhhPeoQYcQK4Vrzc6tWxjOzhIEFE9
SQIkNaLUQSVKULE36yKaUF2l4ZFw2EJhwo6dpqXVmNgo8RG9K4LXwgFTRfVopBk2ApeabhNbzbvI
FS8QKS0L5un/YPa1PWZRIf4cmuR2xoSqO98Zmrvh0hLittrat0n4Ak91Wi44laW7ULedTwzaTejx
iq1w7zRw/HAYZ49VV6AngHk5APooSqOOiQS/9xjAkK3lGCDE4IUCgwwHr0GYr/VruIJQ0gFzImR5
U6O+AnO2mP4UvehM7xe5ttOURr4DNwA+6lxm6VB+xwK0AAY5Vnc4Ge7fuQ4QYvU3gPUFFe7lpnho
+VYRCZfmDztDZIW9MTSVWY8SLcOUSorKAYvptwpJ2D/V87j/vwihNEVqYTYQTuETg26x76sVkVbA
VOQWuT/+KYMs8htqb0Uwy+LkMJMqrKxz/BELpqk2VcCurjr9qcEVlQQPKs7AThObfQ0G05HgZifh
mOZMAecnpQhg4pDHshpmsOlGwz4QTFvG4BOFUL91QiX2So0kdpMT8TRSxl81I7fARFRdI1SP0fHJ
fgiUKwQ+Y2WFXgVIOx44bYAE1J9F3bKW0+GqVlwdR0QdI/C9WV3TLRYlo5WSmOPHu217qTFxbeyw
+p2IVwglf4oBbMBfQ2UGIKAHjrnJpafCxrytYqjbFepliSabPFB1nUydWfzlPyUf25BJjbBeGlHq
iT+wGUVqZOUn79jTh7eMTFrZ047EZ59dEtHiu8dzo8X1E3LDhOzaedQB5D89M99/f5BbaH+RAixf
TzDo6/hyihRRHPIiruGhcTCrQEkx9DACFW/ZvJxeOHoEi2ZNO2D8h1S7824WF2xCqO17nODAiLws
Lcl5M4EjQwo8Sr5a9vQOVEplfMMJ7jd6f4rQBDrYPC2nLwr+vpd+LHEL8n9C1HMBISiIkQXO2tbF
OVdSGRpxYc+i7ovQJdjJCjgm1pbuKnlrWl0b/vZAo+vTHSUguINqqaKSrdF23sdZQJ5KLn7kCGKf
zmhNYr3+NdyrPskomLg3P7ei9JsHzXvHPu/qaBoO+Bju50nD/a7K86pQG0UlEZlvq4HRG7ugnBYE
VfX8+4EchjvZnJTpZq0m71GpstI0vdwd8LXy6wy3jSIvC/xLj2uQu2jQdfViSi80BUbU0f8q5Kmg
Q3jy/j4Eq4pMgIaaRtAOM4G4URXoACh9SBs+ZONdMOmSWJUKETtIug/P/d6o+Ewmr+uiR04AmP+b
khAZIrObn/yMA5epSVnCr9yzi3glDIG5Er2I8HVOlWK/21t1m0BnH9xUYcENFoztA8HrzP710VMF
Rb4JeNjVCfN0SHGJn9cyxQYs9r2IGBR71Rl9if+DiA/XupFVRLY3Ik2TkxrCpN8dhFZ5kC4cQm+E
ZbDLuhtjbcgLbAlOmqtkOOZTRsroglRvu5mDfEap24JgbH6VHkuQlka96T8oB9orictdYbROURiA
rwVGzOS6wEeeeoTbu+sIufSCeX8deqaCuhNA+l6r6OCjHWZc2aiE15/ANF73pRPRqdMjJz++QOvC
PnB688ssKEpjMoa6/zlTwPC0kJf2roKT33SgiekQXB/YDxkB+dBeP+PzWRPHkk7OsM1rRdfcFXAl
H1WJZb7GhmCleB1fJpcX5BW+qCtxvB4Pq+lkSJ+b5/XUJbZgZng90lbZFdetBLz/Aqvoc+uuvSre
wfu4Mhr/Hsh1zMIn6ulGMIJjF2XFDKrdK1auOwgHER+TQULnv/BTbz0JSu0WWhf6bYUc65vOcAtW
Pb/hDlfW69DDHDFZoPADsHtIawQfGUjhsDPC+D3GzcClSlmJfP8zlMDCUIjlysq8yFMAONVZj4Bn
iBj3rdxydQJ3x2+6fkq5BNv8bkjfU+GQQo4mpgYOXk1PYo2WRP2sO/WF1K78RRP9TJ5BBVbphfQ9
bmxDJVckKMs2FfPfsYKOz32u141lgCy2/Cpv2czcUlVHay/ivADQsxs8m1cxuxaV83Z4+AU7ruEh
G6KKnSQG9MkgrW5b4/+7Te7FECUDJdG0wtIc+EGRnXsGx2Ri8saJIPOs8U1Ijq0vTOO73UrIAd5U
5k7nT+iCtCjEUt9B5bAdJkngbGWs8Ummo7HLQVYSbEkZj6fTrlVmZVyfY1E4KwXH/dg9RTDxG7Bj
4XiEIURd0/JG/33waTNc4E6biO6QwHVuSeuevlaWBT21gyeUfxKvZ6BNb/yiIfGlOOlENDJcXVYE
v8UgCcrOjl6oBgFcBUujgAroV078gkCpQCghfz/Bv9uRVosIRAL4FnhfPkRtkL1HvCP6eMdS1jbH
RF8pxJGjOFq6xZ1WR/OsfOw0qVu1tLTOeSRSP2AsxI/RGxjjVKYmnXaglSSJ5BIeJV1UW5Tpoyg5
jmLPhjmG333SaXWpaK1iXdD2xCN7V2cyv29FWW7bvFUiKZTZKVk0H+THhkoaTAsCMhzW5gpKBsp8
VvtTMrSzxlBxcOnoUAlEpLsHgThtMhRXHYpekuPEwQoDEJhySz+g5QIoLBaFCGgAU5gVgO38SyH4
umZN/gLsEBvSAKIuoklCR22SiRHOpbcQf3wIjeON/jh9DlJYkF+xDqOQqE4hCYiEJmYSwPT57JZx
iiIhckaxvU9py5wFvvwB5wf9rIV89Qb39aWA8mYIzR8qHX/4/UH1NQFvkH9Y/plFZyLRlyXHc5Re
Xxr6hSkv7lZBRfZvtgHukyNEKnEuXoVGSSOK/OCoj+g0TMjleq4UC7ge9+Z/UGAq7WNlTr/8wxOC
P/6QQanjlukETgh78rK/a6x3mNEtKj1wAJgKzXg3fbaCvCyMG4WG0pA8Jyb7szdStPnc9X2/lobU
rao0V7f74dYiVBOFysxieyKoVHUOxhef+9avNeaLQoEWjKLg0s11sgcQdF+yD4EIiYTWTXBZZUy0
A4KqvsgAqz4D+vb1FZHdfzzCasKOkB8A3PE72BvSnkEvh3jVthFU1XsxC1iZgMCHn85jduHk7J69
xFCUmkV3HYtYas7a3MiV8718avGr3l4bmPixe9RUCW0hIhXsFaKVP66k+2zIdTk1UsccdGUsTaUM
zmFwFk/fkJ5IYDciciUIg4fy+5NXT8kBfqQ7xmxAit9sDGpY1Ka2mhFdh0btZj++9v6wjzRNQRqC
Zj1do9kaG0fSD9S3Y/id8BhBbx41/DAb+O991+wgZZjbxhk+1l/v2RwUTKJRWrI2YeZqnFlaIYPf
kntLjgjvzkvzS6CPeS13x5WKds4PbIFKpbYxpole0XzVeDPiRlIT5jrz4rP8z1RzabqwBjaxXDI8
6i9oIXd85oeYrxf5QdXnKXpt6uLUFUifGFs1ai2g9l+3plztYay1Pp6cokanQzryuClU0G8pFOxF
YVTyGt+myYznCQHGGdT2LhdZLNA8MxNeNnNBuJENnJOGz3I8hmEhMnt6cxoGI9UAYWTOEZIuGilg
U/WSKK8ajh1Si6NWky20UlY3G0jNLL61R4bCdrJ9kQEAX9hoXrYKYKj0d8vbeDeZ25+yiSNGBVdl
GGBl2RpoNhqCQjO3swGbhIRBynOGXCqx2qVWLBQ5Rl6TfMBptux7QM558PI3lM28DJQd35jTdSo5
YyGD6JnwkNqhuWT/q5Lq4k35uWpJXbtE3rAzf0nWJugjPHc5Hjwrmhj7SkAP74hqCodHByAK+CAd
lxMdrMYVsH8oBGwOxN81MiSTD3F5/Kg7HT2fpXQwipcKPK9FiJm6jjExyFzENlo4XPlQozhRc9nQ
3ETJDnIj7w+jaHRkWw/U1n3M/uo45yKwXIskrk8uqypsWlzSO1Yho2UvSgAHICAHoamGmDb/DXdq
cRYPM7zdRQOoxNjLPm8BMPbhW42HaUAUt+G/3Ak0AsnCi1z41dXfzBXGyfUN71ZYBPFzVtjFI1ql
8N14G8Myx1wHzeE/y5SYQ50CbA4V6irEC4CX4KgJ2P05AnGgP5FuP7RuyBwHZpbF2gcHfDSaeevP
CrSIACBrHbCA9fpK7iilVZvXhQOHnqsw84y3Uin3lLPR2ev6XDxJCTM1s7RAOhM39E6TvSl93WYe
PX8tY96T6wr97r9nslw5re5D8PO28cbHyl/b256fkj+Mx4tZ3y/gI5kgMFdQHYoshPeWPA+H8tz+
a2+rwbonCrt32za1Ks9w1ts/IO2bhptmSGcy+WzEAIgktI/YWPzBlE3ACSCszyb2rNry5L/pIbJq
O27SA8//4vYITvgCV7q9g8KsHDfcZXhQfX4KQWcI00bqUu2VskcHfQWO4qmusTECzYcTw0k5yzGv
JW1O1aQ3NMJIxyMY88VBcdNvynhahF+HVakS6agFpElMqcA3FrA5Q48m+BnbNJXh2QOPjj45YGt+
9Vj4mNP5Tbjhv0jf6wYC44mwuYPo6jVb0jN2/ktzNHmKxP23PuH2cb21yxVpZtaDembi8WacifbN
CgVQ9ZxBY68VBN6HtidGO0mMYmNfTtYP9u/W1CRa0WFH/UcQVAyPAhdjpm2M6zoqWdcg4O05Xkts
DsKzhHaF14dia4tsnkKwst/4zVyVkMKpERwPlAOqcfMnDNMg4oZ2Fcx6sy0Ylki2+eHIwThW3j1k
7jraTAaKTqA07mErqL5grjNcX/Iy7Tr9Cu6qglgquDdxrP0YohUkdXBhtGk9OZ3kLKtJDHNr4ey6
SIOyPeCd/RIg914OtYO+4Mdr1VIIbrUfaqKyXjzxlTrSy4puSGIxPJxMQs7k+3+KaQ9ennTv3cNE
b5q7O4OJfTAFwo96HqeuLlx76Q78y66v1U3l+DOHwo53jWHDBqpW3QVvliPUD4Jk/rZJ9kE9SzlC
w6zs/wotO4N7c2s862O3lj5Kz6Vzdwfke+G/IUYBhQwecau4NVEinMwu0YVSCMagl8XWqSlxOuVE
bGYv8Fc793txmGJK2vOwqNHb+AyQsSCpf9qLGMQlrY/OqHHxgtC+FnNCFjFFBLaAeZ6APN9/+MUY
MtOO4csRn63vEvvXHKxYF5Fo4XmsySQlxnm1B+go0zfMp8Z4ygG7tRqYYYHa2ne3x17snaMEaBuo
k5M+sjgfXaY4TlUoYm8PeEMBEjNEV8taZGSqVeOO/9Dn0fS6FR4aYEJdUuE30g0OvNBvYQZhVYu9
3gkTcZ1MsecSCa3S0gs4FAxpTgjy9TokMOMbeFNF6Effyi765DuEyQi0nvWCGE41Lrn/dXZVr360
3dFyEPdhXQ/FBZ+LB3EKw59YKyZs368PbVw9thNrCK8siPXRxRe5kQmvJ8zB6WfyJ3UvQC7QjENZ
nkA/QxO5rKAliCmTFqiXqPcQs/Onj+VAiQfCg3DMdaMCoO0ZDDvpirl681UmpLM+MNjAHYUzIIOg
TbV/lHsv9tkxG6Q1bmjg5BqO3JqFBLZLoukuhfPCmCM/nAJyYxad09fTEHGw0rvR2ZFNhxD0BcqL
EpVCMg00ucNutpOofPJYsifxqoiyFI5ibeME07zi2Hkh7XopenfIm2PwVlRX0JpgcwgTV19DjKtm
DIsaeOQrpKG6QW9SZDF5dEIr1RYaRi4qUWb1cg4I4c7NbmgSPki0MJoI1EPXxw9xSEr6HArN8Kik
ybhYIuJL1DyicNUzThBLPW2O/RQnMULD/ynKLw6e3FPImlSPi+oWN/kms9i4EvdKrfDJipHi/BZS
4cza6kV0qpaEpFna1Z44Q0VII1BSZQgRLNKHH12ydNdBpkEvU+Up5qbXxbNGkWFJ6CGwaInp+XTV
JDOzBSzMdsWA0VnqmZVbgggxoWrRSm0/YBxLpektmU30FTGQy3XQ4QlN9ZM5qm6/VO835UVw+VPQ
8K1K2AXN8B78FCkbyMegu2lmMzsyD5hluot1kG79q26dh5rSq5qgLnyxtaU7OeFuga2ymUJR93uE
+W6AWVBNNIBm3UZHvwbPjgy9Oa6JD9L6/rHYbAtCHNCTcBets/rPsescSce0rK4dT+fkvdoeZ7TS
NokdykcKxO0iVAeaEnQFnAlUaARo+GiT2dv3tNYcsvd7ES8cUgvrgbuTWQKXQLSn7LhnnX0tUlCR
aPgMh40oCNguV9geOmD7bwFkhZ7k6C8yj5Rzx5Ufqdx1guUbmzGM/XrYVc/7J05SH+RF/swHKtaW
VKqSpGPyH6Qy7HZzb5yWMoFoxS/wYl7Z//YvHQapWyLRgSc1Pery9r+2qJ4lOXLxpAU6FCMjRdUc
8AhPAVuv+5psZyxMKaP1Jb3skJlOZmCPPoHfcvJmwMWwCPcmNuF8yLSOuNpfLo9Ivw05TkKk8OyX
NtsfoBL1uUJ1K9UK5JN8oe4qWV8JJVerP7YvzFpUw9lWqnPPAZFIXtOS8/0fiqc/yPxL5zh3nVrv
17o+zseBpoQJ9LyGWg+wIhtFn/wroJFf6e9wgKcAKEOgCwuTlxfjkyoOPq8yHBINbu9Wmy7qZWzP
lVTRw+jIGjCSYwhx6EoGAWJkfpLYmuhUTTLxRcbmgx0r58BdTTtl/Am/9yfkqYxXwiRsvretEI2B
0jfIvCw4FChjfUEnevRaWQ1j/C1YEJafuGiz5NBfbmgES2MxqrxZyS3fMS0rMP5mGVAoZAd2Hpy6
Qj2OFgJZDZKa/HfqRIVu2mxFGgqSa7odlGp4jJTl3fOVLIkSgFnd7lxbBaXaT8ikBzYpXbOby0JX
S34hFB82wXi3SQrh/AsA2vhPwHRJLszuFfW0N8wOMI/ESt/8Gb7gw/mXSC5YYS2wbvA6rYzp8ie8
yEV27Fan9digZI7DQyFW2LN7XHTV4Xv6Av2E1ADAatOa3FQLMjJGmVZ7NrROtGUS2fQXzchF9Rl2
ZFStvLqkwQmvlChhV+EVI4eo+rll+UtsITt51dzujmp26L7DaZFSXVeXS0hBpnb4+uJdChNYJFBk
2miDAaOLoEuciTa6b7U6tzcs+obh18zQJx6PbBoB+FMcQ3KwWv1wt3wDsC+pO4bXDGXkwRiuoHhW
P/mT65UK1KtpTdAUkCs9vtipMvmF/JfHloL9cW1o7BFn7cw94/IZgGXwVQEtnpqu2Q+GAVKeu9SQ
Pex7SRbmkFsu1KelzdqF8JkVQ7kGoELeEnG9KSJIN2Fu4LPrmp0VUzHi1gD2ncvWJqDsRZbzDKlr
no1vGVrBxsNM8/U79K/XN/Natp47KHdfJLtNajsiI2goVym3p/D9uSrcshR4nxOeVEtHtH37xXpu
ClNp7MjdWxBzCPlF8ke9hOKtX2fCPRXGEvdOsRM4cT/YN2rgyLHuAJqE7EhzMZtGu4RRrmxurq4h
TTtCA7lOXZmv0drXW7gIsTsWTXK+U8TNyqceXsuxlRCOLwf+/ggRCGkBbQpGudI8Sh4muqL4j1zD
8Qp2JUlAM+ZrxpTpf9VPKaNpdN8oL4a72RUu08Lmo45z7eQEpLaqBWoXx+F4V0TBgZ1EaDrZI2OE
kCpEb6sIWjcdydxAXOo9XzRzIhYaTJaMwW/YPK8ookoH4WACfjn7GpEU7CY5GfA/1PEtl0N7Gshs
YL5yldyCB3GG6HkmG6OD1xdpGsURaxls1FTU+x29dizf2XG/tn7+xyoZ0wUdyH2r6wwM/Gu5nTSZ
fln+DWQZm6AZKhwn0VmyhZKGENH3/197EfXnTz5n285zIjcrDVoOpN6m2k860wLCwuRN82HwLwHX
FMZxLE8wz4MGWmnHuvN2qDFHc0SsAOaEs7fbOgYd1FemrReMHDQvJUPuomtxT39wE2FL+Cift3+T
p0PoQNvYRlG73RQ5+l2K7Vl8963cL83aJNKgYNI4Gk64fcAAFDLJlvd6huQHf4sOWFeX6al2In/5
OjFqq0cbbTN8ohaaT/HqtgX+z6ckCF4mCgqPWqavRT8Y6pNryNcvWdiBF0Kj32avyAgljU2OIhZ1
stxKl75KFgLskYMKjV5tWSoWkWw4GzIG3OP4MkiWWP76dKXr6cfLqSibIws40XBYnYxvJM51DCsj
wOlbuYTjf+85FhGIn13h0rXxVP55V2nglTaWGlBlNTtZt1pBFVnhXQddvjdWLDjCnmMc4901AdEs
sbESiFyxibdb5dPqvRBZTtydL+PHq74KsL3hp8x8eUx+tL4260HjYK6uxTDDiVm3P7Ab1yPt6f9N
v45QWYcYKUZ0VodqtNWxBH5kYqZNIq7bi10bmJhKqzfYj17dpYSdRAim6VD4OSITkR1RxjNqXsDS
TfS0hmphc6cvljz6/82OW30uQH01DumvwYWoGspJTSb18/1+OXRnPQiPCieaNlcgRXzFOWN/Cv4j
t9klacuIhk7drMMLJ+rO2b9oiBkdfwE6Gr9nHB1kcF32EjGukZsh1LFTR7F5AXYuyuhmVoV+O0a3
SBW2bgxdMOW77V0ooEoSssaDV3F5Tqm1SdliWGzZ8BTGLuHCem76xEbfqpiiauunAoETbOs1NS+x
IniPL0fiX7Q+bDBLLN3syYkgoO7M05IEG8ZWGgasHkLdomVtbKsDwI6y5itOVoJT88G9XjXIXmor
rHiHksfkp7cyWDZWfRbq+0zB6qNeIi1vVgt+g1J4P286XxHHPoP+BI8YtnZ5FQd/4hT3wg/xEduk
wwNUCqgEBjFQ6H34MHG8iA/Ceda6U65YHdmiQ/6MtxAeARV1KMDCNkAShcoLSmgFlTAdAcnJZIpE
uBr+eJZz3TNUTGJCfY5lxzDNRCc/L2oC4dzSB2r78EEDeEcGqseeVNKo2QFtHJ+Uu+FVACcCSKmU
bGVi1STuRRGOshU7+bqk7YsUDICmATmwxcbgPHtUJLRPhUgcFIxP2ubnJU7qkpD7MlpxCh2EpWcb
Ji8q2iZh6Dr+lCdeM9njgomed3tsR14e6L4ThZvSyJh6g8cxbIlax+71vY6bMQjEoOb8tSrjRUuN
aMmgf5//NsUnavOIyAF/vj1FisaCFk1whR6wHwtdJJphApge8fmT9yON6LZ1tejfteGsz8RcE5db
nK7FoSRj1jFCCSuNqrX5x0pEcCuGGmlYUXrEMbf9sdIVqwULZDqeCJvlo1asNvVFSefcc8I54mxy
N/vKe1pVTFDHAHHUtYhCwJEurN4nzbowfAN7pUJPQy7LPn2QxhR49nEykiyoR7Y2YU2pwgJNfPav
x/ExQT6lrBRRUC52ldUCs/TYNSKU4he0pb+xrSAea50kkCWwtZWiIqQ/zTGRejFmHqRwzOay0R0w
Kmpsv4iWXtYGPf2Uguz/dQ/7IXj0eP0mL1DKySfAcBBmVRFNvPJeo6O8WeRVB8qU3sL37J6jSJNm
LYXFr1KgLQt3M/AIZG23B65BoZD6ossRch18Al3HQvZKdpPTIK7pLemGNxf155yw8S3N2jLcjhxB
2+x+rXyU/rDQVhqiFXkeyNdUZC8LgpmGtEl2eLh3jhnQaA9RlSQWtluemPwbXHJPqJcR9mYJlyOy
PMWEM2gdEwaTTtvxbaO0tqEgdKOSLkXfxwOA3q918qo32HuOiG8ISlsr/jDxKMpavbRmNapa5IC5
SVQBeRstDlgUQRTHs9Vmu9w9++c52u1uxGepX6Mw5xEs9R26XbChyNMIfdojlshNYwxPBOKkl/TL
ctiLF9OebaGO2Tu8OUk+ea0TiCiZothqLdcUEAIH+CTgBSLYStOwYjHXofSDfwP1632hjR3BLPam
6nJfPgnwWf1pdUYkKYi+LMps3kbBaMrkH4k97bd4YXHeGsU/7n069z9MIbCO8YrqKtJRbJaXj0CI
eX8uJn8YbMMIPZhu4aCtT4cOr2j+bDSX+nG6x8Py7wKV4bt+RGx0i7fy1Uc8FURmXSQM9hzSWNPv
4o6lnVb8nIizfnxIjbgMn7A7RDGzmjwHqc2kM/TQvUArqurkGf/kTLt0k04QsYm4ufdm7nBziWOr
KvGDfwrWcnFwP687oRS57IZqWz9CV4oYkCWMwrF0AnHpYjM7YQ0ctgJYcBiKCpHSdEdvVxank6eH
fDICSWSKwsjy/bpc+b4yUd1Oapw8sOhXXGeL1W13ZZndo2E3NjiImduZN0+GPLMQYRolEiZJfCue
AtnqOPOJ8TjjAU61s9G4SWAUJlAIG0uBkPTeRFSO0sNcAbneYPRwLe0oR9mK0e29PWiCWNnwXGyY
qQlkQp+QwBDylQeMUOVia6AxHOIgzMu4CkINhTsokl/NNIfOpgGV7qR+rvR98v9P+EHncZfbbsOA
tWaJC3vpMY+s41/+rLZ95vEV/5SS9dseHftc3rBi2ORNmD12z5c5QIdEqj+Etui3f91rhD4H+JBn
lSplkNyyAGXA3j760JjZIcmLQE/ra/l7kVnoumcym9d3rcDy54Z5zkPnCvbwj9iUpBcv+uiP9Xpm
FZctC4359yxJmbyQPccs3t6pt71KHZ4xWaWelQuNw08/MYPFJ6BSCq2dwNNo397pLnDqAJzIc/a0
WEJMLp/pd3H/V2tteXM8fiELZE7dqdVKLT0kgQY6jYynyCfp4/jCvsy+fa0MDAbIv2lJPYi2xdxE
tqNmrz6tQKsKka7HN+uaMZxm/AWvqFEUwccr/Y6ZJJJ4TnFDzcYsPujj7xKMqGZehNaTMBCeAB8h
4Ag65Qm/9aIhelKhLnxgvmGHKYH9mgCVSg8RWORweoHlcgq2QejI+OAVbov/8zk0nlJEWkLXbEQ6
FgfEt56oF3AdJn+kkIIHpo9E14TvmwktnxEA3IVr9ORAyiGS89aFbGquU/rx0a43df/dcbGNjUfm
eUQOSIuFO0N0xqSlvykEHvtT4bOVl+cQiQQHTL+0e1AeFrCGp0ciEBemSuukkQdnyeWnROaJEfZX
+S5NN+0qbq5m8kAOwTHtw9K+xA1CWTeIsChRVpH6DU7c0zAeWMKqn+8Zo0lyn0KyGg7agcaonPpk
U1oPubtOnrP73go9DrA3cv3bs9hTvryFocCMnO68aK9gvs+OvzS6EeLClHeXYbNWPgvSMlRYo1h8
9uOBH1Bvs3+rb0kzbHuoR13LymQPDNuXmoghm5bbVj1PwrpAOwpHKqR8koVUgwSlyY5a7w700FvI
6XTi5osbCxyXhd7uWuNFtAkyYbFJGB3emiaH3rH9o9cghECAC8b6bHpn/JlsmNMqSDju2FAB4C/w
tjGuWUfTSdmwsk0tvP3MlD3612qfz671qHvnQvKv0nzIbI32T66RBWIySmtLSARtM08CU+yHSPAr
kfBMSKc5DTh6KwmvlkPVts+cIKsJbWFGj3bJ5lYGMKgYuBQJZlQdgFohOE/y7HSvQT+z8wAVsyFh
oTks5dRj9Sle289yqlKqfyRy0iARzqix8obvI4z7arftFQwpTbuD0uOnMEnNxcgWG6K2V1t87PAr
nAlbJqIJq4TzHfJRezrgkQO3oLs4jNCAZc2iTPlSfLlaqx8J7c+5M1AvkLfh7mXBklWl7eHUZ/dM
YmgEoZmMY8be5Ahq31GAZYxZjI8sH9lrGaMWHgVxjGdkjz4Q/xutc0EmYwg5Et/wtfgKe3NAYhWo
kcwg2jsB2Ws56d1HHANimtgxvQdJNnGNx7YUZRa+Asgh0wYTx2jyn7XFXXkC19dtBnSE8edFKSBZ
/1/lysKYE7UuFvQQZndo8b5o3x3iuLUcHT5GRZRnrUDeuj/rcTeVxdrYOkhaBFsLqJ8Zhiei/xuk
2lY9jKPAcD6TSdRQFmJv+RICoQCXqqAPZkufgxQ/WpI/3+skQvUMBPsLvf2jZzw44z3o3IY9mTVO
+e30D6rW9d4xyAGRO6pIcETx4TRTjCPH3ornbXq9GLmTPULF1thLEiVJQ51iZQDYYMeaiJV/KbuX
jkMAjhHOZI9MZF6zTj0RPC3eJGTYcdfN3cXdp2Og+Kb6SzTCKIH0uhr2dLXSkeNqAOutJaiPfNv1
cp9TnSzuIBY/kJkTaJdy6KwRdprgQtxF518lAWVieUQ7OwozfmjC4uzrASIT5D6vqN9pfQ1gtTS2
E/RSAyT7Dl7Q3FMjWfP5AfPChpUOetj3sluvZpNujMK4YzoGUewbFaVF4t6uhS2vV+Fbpu7bNVQe
hOiObPFk3nxFWQx75p4XcKw270MQL+6r9yDamMnkwr7ydEvXZi9HFATStbQzRYlPlP1DeU8Weywd
xvd1t7ndrt4v0qVtnHAqkShjsUDbZ2LBDapmZqMrFkV9TTmbRpnB6OpdMR1ekH8lH9d4e9SugEMH
penH9WBZQORbo1lhKuQ6bWjDzEpRnxQd6Va7SWN4pJMD6dqKKn+PRjLiKSLErPaYAT6tfMwSvmkf
+8nCSu1nw7+5iZ1kpDw7N34Mk0RRxXI6naBMUQjzhcB20o3jKZcy+YApMZu6NaMyr/bKbVxmWVXi
kpkt3bLGsZJsFW4+FU+chTATAZPf2oUmuyWTIcSM7M+MZINCKXpmoQxoMSBsmtnbW0NWGW77V3l5
XhKgyoft3wyy/ypWqRv2hlP2Q7l5Ndk5C9KvOkGyoRZXrww3g+j3SNn8xzsv9hlYRHKFjKRqOO7P
cdo2HLxvFj5uU8CxlsEhnI8Q8RNjqYVxgP81fkgqBtGNQQ7Muo/fU8WNrujTMVbGXzGlTKf7bfJk
jTiXO0+daVxGxw68Gi1BbDlnZBWSummO7InTgf3sLnKHBjp2FWFvPXFvv5WU+RE9t/wR+uww9f3S
7Tt+giA4OT0jiEsqTRRfGUPJJPxj01vZIVKvBnShnNi6IxQap/Dj9AkqlkPybr8YHv5RBOSv8t24
vvV9sWBik8gaFeMfntKTiY1aYV/ngd3uzW6V/H9tjhA8z38HtA7gXCLSaaMohWKkhhFf5lLrU4I8
jcRWMBp3stifwD7mURIb7j9aKUu8fnqvKReJTO9ImrEt0E9JfvB+UZo3gd5PJrjtvoYo8R054ET1
ZYaJGwbhNpucLDwCioU53jV/a3kXDbxk9EQ5Vsl4unYs/Dg4ZcrcCixJnEUig6wyuRSPam8W+8rE
vNzyOcSqRFByVCyFLZipuyxgdNf2aKVHdxLFp0fw5ZJTr/TAbdnYIGyHMRgivAnA7+fLOQhLy/Zi
sOQpXv87CsBDn7ehFT6pWTUR20FZzTBZ1wDtx5wAQHxZes5n1fG4PeoWTWIX1Upd97ytK+5ycelc
Uo12fP0uMZAQsVq2Bpdaq+Z86RJmWoOe96dCpucsXOhGVoz7OxtbKZm+aqa7ZLLYXmKSw66bgKec
R4RR4WNnoMQDAwzdxfbH5/TVW9zt4Ojn6B2AC4ReQMczm1SCx1L6rZKTJP/aRro8FZQi6AGUMQW2
1r/6QQN1WogPMAdhXEMB2kno0vnNSpz3sL9tUY1bKoBSCPOd7YTwFCQyWVeSw9dZJ3PVhRpehtsh
dl6x5MqptEEsTps19sOxHNKo3z7LddYX1TmfzpVEGc8mFU1AQTmlfE4xx3mAPw7z09P6OAHEdTZe
QynXjQtZ6gZUZWCKUaER7BrXG+iKN6kp8e980GoJI2lRILJ3zysrVBvSAZGqJg4ebFMrwIrKVFTa
jDd2HJ2znvNeHHeEw8nTpxJ3ssdVnJ0UlmG3006zFRJl7V2k7wZj4Xxu9LrAAaz9TGpUSlX+pFsx
nDAy4RTGYhNVfZuGZsd9Tdb4F/4nODDrmiintlSlW5/VFBPGaHbvicvrAzG+WqyLht+fRiq16ZYc
Jb7CA0od//dJvk4frIYFPmTn58YLhj1H4q15MabWuuvMdHYkBDOi4DZuJoiXzHuVdkxtisVh2hWK
QGJ0XX1E87pBaPuwPBoNfrmi4r6StAWo04MWvZZDfMkVXsWRyaqHduC3h1wsKQJbAQxNQX+wtiTd
qNkxcU6Metuc+BTxJTTjvhLU49pu/iQG7JDmuumWAkWtGPFou4nx61mk6CScb/G+5u+fHgHKuomX
/smj36zL6LgUt8XvvLll5jAwJR5+sq4u/D/ANPz0kAVigGAj4NJVZGLnmX8/TXtJjTf2Zx+NcOEX
p4VkfQBOenyZflidaa1h69g73atpjSnZSuC4xBGJuKTI56PSWyso/Dj5UQJE+W2dPERMvkjBa99V
pRGw6wUGdfNnbty5Fp9GPWcV+IA/S70aoIJGM0yDXUXWg9GyFTYxj82nvNxbYig4IJHTLVBgDayb
P9ofYLay+djgjqHUbCcZiUjweCRNbP/hzsuHYx7zZ7I+09i1IyGew+73RBJ87ZkIlapM47k5m45X
5jobtPp3a460ZjMy1wN0jNE7SG6bBwP+zHScbh5q3yy8nneDpWrbyrlti7nX9iDbSauS41vOk27o
hjNvcOBra9ITHDG0EiGQJtznAJSiVS/OrpV2MdYmGxcgrPJ88Sh/LkYMn8wTXKJv5NFnMkvKBN06
GX4ylq2fGelpai2UDIXkH7hp12/6i4QbayAB9ydCCw9X+5/X7JrP0jsVK6xfJtJEUZmt6mctAXlO
JpVDA2O8ufQpYxSKVtoFQ9LCaauxaKH8p7CYXJ4HEwQyHuwdbp3xI0x/0aW89rNOFhbRvVlLEFbJ
zlgF3dEVWZa+hxqEt3EeAS+JtVRZ6H6z8FaA5R76SAtR0zjyp/gIQadbEU5tjL5R5ZBWqUKXtSyB
iUyHBdKqws0DzBxrAtVn3HAcHx50OCs2C+S7UIVuIXl6vhHYBFaLtxN9MACWEKhoQi/2LRlrmxuq
MCynXN1VIYINFjTfJWwdyYhohoQEKp+JN9x6YarODsF0TXyu9ZgkxEiuQOR5qiGL739JJW+RAyk+
L19KR48GcpsOSr6BIYOVRjQrJRfUyxoGmBS+J5twdE+ujqWJ81wh+xvjE+5DKMpzBmI9vstZ4oK/
lem1dVduxSEiERJD8403LEZF2boyHpPO4GiNk7E5C+QwK1yfUPItTAB5+rj4CStpPFAG3RDEodEx
qJ/Z7ICmatCO/rZDBhkHUX+FBJrSY0w1qIovzTRjZzNYTWpURZsxUlmsY6Bi1TI5N7TuDOX4R++e
zmwJZjiPkXUsglQGuYH5afnm75r2BGZPPVCnneeYYl4HixziZ7U20ZRGq7AsLAfaj0iNoUZ23zgv
LV2eJKLWHrD2SsNae9fK7sBdMQCHzEHxwBWADEngO134cYE9P3o4Md59p/lrLHX5NgHKcvvPb2r0
1ZtT5DMLVCqYDQS1BVJTcnqzz0HgCNLC3p2eFRec2JevlSacKIE2uKLeUDkRScFe03vkjLR0sH3w
c0urQIefCtaxfm/8O2SDB5r3dqtPh2xhYlQ7PSvQnYYF7cQ/EMwF6oXPTanhBZHCEOzzzRH9E6g6
AJK2ZpVKZc9q2ny4gtzBh3fsIJkhptdpGeaORrzP6C6jYpAl+fB4+0RzoXq1lNouTRH+KccY2jZG
IQtsLQF9pjfcnq9LHKozgV9ySQUYqmUqPoLJlj06TGHSEUx75KCp37qfc77SvvzzaQGnB4hoRsvK
NsBZ+smts/ufSk881JPDdhs/wz77DwU3mWA3Gj7Nl+WWW9+YRIsTByllSmMVoSefZuXXhjtOWMJw
DIb7M3gCqYW9aZxY47Y2IqJi6Utm1jdCPQN2Xev/kiBupyK/zK0ICxnx7cvMJrBOZZt6Yl2SGzMG
FAC9BsMYQeJY5BSBMBti6cdBJgNzjIaBTdU8hFqoJYnXkIR5XU3OKhv/bXwVqEbb63hFCZWOkWv6
1nPzT7nppxrIxn/m0Y/bRplQhEx1ZNGxRyICGa0D2uWq4sRVsIj5hVycnnNkJ/u520s8oy5+d/vA
atYHaKRYDh8BWaNqKu2j+D0uvfHbeLaOPtoVaDTwJNrdAmO/kujGPJJSeHiHVEn/v9K3vqL/Wt0d
zXjw86TbAz+RMqI5ii1NIjb62L+8GyWmoQQvnYCQcNmRRkVKp/DusO5JNVdMHEfMutU6/LoWbWyZ
syIOTYTOwhJ5JdFRkfi1eNQgXIGbSfDKCQUNt6uMSUUIwqgjDcqVoeNtxJhIWPaUQSwhKmkzKetY
8HNFcKKUlSav0yajJOm+kB6y/+/wYuIqRLO9w4Ikxe6Hg3BJ70IPPTJP68WJsCmmF8t4/6oYXkjj
OzUA/hUs9DfMevhNI8gBH9IVc8doBUxF0/z8b328c1XejyCtFadEne1BjMbxAvJxQcF+501eswUC
5ojoJmwXjKdy4pEWHWmiwwqS6daIlqjbuVAFYDs11Vb/m3qoqgbCIm8ROSyiM2lNB44D1IhYzz7k
Pvm1yxdXoQho5EIndA4JiZJt2EA5tDCbaZ4FWDNKl+luBJrwdObFQrjYgwVnX7EF1k7ruGQt86Ky
cBNaJKIDhLFA+3vrIdF3rdaDc157zAlTOCPpaB4xbLkvnVOjygzwRC5MjnPZr+GbQ5DcmP/7vXaq
J3kCIQXoYgCijGOvkBufSg75wmjY2dNYOD+qV7fuWklR4HIgnxnhjv4tvCKmQh7lC8WgDKPhykJo
kKPApQ3FEXNt9UkuM5R3DWX6hfO2SK6/vVJWC8RDSVC5zAtQJURAbus5SilUm8wf67U3PsMJnOWe
qj7GI4Odsur876rAtwiL6ARD3SRriMkohBM8qiQosb8vEgl2d9HcbXTq9+IZbOazgaIPIGsMnsn3
jT9+azsXEhOBB30rE9wFGuwf9NSORrsSU5I4JjcNGCRL5tZjd//SkNtI5z0YAtCnwXgvrR6sLZGA
bQ6smjgJ+pTYixr+1rXNRgnEveY6l2M8KUjwspYHEEoNnljLW7BnMDibbR8zE2F3zefxmq2A+wlj
zF7PNxcHyQP3zeIpeA5jULX5sFFI6WMV6fJS5WfAOU0gYTIbcTYW360jzDvBRvwk5bu3K3VdvCJM
FzvcmuW9RUiVzIf5Kled7Pi90RLkNoOoLh/KUA4LssErOq1WCo5v9P35wuv8bBFk/7sW/vYNrPLc
JbanOKfvKf6N78ukFu/1uX2SWaPE1qA9SN/RC9UF6YkTntVID/rGyBWbGxU2OkNrcy3O/W07/cRn
PDBsNCJEID7GCxYdXFREIfzRqGjYuNdnOpthvcKA6Q1grYJ2CI7N+DxxB09J0LD1s6WKvNraHoL4
msCsNLb79E3cFs3okLEt4nxl5eifrbH8scykUB1A4RZ9ndstiRWgCwuN4mkNYsmKlGQN0FfuUNNz
KYjw0rnGBRQn6qBozbwJNnarKb2xlLuMiocxt2jE3FwPmZ6QuM5A6FYluUcEIYasYLaFlgSmXL0s
Hcx5n8/JSVh7lBmhd71MOIkDJvvg062oFjV90FVNQDJKM7+QAGE1g8JYOMihebnj+J2fTQOHHPeU
Xw3NEo4iohRz+ezQVFKZqa6iKZ7LntNL5cOfTkU0IGbu7pehAVbBVxwpXzNe2Bb06OdhA02Nq/Iu
2BY84j8Y4jQNeTZ4D6ywR8v5H6vgZIMhmG49+WnlKLk0mqDJL4u1CiQfV5f02z7bGSmLBLLGbRVI
oEt37AGbEonLU1xriyQbRrynFXHnlekGe4VavCajg3F3WQXiScZL2klC0By3pC4Mdz9OI/EUqcBM
BBQiorznGKcz4+kdPffpDMrCN7zXxclH40Fh0NLPrna/lUiaDh1VAxC6azkoTmolcYMdTuSHejcw
5RdyOYs2i+7tDwUDaMElouyN9QnEobiM4tPaPXYMjPWOJ/fGDBgA9IYTTqpfPqju+5yZhjRP7fnA
kwwxAlMl4Ls+38qZCJZPSW3vAhYW8+1R3JkkGPNIwGIVm/rVx6CHkHi3AxI4soIeW8TxDGwtC0+P
blMps+rYYTbbFoMXYEpAlo3uf994DEWCiVZEnzXjE0TTJpdIPOdKLy+EAY6F2idRvz+iJejzzCcO
x/Hz5g9H6P/SWXssBbF30U20LSJRkl5yRebB9WJjHUKbgx7XU72b3cg6ABT0VUtR8t5AHnTRGBD2
xbZRAz4gpEzrd1vdOcrZ74QNiQFJj54z8R6yrLLOshCE1QwHWW2VHO2wwHpCcrPYozsPMT9w93wd
uClRXxjwBXkZwtSVYnOtzFM2osuknmylPjStIpxpDyZ/XgGh1NoiCcXqMM4EFHF5qjMA7a2V3fLO
OhCE0XK4Rl4/2XaeCXdUv9zw6XzK68qtRm7h7O7mik21dICAZo6WZvEWgPaSwu0aDknyInxmiGiZ
wC5cW4GJ7F02Csf965N2IXqeGzjb9uM0zTmXzzUItUT/aos90Ll6yEFWR8CFo+QOR40YM3bwDLzf
ddIyejPKSeOiZa0AbbtleZitxaOUaBjO0jiZ2fU4pa7FGqglRgUlQ6l0Khj8ivoijzadb9oeaaxJ
x4KnFDxRAD2HmGjve+5P1drzQM+hxh27YFSTqTL3yHNEPIxj18g29auyqS6Z+wx1Ch1NSGELoswF
AxNKwZXjD3YkCdvsvwfvz6fwoMQJcL1zJE5bxQja4Nbpi9REbYiXXVcyiPQW4uQTHPC17UPej07M
PFdwlU5lv8d8UzFrPLA4q5DmEic2B43jDR4K9ZtVwVzg1ZtLc2PzBgcJiiOkrMygs+FKY4kLmaOz
oiqdG5OGzmFMysTP8H19RafofOxLcVV6yO2p0TGu4FpoDoT9KIpGZrPmLhUI+K4J4Fy8/pgRAApI
tCZ0MAz1i0U9F+2eZkdjRwkcyZK1dbcZfz4oS8UzF46tGykUMDmTCYx+E1c7BS1q4HBJST5p1p0H
3siHOWshRTdKeG/pEEso+BtkMFmUeWzwCzP+jObWhzCYP10rTetK4cFtTeSKhP40667EUy+H3CUG
fdpOFFA1rrymbieesnJ12l3KRNd18dn+/wVhlBdj0YMsgVuinMEWSv5cqF5eTlsSVPEuXAInyvHH
MPv9ru0TwA6kB2AURbpOjtnNME1c2j4WyQeWrfOjNi632xLcCN6yHNOMRxpOAUz3uVUJnrrLnHE4
gZ2C5j7nSpDhrspwGlh4jQeQfU00Mhy85MfByPJUMGDcJB3+gI5ZhnI96gxvp66yecUfjid9yQH+
WGxc4bxHkRk1OkVQmqsUDShzPARRTEFkDBTBbgYXKSmi75ElGAAq7hJyj2hoqQ+Wk0JrsP63MmFF
o3+JfPvR+4lgR7IaAStfIMgfbqppFrdgivXQl5LPOP6Vjm1p4GnSwvE4Nk493lNJglbjQ9ItW1Qj
AJSjXu90qLNWgzNAKmfBagrBua6gl4ZYDrv3nitP3mIcsrYZ2rBF2F98UTMandeDKfR+3x1kWyR7
NmNPnn/UGBuj1A9Dc6e9QWMLNE+uJiDX9OocpBURMr0SuM585NNeWvXsLznbJ2bWjmCuAtxHaonK
qFmMGtcjJlLk5NB/rf4rGyo99VHCclnivmmc6Eu0ziBqDHbMK/HkQRhC6CbZ0kHNri44Vu5fuebJ
yPabcxtLxxzNofcIFdlQbqV5sdg3aoJIf9T5fgNBHakDp3P+AY2FnTZTD5S5Phrr2wa/WjNBdCWo
CuDCb+UaDpABsgS0xEv94OBV9C5uxLzSIxnn4+bdov9uRRYflrPGMuY2ta70QVrB5KICxDpFPDE1
EzxQisgD2dFF+d/EGLoF9kdcFYxh8GOgp3lRTzKLs2H6j875jNmS6tnMXDFmbETuh8rPjp2P8xwV
dSNRwkqpz6tZyZVrWcNOhHQx6EC6TnoUS+jGtQr0Ob7JW2ov5JnqtFXyfA3eDrPKQx6Zv9O45vml
NGgA+jmhMlfyZAt9ybdsqroaQH0uw9FvzDD6H3P8ZLrQH7LMX3uVQ+276MdGr7Fu8UKVFs3fxSsb
maWfhoVSPqAzuZIW7+1zh7d7EVBemxTlwypoJKnbmUUaCG4usYIhDeiyKGl9P46/LhMTCZg4hfx+
dlprR4hhflTUIoyE2EBa2bbYy4NrS+EVTPirSuNvB9Qd85AhiPdi2mAfuG7c/Vn+fHT4SNnpuE9o
pVms3Gz7jbzcD4YcWk6mrfW+U0t4S4M6kHoHK21ySokgVoxfHALlLuJyPkj/JISwHPbrY7q6YySy
Fzg9GA9QnKE6o3FeIO9m4Di5diAyyk+LUeL4f+0wCGvJGn1tAeJoLa7QypBLrEw200oxQcmtOZpN
jzTTTkt5n6hlgk2KkrajtnGkcPwjq+i2+EAqK5NFNe2/ix0lrTr1DTdi0ymkzmhipfjJyjweuKOG
S0NDyQHlDR32GQvoiAzsU8mlRGOdYPYBS6D1QKInVjzLrrxpC1rwEKUb9ieOYr0Gphg3+ouFNbeQ
I9VUjPkRwIyKA+s5vRWVpJ2CT7lCoA1IKXOE0JjcOLUAdlEGUDSQXpRStjj+0WhcdNcsUPQ6lUcf
nebLY8oVRohWofC7e9mVecGNrtMBP0nT9bNQ/fiYe/LafG9pkkbWnDP9tKbnQTqIdCOaYFBlOnlA
qgx7RhThpbcIisJMI/7SNJDrmkmrvY/SzPitn9zFA7UYNjNsLy4W1Y36VCvFUcIlppzVT6W9vP+T
Pv3IEObSglAL/crJfmt4lnhjcXrA+VDDb+57Wp2jmr0QVxTBdzxkOXvcvTzgZUfqDmUZ/6xvddcx
AitACBSr2j32o1CGJHf08OaB7lDw1fnXToyGRfSKn8hdx0IW1J9ZDl4IXtqfG9hCw9wjLqcHZEv9
8mi+6R12BMHrMjHJ4wjrxHWln6ZDbiStBmuyBJ4L867T35Zsmo81RZm/cCgova8Yk6NtW2Y6u0t7
pRo3a8MUeqdbNF0J2AIXQ2MIOHAPvJbLLQ35oFEqhIVQqXjuczDo0OnHcQIGHauX6DAk5Vb+pPxs
POvrDEhIt8Rym04ad+5ZC0nlXDZ4mmsvQNCLSv19EhVDrHEtHTWyABiPWsr2AHJCkRULgrP3vQqG
XEQsPbj4mbQGKYlB/99nJyQvRWXJvgu9Q+vgjGxfDQv3/zesLmfN67GMU3pc56A8ych0llyeY6P8
1eGk9NdwroWgFmQWffAfem61Aw9sd3D91C2QLuUGC1uB/BYtTdlF7jGbbxh29+DBVecfTCOst/Ot
ws2lh4/cBU/Eyp36qFuIYSbyfZttOgW+sj17756gFbCZ/kuR/W/bVeaDx0spUhF3i5jLCSRgzbQ6
JI0QrEH2cj7Goi9NctL2JnNrmjV1VRT2Th5xfmQIzLcbuMmS9m++7I605W10Caq42QiYiQNudi0G
V7s6U2BUuTJm7rMdLbefArvFR2gKDuJeM7UGC9t7/ZqQEcYCf4+DGBp5tZeOJKgUy1cqL49ILyC8
4QeXSIpuaJIkectJnbT5Sbq0pHlRuuZJWgWwilGAYVxyRb31DovBPitWOD6BjNrOOYZyfkEogxCi
75/sp/66k6GyDaJhU0yMnfbgpBlkE5EtMpLCcQpNmuz06n3bg+Om6/CmIesIagJCDOcaM97ZsIeD
osvO2nOlLSDX/5vGxkkMhLNTGh3u1AqVAT1IRuWt3e6mUQ+nPtN3VCwdaJBYOpWm011tVTeeqdo3
VCEMwP6rP83pbCmrSmn5YrqNw3qpDp/wfHXMb7NNUdbZ/OBJKc6XVXtWFQYZBKyXj2pOpAzApqqm
848k60rjuwHPON5a8owR1T7be7Kl4l1w0/hdY1h8wv83ED16OGggzQ+Ij4vklnHaFvq44l9WHbem
nh9IllDVQkP2f09CD0imypDD9INyOLwIcsWuJCmmDz1FaAUVYv+U/NU8iSsAQQ0Lvzdj4Ha2oGDb
C72u/WS+cYf2Lde+8swfJ2H29HPERyCz4UaiWIeWVR6x2WZdR64qgkngphrdxGQUub7i+tkQix9s
Bexyv+9tLo3sk35uW/yTNuTi9uquROtG7jSf706H9hdqPHqbDCJ1IBH0V5Do/I8/bOgPir9b1d5N
5I4FWe01kXbOedrBjzkA/iDz+53+zGszat1Qh2tGqrdiis6H9pMehjRqP/Q7CQh3etTNxXvK9mWT
umGJL0MSl8g7nKOn1FH8FsFAFueLSAb9rR29/vocB8ityBNUJVtID54ZGUTjr1JYpbNAOv6/w0gk
QlzVE3Z4B2zqtPkndVfU+FCsIAvfezZoMVMC6ObgyDRCc7zK67JcfsIo41kB17ZE671JqVB2FKH0
GZWBbXOB7QAYxg/DD4JqbKBzkoHWO3Eva31TunE5lRIrLV6aZBLb3DV9EOQddOiO6vBemvVO5c1x
4UUBcLc0G5fCZHwwSjzGDfH9GUFCvWCJpSKxkiiRayWzewM4G/+7xzbKCnXW3h6d9BVa62mA6nVT
EaICtHVcQ/RZeE+0qLxxI5teOe2HIgDTZb6LRPPBh24ziUquN5JZ19Puy9qUT7oGjWkbZIf3GBNB
ab0VwF6N/+7Z515TmUa2QepwDjHOxznNzuOAmem09IXlwYj226FafGO8YhxznIJqtwOyMbxMg+iX
Tq2ZKeEGOfoJZzkwP2Vm+Wx3neOVIdEzwSAAI1tDyzABYmspB7+WXvhZtob45GLcmouofos/1YSW
bSI6oBRhdQASxYpS6xZhM/V0RjJyz+lgaRCMGz5/xT3Ff1naMMYcUXrANuwUfNkVBHtPfqs2Kmmm
Ae9V1EU82GMcQkmpXZ1McDN/0F75KE8gjhl3n6TPb+xsNgUtqEAsgGAy3pJmpvUtbwbdn7M6rAMv
mcM6ZWdc6EiF2HbMXfeISe9cFJme5ExwMbGHYm0GXcMvFwPtP+TVmMxAkMBGzVtE+hjsoIzE+3rj
yvCuS+wHL0WjFbrXB5Cm91XXvRH7z4BJ+dpD7x7ZvXMFzq09eKOikefgv1LDvvLCGmXykv4lP61/
plGG+Wq6sxBVIpi7iE+JXi9SLvWS36EL4vOpcoI9YNxHDOypfuK9Wil3l2P6njuzOY47aH48nWQR
36xUWMPY/1VzahqWzuznVs1MB68WpaMaXaD2a8kdmSFglWTgMYQGBM66fkOy1o16/3mFpfq9eTl0
+Mw/N2KuXd/RFZajpbdj/vZEPY952HskIWnpNorvaAsex7oESJGkC1w8b/WICKNpsjgnAK29LUZ9
oCsZwEfnZYxvQBStBJjADK5HLSHE7+pTrzG+j9DTvGDNY5EkpOWQzClycNt6RzQU/KzlTvf5pUEu
WuS066jIVErfil8gBkliL5zu0jgtM2v8rRpf8LUYyPl4/T+4kv8Fxkpyen5OVpUkySu4+3q0QV5L
Zrhkp990mYzeVJFpKZn5vvDL0BiBFX1yixC14wwgACsm2ok3X27f0d4NCfp8qtK3lHdLpa4Hy5g9
0z3ZrDuYFvEuiaR/eD9p5kAauN8yWsuzB+kmCOeds3p4B1sj3BCWWCLE6a1ZJksEgFZqOV8s8kbT
zJfsHD6Vn/8c+JOlB1S+2acBQ+YkZV7oaOaYJPWPgqwAjX9Mgl1oLwzWbT0GdOkp4Xz3lJ2VMzL9
AlgVcCdq+4hG29pFs8Ti3omKvqmsjunAuHS/50E3obJ82GL55L+pHyqKcbtAS4KCqNFU/bR4iRMa
KF2nyviyrYDlOiPSN8AZ0qkJ5nWwTgge4qZZhqoZGjUa0feOALkXN611BfzUXz38OFQew9qSlOEa
1ziHFpM1//w7yLgBOu1NcGYTekAp9dTYP1DUDXS5nzYj5LZdOI1cwGfL3D99K9mhv71DdAmBOaJJ
O2mE9fKe0gYZphfAqrtlGbjO1xO5rligU2lGi0uE6ukzmb4NlRtnBRBdje4mp51tzP5Ddo3sRDtQ
nQg86nerh7mjstplFEKQcfxbHBwvN7gKSQcDHkq/0cvAE3OyKolAND7GqOcwtinyUbUr/7gf2aEp
BBdNMZRXd1pN6isf12YY9GZmNIm1SzCm+v5QeusVhkfrnZiWANXjp/tkDgWPRSOTJAjKemBuPvY4
qh0GT2mghmQ4PXO3xiJMOdmctjTZVGXsJmD66Ux4wyFmYz2Wm5kZrT8MwGgAvZmcQFOGOtLuX1Di
JmTeW/QZ4i9UCbsIUlCaU+V6FWKKATr3pU3d2CX3EqWjJBMvB7jQTIUQlDFJ+gw0VdV/UNW5SuKF
iTVaSwjTJIm+BCWQEeJ7dkZN0lpPoBZNCqFPbGhVM+WIohiMU7/sXW3aYAp00HFALHRqSWRtBsxn
F/dVBuLJw2reRpTUKtrpAKrsg8QHzebEJFZZaL+chRURJKCN7XLMkLt36LDYsvAeN4E8vbFf4jRL
j0JQ0wlHXQTMh2ItMOhibV8l5ZzIftQtEq81Uc7oGHLbziDNRfyuSXQSye2NYSvR7NF255zR2yeu
q3Y/OvGTI5h1faCteL/DXn2P+CtKIeKyn6fSPriqwC7bOlYCD7/pWeFmbcF7WIDEEjb+O1hWs3/F
JuhnJFD877+IqXBs6qPPNbUzQwhA3VkJaInkp7o7+8R0mSYFNc3WpJE4uMdAtbD5ElCjjoDf5lgr
7wFdNNntRQrgooTwvc7FOJN0V/yu+T24QFvMm8NpSf+qDndK4MLe/t/ke6GanLAZTCNqKrFWQsvX
akgZA32Eva3kkamk5Hy08eC1D4TYFY23rnbdoiaXWwOg/fQPOM90caDh+LsN0hohsxtjUAqaafGW
Y/W6FB2wbhk76l+5mVYX/KWYjUEYRxh9eXQmCL9JoNspsv3OwMF1uCErURwiJJwZ/S12Z/tlY9Aa
wLbRGSm7cse25Trg6PrQ5tPklbnik6YLoWUUOFqKTQ5Cy2mIwip6H7hK6+QUTfwxIsCRK+7nxmve
mdqaYygPwcFqgqTP6dNCIBbVkoqXCoqy167bGxnlayxTwF5rhHZcRyW/JT8G8BKGjP62wds6mmnX
Fz8P4V1Y6evFqrOXDvGogxvoeYeFZg8Kl/3ovanuMH4yWjJwitDSed6iQ/vbLZYSU3WY+1o9kLkW
r6yxud9zJbtFyUEGiD3nITOUZmHQXZB1bPcIG89vDz7Fd/ZmFFqasL2T10RFSl6nPTECbS1q1voc
xf0c9LXrp23HEa6VvymszTiUwUokze6VFL4exgxsmhRDbdKYF2MSSlpCO+53LnGeUfZG7Ih7Rppy
Cyqhr0t4/nbxch/ncJTGa7eK4Dp9BhYTdVbRHQAUEF7WqiEk6ijA4YHeAkbWNdZu6J4qhZlmD91B
z8bo5Z2RWoRPf914Grrp0JB66ME0JwaaZ8TUszEaoeI6t23eAIUURQ9KrB+S4mw2Em560BYY49DH
LzhsWdFxqBNRfdiDwSAswfr1tObEw4hvndUilTC17WDpmqA4wE3GRS7kuifY9z7IWZ9eJLWqHUrn
0tsEUbEEVkfHP9GpgZtVxUf5TyhzZi3J/zUFdhueRzEw/1m9XwpsQ/7wWRxHShxhD2uQOjplkGhG
5RrNnOLh5CN9Rfx5I4Ic36Kl9lkwgAhzHl5I4kiqGNM+urFmE6pzjnY4dEhsURp5EGs+cSrip02R
TgehQH5r79D0f8UMvUruT2R7Nag0pjaV8ZRm5kOgkJkVpHQq/jtjFGBbaFJ/KgxZsEgvnX5MukqR
Z/kmVbMebNmpRRisun6mcusr0/T658Cz5H8t5Q95zAXd20gyHbq3n2NSuWNNwznRdDDMDoFAnb5X
z/p5lMihg4xPskObGW1bwAsJ38zTT96kvXle5AjoniK+fpnCsCRavg2cbjjnNLzKbToIOjiNw9ev
4m3fDeI61JCeo1mYA9C46rPUJwpLIDZ6LudHMS6KVK+zIsPyHWW+MX0g4Pk4fjE2F0iC8pyTSU6y
2hyTDhqUeMOs0hSAUry+xquzcrBu1a/igIoyz+Aw9YDgtW62wZ+QlMwXGsrqD1jhinsxjlrfgu+V
zk3Yf1tFhmKcL756an6GieLm/Oj42+OWCTjtHKAhwkzRPBi2AOv33fvZ7N7dXIoFKitOVdotp5Zu
Q7WViEI7Oty3XdFxEGd+4SLp809jbTNbXAlHreRML823NKtk7daQR7gyQQaunBNicAqd3MaI06ls
NZx3i1HaliuBUzsr71DBbz2fguvqlAj9afjoLT+lXg5+xykVyZKMNzi+5JE3OLYMyL9mPsXBdPjo
kv3o9gRPwIj/OTFFVTVtCB7zb3mcEt7RBerq5lz+2Ve3Qe7YOCmA8s7ZPcuZkmaSAOlgM5bxIrl/
aIkEI//bKvdaGGpYxttDVzwUoKElrJ8Qtisuyqg/e+oNvRqAANwVhNoACqRcJtSNWMHWXoIGjpCt
YPUp2tblige0jE1Pt05jrlj/Y0MomeKD73PD4BBK7u5T3UpOHrnnJGkSFqKndO9DwR2cXrcIR2Pz
Euwtd7qOJ5reX0VWc4/dwxMKC3WFmkYdvBENXLFrVYTfPGnEwpv8OX3haDEAvkJ9ziWCfCfIA5FU
HpBvTJV1qVsQZTWQ9ZAqJG3pWUiWZAhVe8Va8yQ5d6yMIf6sutysj5iqFCYVQ9V32aBVb5eKTgu6
rOf0R9Xy/F7oPis8/com/0BmBlxWW7AWXQw8vU2nlcHpBVQXHriEwdh4Y4LDatEtv26tcNovKmSd
sVmGVLRFqxMB/d1F6NvrzqQlhe7IG3myMy8TDCuhyegHmEMEjX/19u/OQh7uxQUKM53dDrFg/aPk
s8qg1BQQJC7yIZ4Ez7pDPtb1s/HJCW6AXpUq6mac+0cdgj4BGjaUNUVD/X2Id3qB/T8IJ0bbli9h
NLO6g7myT68xOqerHbggnWylYiZQP4H2pUHf8gWW7RqCVH1FIk4sr6Qr9aOXuqP/AAfq9v302jfI
Y9yu6TrTkV2MvTY2XRtKJe6xzK1B1vv8cFZOiZ5H8kUbkBWnzdMi0LXkvpfL4RZKN4zbMv1cNn5D
ofo856MdG36uYWT7vYoHmXfvuqkBqEaQD/RAPJh3VR/kWaTa/PWVwELARPvJzXEvdurwc+bTXLdT
+c21ZTVvbpGyACU8tyG2Dcl1KQNxCuU+0k0YRYkPIY8kyA/roZi1dWjQy4pJXRgN6sAAOjJVCMa8
Gw44ExXhGSpO1KVTSXGJJWDGl5hfGF6bjuV5+cP+3QhyRvyiRtuXCEUZ0I7NJMouho/kGd31ANbq
ui6bgkUwnusfoMPMBjREV7QQ7IVKVl+xIhbwRWreTtndeF2BGJ6RUad/DkHtA2uaKV1D8XfGO4SD
jZQnOb/sF/9wuxDI1Uxwd8jz3El3XdcxbJ10UC+XNdMBeps7LTemNuFOYuyRNkImgeDg7dQDw19p
xg/NPLeaXS9qdzdT8DLZjo7Gru/XERAULLEDsvlJwLr4yneHSwji0a4c9iPzd6I0E2GL2nt8Wstf
Bg+AZOvzpg0fJrAnSLoee7cEF+E5cVggOuEyQDHaQbslX/zd8DXvhm0otb7b4QHno14JZdm+YwYH
h55kIcV73CGSTv4OCP0h9ABqPlRSWLmKKHWjirUTGVLzSfTpSHa5grY1EAs/o57qjY+VymDZgMmr
dqHZX3ePOsY09A1JgHLkABtFZ3aJjLMZvm+HrL8IUiqfH+zqLn91sGk37XOdNwLctZ98GIBRfAT/
sMned6d0XSx7xJBzivdbRjSdOxMdE4HE/7ioB/FH4tbhPzifREXRiXUYLetLjXnWpiZ8HIgri+in
+IlnYkeP+kAVldJYEe7W75M2vRmhzSKykbg1h/dMqbrCzxO8IE+lX1Kn9TsLkpMPJyVjGhPcxKsd
aerZXtED/+ExPWRGwAn2hhfb08mzFjdUHBT5AVktr8acM2iSeEUW9f86jdofNEGWC3BvtR4R1g7h
kSTBGwcaT5itA2U/HBD47PxYQRMD6G7CV0wII59tJse/o7KIc54Aa8DYBd/qolZ0UbCfYuhxQHyS
/jeiTmB5ZUxD+mCbqvqKTiJGglk1th/UE5KrtpRXChf0GpCqDNdEMMIQvnn+Us04V2Xo20CcEFOd
EGI4MpdisQJDt9DRs8RkyzGS739zsXFcJS3KH7OCcMRbKjbSWDSYeR4OThd66/2mRa+J2yiVNZec
aYtDmRv3swzCYAfkFsIG8XRhBlw4h8+xK43vC6K83+rW5dy76vGwQHd4Rqg+y0B4gSqpyR2O4kQ4
vjWBIRwC/+ZRTIe5WoKuoDAmsRZN1luRzZayt00UEtQlV3NdvefBk4fltIOepoE57buwi4b1H1hY
2jJzzkrdWbfiNICLcduWKPjbin+a4DDqm/LlJDfbJcsQJkfhfuaMXzeB3uADzaTn4FlqXcznwixe
Oqq5S+yLHNQsM49DU3iOUH/xcS9HNCtGg3zzCKtb0TnqF7CsuwuUItvFpXxKgC42sR1q/EtQePM1
ggU09AItaOGx58LuiyGe4von/IJy+G4EuXv3sT3YbW9LwumtyC8qB/cRgUfJlMT6SmhQayJpp1y1
nWdAakRAsPmvMr8ai6mmb13ORSICKPWOqQuHBRQkwqyaWHmWmwQHMwbqKRGU+uU+ZZUWeFtX6l4Z
SvCx+HhpK2D3leiH9B4/9T6NQUpKQxU7FI7CGkJSHWBi6rWOuzHhaXDskpNtl4xIGjkHi8bCIdoN
hfa0XgeRX8xqrK6hv5EXUQI6S08jMLo0ma+rCVpinrJP6c5QVcRKrsd8jC+7WiWN5dGpWuz3tSr6
n2KylVCd6BBKKkqCOXOsQ3OsbNOnOjus/GkBk2CBxsQ8czvmP78a0LWjF1vfYOs+WRijQzfBMPql
bxK6xavsltFVJmAoLZUrRCKq5iSBce/cwXdo9QMyBcOyfhnyRRoftJ5bj3SFHAFPNjRUR3oQ1asX
d20UCQJRwaWQba9Ggz7aAmkwDZo/Fkrhg5p3sT3IJqAJSGYd4oxfblt9ZxuUGFIM8pIdHeTpi4AI
nwfKljiYkfnktlGxpCS7CrPk7P5ub3yjLbHZcKO89IP0V723BiaQYFfeQHJ99juhnaJQHTwBF7Fm
H0kXxoGbYAmm1bAHaOBrtWuDUft/cycvHteW4V9ZT7YULA+vmFTHsibT9OGCl6kPgRRc2/KjTnp3
zx9onJCZrm1b+rb4/1JmjpsFGa5NGeyaocjcJFNDN4yrs8gzR8ELF6nSb5nHDeOAklJ4menpIN6Y
70Tp3rQ/gfRmV2RQgtd9XJmQcJz4SXygCV1lxmntzWMAqo7AVO+3L8z/gZIUcaEY1gITwEi04T7V
9o1u69Il9hIQLdIISMK682ecvzD8Jz4Bt/uFce9NwCgghzFqHdmISRpQVPGVamC2DQY4vBnIvnPU
zk2Ut4oOw1qVJY6hUNrFL6ytIj/GKXwbfqF4vSGlVkdW5AYytoj4rFtZ7Y0KcNXYVaIkCsZoW9kb
F5SCYs3CTkIcstLGL6jliG0uBKlsYuwIOTrIiTRq1CQT/PmBu5q+/Q3LTeqEZThF1JbsAp4xMVoz
nC+rtOgj0CbguT+nKC3sz8Ij7rdGFMS7JXox1W0rg1zOLzwrSV+bH48AW6i0OAT+O5tmgOEvPJZt
R/5AkMgbYyPWyao774zzJAJn7h4IRJsF+01ojAUac16KskQTiFduKE4FTe2DDJC6V5VtV4QKZPgW
58BPkQKaDQB0eWtrufBXQehrf0gEk4gfeu+22kN9PDgPoruzBsI0kuUkGbMOSVWoQyPvc78jU1Qp
e+JUVtDnb5s9HsnzXtIpyPLLWJiCoXLHOifficyWxbXjMs1ebc8e0BBbI/nSxZ7b/ODuub7Xd3Tm
+MX4q6Nq4UIOZHgCpzq/IwvFcdsFuaV0apV0VWx3T6GdJF1ceZf4hruQYWlhHr9AgXLh9yfALndZ
9JRi/tlOpIs9QWvaE4AtFz8ZQ1EQ+mZiGPpDK5VOMZgSWNU4IuY+tPd4IXOjpE0ghXQjnctuPdkF
7gzPlvKtIgBmfKIAMab8EVfQQ7gj8N/Hr0kQm4KRNQ/9kX5v/if/ySdR8X5MKiwJyf4/8ERePYig
BoSbTE+fqJIRxKEgOd+WzlCSdJ/BJMLE91IbnIJh2phN29SDcedMejuKTCerwrw7//lWTT7YGQSf
s9OQpbAoACiEuPCmIQMlYZ5jXzHR8fmICy1tKtgSa8spddHqnqe00YByd7RjIFe2jwwzu0T+k+7T
jV3jVyXZ/XHw1zBgqaAK3TELLqvTZKI5cxWVeJ12ImO1vmr7/OMpxhm2p0fZEpw3b8QepzixvJYk
oLtqYR9nLkohC5o23/D2+t2vUfWSoq1f1PiCDq+1sRsTtLPQY9lxSSXrTsStP4pAa7WThxeD7wmo
cjHYZHxk1C9Q4be/Mmsc9xd2AtNsHY5214Dru2e5F7NOIGLJweywNumLm/0eu0Vqs+3Pe1pXlAdO
oP2UK4hZn/FIFz0fGU04dD0bBB5okIQcCS5E6N0FOXNYVY2tU9J6z9DQc6dFREXISDzuN1Z0ugtI
8wltFou1Eb0jc9kG5/nIFPZ4Yqv66uP8KxBQW5pA6b5d3tapuWrgVsR0iDsKJs0m4+iCg373RGCg
yLMVmysIaDbzpJ2lq/1lZC+00LkTDQcTF3+T6njWL/m+ETF0X18lZEZnQuUCRUgIZ196ZE5Za2oN
/0itHdoREUIlVIcoI67QAjD6iVop+MWcCfsI42L2XKlarAcbM8xRIHUlfI1odQ188ABVgo3hoYHD
kDPysqS+K7WjZSlCXNJt7Pc9P5T6Fg7ZNsY+ICD1D9fPKOjtbIlFJqwg6y/08YJ5BkvNP3I0HYaI
OVvmg7G6Li2hAZFws9NTt8mew9AHX8WULYNazgy6Ul8XZJA4NFmGlx8Y51sGqaCMLidO6oRBbUwV
/dwYotkADDUUG6AVMyrDgQVbzv1fHK5wBxHTnCeD1/EGdOERLNTBhEr+8TQeoPq48ibHNYwnZP37
3bDtfrTt+9b6Cqn0IUvfWghfAo2dhFUcJElrowR483zqv1+eqFq/Mm5ZrOvTN6O0yzrXHbBFn+JB
x8KQg23pICvh16q0HKcui3oN/am6f+DkeH6Q6ejHANzHhbyCpMuGeAnzg2WNKH2C6k5fV383sYYI
I/WMI6ftf4v63YJeLau+t025HwJB0kljlNW8KiXEzL8QfAG3+7kOWuny3OmdE9+CKcZWVqC89bnG
PUbaIHI5l5UNFe83MRB55iaCBYXUpFvoaswVaz1jaZGfWx+wsUfH351GUtz99TkjXP7mbyNIXLo8
dR67lK2J8cLVdfJwGK2jTBOU5ozEdOU3Q50PEj51U0XFeBxfBKjudRxdOqtsSilEPLdHoc9KvSe/
sFeKWm76F7lJ/hlVsDHIAaEV6KUTaVotOhMc4y8Fw6LMz1bLzISjH8appn3mZP4iE6s6En0hAwSm
ExKTxjKX2foivdd5hrHrSp/1hMatvGkHqPS+0M5Ef6JeTEu9n/fqEB1GrEZE99je3kYMy9u1GaKH
RESdQYKYoor3Ymawvm0+583uTR5zUO6JsKTL2nYsWgBtUd0Z3OGWayTb9Ig+HM3yzh8ZU5meArj0
jxsEEiq8CItwUTq2h1hpOAvXmn68c9Fc3rc4VBI9iXM0HJMCtBGKjhZ010Un8H6jxVHFuPtUkeCR
uvMjFb27JBPM8+Q1dgJowkcG6PaPIB+4wEaHTPID3t/AdGzTWd7hO0sv/L+bDYe1hbbgwskBf3ge
Lf5Ebd6OhLvVoRnwYD2r0RTdBw91Lg5027aL4qLe9TmgP5WCUg/oX7GpnQ1deLjWgH2xzVfZYgsv
N3w7lWTprQV/mXH/xMAbgEfgE3xXQ2uDgndq75SJsXTpPNrRpvVoc3N6ptgJbMGslVmXwn7sT69q
ZvgHnJpawwUlZgllrT0MdCi/n2Ocs6uLZbYwt6CB6uPFk0dzLdwtpyDyIU2xkabK0E3+hFXOqCgh
jb+5NHVqk2kWXUn7JNBhuoOAxXp6aztDK4xTwQc3wVPIY59M23BAoA2q1ANJTwQ+tcNoBsUQPTth
oE60bgA2TOOGC6eV4gAnnAw9nXJEUDOtiNuK87+1Kk9THRQu9d8iOrRArdgyl/b5Sp3EIXDUyyDd
6tnSVeDixJ07wrsoN+bZlqC4n+FwiL7DsroSUoZzLKcs1Iymp4qTFeFqhhUkH+pd8Q8xH56Qbluu
t6yiyIrn2wnJDzxFFwoXjpETY/BYgK54f+LEFPfVlUS3Re033BXVSUn8iogHaGuUZvcpgKl6eTuN
qSXRbLaAG5j13uuhOhKEPPOCr0rKHSoDLx7AW4OoG9UK0AsnDxCUNBqjp5B2VliGaKPwFsbx4ORU
N4lB10C9PWNtAYBQlLJur2NkgYmxf3GQStSyFabamPPb1CoRyicLFNfhAZSzCtqTc3om6ilgFoI+
vmf3skiF2MhxUqZhsVDTKRs2KN93gokonc4bH+TSbv9QjB1/ZIAYa5LwxXYUPfxw9i4rmPbdhMT9
fVDTzbvjXmcphH3WxT3LimRX3oRcO3XHNMPSlqr1ibmbrrekA4oeoTSJJ338txBWesEWnd0tzfqO
RwqAnol78yFucylM03YojGWitiEv9HepFtdw6TmR9oO0Z3HWhu6wl5/ZF3zbKij/Vev4NQY9Fyvo
LZmVLgdiwUDaNqHZnfwkfGNbSksSHwHDS+Vr9RxyitLv8gEnAMwUqi2lMkn1cKWYW66y6MWVaPF4
smU3ppCviw2XypsrEI2ENOcxGeWKn2LtmZKL6JSTvqiGvZsGzEuXEjfcZ7qjYhdqM6Ig+QBn3sEB
2Q17RFkKxVoHNmChGePvt74ogHKTWSVyHEkwXPKLMQNCp0qthdl+Fis1FVjUKbnKFkQ2cP65VUex
ZhAV3ywX/4ooUXw1VCSI2+s58aGE5SJwWg03eUO99uBprnCRClh0ygNPl40LFrgeFGE9LS09Ud0x
9ZuGnBCuJZTnCQ9mud/h+9NmURyRLVYLJutrjZGiOu6ZNXgeMbqt0MIxOGldImFX6j205rdqg7Gu
WKMykP9JMAjzgtKprE6lFdrQYptYpd0U3/EzTkQXx09pNh7Fxev81LxKLMID4uLhOggvsZg87vn3
UKO8v17DmWJRkx3kTbifxc/hsZth6TYhiykGVAIwJbXlGhwOmvDAf8X0xduH3LUvvvbOnuGf4rW2
AxAPY+6EfhVvwKaJWhjBC4Fv6OS/WEcR9rlZFqIPZm8twxlBd3YuHLyZpV7d49IQusqpKH5bsjHE
wKAIl0PtB8kwDCFRzt/Z1f8DJ2j5LGM/Pqs7dO7VB39W0gYuG2pYPucNJsY0alSew0ib8fO29DvN
QZ752dAJTdII2r7BbddcLSOfV0qRZ5xTfo6K9qM+XJ1+1cbPuECVOLtwnWRRZCCeQ+IPF1kLmbP4
2GoyWMyTW5uI10vB3a7aQAWiMAD0EhwHKJape+NdZKQEjSjILUGOgOxcJe2GbmxYAIVieLisCWer
XZjBmJnsl80L+Dc1Hues7bphauXaRQd/Ip+cPpO760Nae4jn24DiNcKC8R/bZbKY2Tdu9Q2CClVH
zG2Z0kFo6fyGYJnCuk4/cSlB0Hzm88UOZ3HDts1Qk9v/VPwF0vunmt683MgXIuIjt6GyTqRn/9UP
MqBikJsJVyw5PCNCazWqn8gmsMK/JAR+RWFDBNbBjbymeX+NV5fljPdsiH42pqfyHyUoIcWpMltD
4J2dDr4PsXRUYmY4YrLk+s5kL2R1K9U26ztw6wDp2TML04ZZ4QUYtFdeOauhbTZSulEDv1rir9H8
WtCbqxugYnSLrG9Pi4TWAKRzPb4JQfv3Q0NWK1j4LeZVgJthC761uT/MfTIeSEr5MNTBKfK9cOF9
X2Xcshj4KEMPrqh+X57FOryXfbpKElj0yQH+nf2z+DdDFB0+RucmAw5MuI2w4kNrMukYEgNY23Gt
uiQabeHIBDOa4MP2gUrQOP9eClQ+pFweVdYtyZLdX+PBzdfhfCDSikEbbYfjJHsE/VEcrVOLk4sv
ij6Kxn94Yg7MOo4U/iI0coxdio5iuU0GS6cUsQnWK/8f9zq76Qkqg8cK7ZthtGtHhcB3ePRhP18r
DPdgBve+9RoopEiq42eJQW6iB1NjibexbKmj7EnXLFikoMS4xne7cj2hyk4/B/hdEnZqH2ev1gU6
pKU2YA3qKY/Q7VdNd8l9m0Q2xpfWqO4lUV7w83NioPk6vbKOgtEtdwEbUo76in6eseE8tQiXdLPE
sV4gwPL+kF2Rd2KsQH3QCUSabruuVqRgiOvanNYwEcCIosDpH9/nKniCln152u8wm6KftlLR/QGU
wIdcaTQcw1vyStQUwXs0/svZVDFSyu7VeC7+wqDUPPleGAyQKpafCndyn/He+axSBt5zy+J/6Glx
8xldf01L/hsZHFXXbvvsgdlVe137tad6EMW+hx0qYhsJWB8CqdGBmlvuEIl1lBWzDpTsZpBkhlzq
aKyVTyB2UWs2ZseYFm37c4l3WYwMF2DIXoYxPQSI6yUTPlWUhsbuzZP++I0bzgznngsrloDjCjCj
bLMfduuMbouSknPitlVeEOQ8IX8KV+qPUIwczOKGytF2qT++kYEMLGWxc3+4z0bnTF+oODjlaP1M
jkBLwyxlfKroCp8b4ZclEa9VrCcAhYtdHRWV7Rq+Cmvh+8YD/idfDFkq3/PlrI1WbupX3BmkuLKz
wbZwQMy5j9B+UsIiqyHuAbV58BOQe6DPVo/ucqrdPhXBc5fNbFJCqWWePNBOos6K1VaE0FxgZ6/R
FPntTL/cq0Nu6Ps6jwvJv5bUl3sPnQmXaYQyE80cEfIcGUPSx+6IB4l63o89L1eqeidoEj6nb1Di
YHlqKo/82rGSnbt3Zri4X0idscD+M3HFrmgXaTVp4QSKdqkXugbL8aYwHSuIncieIt0Ybeue+qap
MQf8MTot/HE3hvBT53FbBlfiTR4mMSvA1TPkpwBJQHDqp4GBXQLO7096//IVdf0pYghsC73eRckN
ZRMHCViPNNfDpC8KH3rTEpwez/X76YMTUEnnMK92ULxR+8fSzqz8R1xrpbtD3bVwBGVsU7D8gvrh
yiXgLAueV9Uoj7i0YOdvLzprUFGYoZXz3wxYcWtnePtHuhn1tLBVama3BxYbGVsZVRfg9pzTqC1N
U6yACFqT3s2fkaV48975+m/3m4rBxdSou5OHEg3snbQpJWWzTVv8VuOYJaP1tY4QhVR3OlhLu16W
RF1U5OAWPheGHyDc9r9GoWtrOh+RK76GYdpfrvpZGYLKDO8op6csjC8AQZatP9L0rz/AlJY/1XlF
CXwYDmFsVNys5gMLRM27zL9CkY3pbQGpqtq/IybC0AQYW7zBPSbQC7IrQz2uJHZNpDqNuvskNr/n
WT/5hwuXHHQF1gtrQbMbKArjPPxrkengDxkOSAr3gDQcqJv5Ls1C9iM02G/TScnOueq5yaM/b/C5
6sOqr7gFN8tMmutlgvT8J2AuPTwUgYZvBDkx0QRIowRIiCzm8HBwvPwrf6oSyYAceT7U1aqkx5YB
EGOQffn+76LxZY3VGml0xxXGOfVjf2uN3U+hvVDowoQno18SBVAoIcYpubQiCJMN8ZjIG0sc20Ab
Zs7r7UMPuzEU+BUe7dpNhTZqiYlNUi1ZcuJXFmV2iTPTWCiNCEm7X9UinROW4qod2JgqDoJoVHgH
j+MVEDO0jMf6VVxdJGX6N7AmrrW95xZ9BQj6p+uJ90pu4mTeisUVxuTBUoRr5mN0KJmQxVmjSazt
Y5Q3BjxUWfuizvvN1mQgQghmB+OgMg3bkyGN80omqh35jpP5E4FWc8SVOBsFd56cNfnEIIyU+3W+
Lrhmehb0xls7F6LW0at6ikG0eQBvJcnktWpz0TypeBVaPk9cQQ1WeMFtsdSFzHdD4Nt5VYoCpF9M
RZx7Y7XLO9WvftBEiwaNoaaAVt03pDRYg3l/ISUXoGrJUcG9tgsIXmGj1vgGxfEJRFWnSXpvL26t
per9QLTknYo3W7Mc5cQvtDI5Z4zi0j7NhyAQj2EY2ZDYKrwQZfm1pPbVguTaJJQhFuqYvzx60SGn
uRc+SfopopFCuBnRL9JrgziYsHp2vmRoqtskGOeXLPmh4vj/O6K/ruTC6jWWjC7MOfxS07+1M8SN
UawOZT5kV95k4ZKQ5zzqOURdNwJ0b0dX2htkUhVrtWkF+NjIy6Muro6T0lWJwiarfMXIGtdbq88O
36OaA/hwlDLg9B5TGq2MBXbOKhkSL+0WVF+Z9efVRnYtd3jPieiOjx7ORwM7q3IM9a6dB7/Pc/kh
kNxgE7+HR0upiZ9KruUjtfGNW6prdCjRTJMUqm0zbSzhlW3TyuIu4lt+x6J5UfH9FVCHwC7GrNAO
xcITQ71EoK/6x7/BhZJLtMGGAnprvSt2vSTSuJisTFqHwP3ACpGwfG0qJJsw3oziD6E+1Qp2Q/SU
62gdKn6oDnARzM8AEBt0EWiw8OLjxcRvFaKzPG8xAlGC4YypaLuEcKaGV972VOy5wRKJ2k0Cmk/c
R/5XWId0XzZ1cCc1UGU49yFpGXhYDBoqTR6yI/a5d9IysAjHjVCKq52MtZX+s7wzPotdYeEgHeJ1
spB6cS26w0i4YfoS/QT1EUXblQ3J3bdBmldLpRxzO4+VxTR7QHqE/Iw9RhrNyXnTw19ebWeEQW5p
xUFYfRQC6zQmK47Z5YPaTYOi1RBEfo0AhrZlHvKkKAHCGiOoFHgG60pYcsuoH57qvEv5kXQlSk9N
fYUfw1xwst5f1TJc1sCPI+JPshkUGIyuymJ9nm9kYSLUs2ITXgBABTPbjWQeR1u5Nuj0VY5/6r36
NSlchvsRqdj1IEbWPB/dAARoM7N8+/0UOE/RnsCUpZHZQGFhkSqL8XZywSJtNKuk4JMk47DRmXN+
fY68+cb+OGSkk9YXtTyQfeTzxTlBoqph7tAlU4XzsIz+cMdJhW7Wmo1sTeaIz8ruoKnoDhiB8o3a
7NkD/aeQwv8QbU5QtWNlNRhZU70nqPpgYiwkNzLCFrK5gQqdC6CRrzX/VTDcRdtVzmHAxt1PCu9i
ZiMSOsf7VJVSyH0nfNnXOLGXki+yr6S05svGobSz6X8wRrRrSADx7aGIF5Onu+I6BtvXnwwaqNvQ
7ofwCtgPD00QFS2GKC/St+thVbroWdfebzcKBLfcvgxX44GTu4fQIQAxQG+93+b3l44yeJtTJ8vq
j8Xr80UNl8jsPY6Pdkrz7W4SNHwjiUF0HA3KlZLPLNtmxun7CIpHiie7CfqE8/8JUP3wfhYfv1uV
BmUs7NW7IrSoKElsRUOJzY7A8CZSo+3esOpZg+sdPmF0YUvJOAL8r/h35J3RdU2qu5aJun+H1x7Q
BHkOkaqdYqyHvOQ0yRn4fYHFygghIDjDF6D59XtCZ2J5IiPEzCkfQR72/LZ8eMoNixjRE12IRZTo
w3rctkF3Be1TUYHwwP+P6Bi06yQD4U5NKVBpKRDIhxX/jGnFRXjNKIv3tiw5T9rJbyHMkaqsHuPY
1ffH8fGidqJo5IHvfCKU0bJjAm60RVnC9myiDZtHwc/GESb4j+88h/Di9zedbnqyq6nhhXUhMkEJ
ZbQoEAe4itC2M7FpPl7YVRyS+9FFvZgvEST5NVWKTz3V+IFDq86yNph6cjme9e2va7ajOlT+tCM2
8jVIKrI9FlK+HsR4UuIGj/7az4Pkpx43zce1Jw9u/ZlaVgbJzBQ6m9gMLoP/+yTQ/Ld4sstYeqdM
tg1XzkPx0KYXT8WyE5/pxzlk3fWMWaeTjooaDNmm39z9UDo05A/1rNSKmWGYJV7GsLyDXMFAyCho
N5Ed8UnXGLHHZYLwMQODTyTe6Vq+wyifPgjun5yHuNyDUpEhSvmWZHY+wlUCWzuneuN4I9SFoomU
leWv1eYRZ+WE1u6FpbTkO0m+1nRG2YIbb/JlYnHDK8qQpUeNvH1jAlmfqAAlywCac+zIgdMYs+ne
2mXEXeyhXYmSh/MYgfPjbF+uRN6F5rA0h/O6nnaqMp6SzSE+hfEgU0S3NzSAl+hTcZycUAWIkrIA
FFHdgbJ92oJbR1S8bEYG4OTXmMPbcEDD8H0imX1npT5+Ns7HcMRwtzdL7bW8gMub9TU2z0tUOZM5
gIse/YbKv/hMTnb2P3zkWYzEtBvLnAYdkK2w8Dqo9pirdbKEo3OCPpEBCwc642OP//OueqOqYd3P
FwpyOdfK9MGWWP+q/2Jp7W7WSDDG4ow4ArcbB0iunRdyTs8scGKn8XPpbGvkiJHQuju/Zy+c2ZHU
YUrRMdd5diiyOolpxCITI0yda1N69iHyqpqtolRi251yYgIkDNJSDwScx0zs0Cz3Uhdu+0VBfP54
DgGzKFORCDShzSP9F8SbxxGu9WkWyjzBKh89wMUSkWY0vUmGRubYDPGJUWhdx1cKezXdL/Ouf39W
C9XS/8isvJU9JbZ1EMBmHsP1g/H9LiZDB8umRro92saZdVMkPLRiV7xAS5ql6B6uAMWwxIWvlyNz
6rY8cVx141iQUfmBQbfWWRpm6lDBYcRC9wrBdIQleOdn/KzvPdcpLdyQ8xmuGDGuoLDRIlZ/EF6n
0+nNIoAozomLfCe9FJbnC6KL37pQOhl2db5Zc1+cxD4asUftPGlmOmyuyy0IsV3AQJypHvicCSl6
IEkgesDSX3MlkLsK3sFHMlRoARPllgGI/oOSAEVxvUDLHK9TZi0DRofaTLzy2QBWcvg+JFIbQkKn
JY3vlXIXDQrvZafQTzAzrKK9Vv2cOYt8dmQipbgVtZ7kPkGbGpQTUr+mXjySsSLMZpfmuMpr6wx4
TBfXdxBRHOscg45OH8XX90DwexZYTHE32Fkbwn4jb0vJ334HZGseBNgLhgW79/JBAAFRt2jZ3W3G
zoOU2RfeGhku5iUSaEPclH5XtdTDhSkaCQsJz11JGO3PfeePHaiNn+N6oVLUcTbBC4QIijoX40tt
pYa/ExXBMCt35yiIdxd/c2COA2hKJMZSfaRjwbxbkWe/fR5MNxmQ82kQxaMhqkw1DONi6sKatTtl
Q795xym0ASOT/fuGhUxxkWWftsYYNA5pOsPdqi4tq6ZvfJYJCXRD1zbg2tKQ5gJMELk5t/oyBaoR
ykEhAJGA/4JI+1m1LZ+Uz5rBXIzBNvgrbZ4AJfDp68I7ts3eI0cJjuoWBDWgJdyx0su6wEpLqCvH
zLnmrilxy2iviPjcvXUw+Sd9dcT1hhixOxqmIdFfkTOw5C/yy/SWTQ25vyUPuldemvN0kxqtvQDm
alEBO+cVhsh6UrcDqip/SmLAsOd/2m55NBIg/M7af608n+aE9bs6S4iTKKCyLy5sbPCwqzqJkzoZ
GjvggkcSaogOn0NUlKx/ytxgXa2u7PYi2tbkiDiwepWnO8b8KvEjX+dlWCUqDIWX5m5oEnIY3JaJ
b7dLac0Zos/pckvi7/mv+0VvD9Ls/KO/BoJQL+8yAQi8Rer0z/Y4cJaXYFHSMWXBTUaJ8IwgwiCI
G0/a8iSe4F39J6VqVadVLGHtvgOsBasCMdFyXVHnlEpUelV3I8yZ6lZ8C8zHYUUQufR5vnB9FTtF
bJTy7jqiS5DAJLUsMGNPTR00oyKjQJrSCpl+K1xzlOvhvb7ABA8B8PUswop1+hvmJpCskzlz/a/j
1pRhpqdJ9B3W6r8wDg/hVREhkQOnh5NlX/bNSVXoFYT2VRcL48cFH9xQdDbbDkIrpINQiLQdN6QK
IkWQngJjmEXY5XnJGtJpo2ORbtIM8SRyNG9SLvbRSlUj8M0KSHaEDlF3Su/bz/JCGqLOCorekQLI
zTs6DSkE0YP/t7PXtfWmFEge6rD2TUL6qMwNtHw3ncl33QSYFITAClCVn8ScUGw47QMO5CEJvNPb
7jSHZSPuxvBGqdVASOR765op4xTOSoQ2oGzP38ZCP7XNQk3pxG3z01M5a3Jyyrgi3rAWL84QVBp4
Th+oimSex4ciVLFnZ9F5M0yydikcef+Ax26WUAbwgLnP78YSg/A3vT376EZpeHSfU0tvyMWco7rr
piWsAsizHL/Hko5B98WfQtoLpATmwyxEVoFz/xu+VlZfMZZEzV4u0PkjQRaE3Biuy1V6bMDxzekv
7wb3n6P+aSn+dH+jDU8+n5xo8sEopBryi3xoaPMA79g8jd3vu+aCOu61KIH4wEtAZihdvj+PSDXb
sJbLmeNb7br7mLQ2FY5+DSjzKNiOG/EnOtPIAgmM3zN0Z7dKYPEvKRiTbB+pJ50UTkJVZza5/huL
z9tb9hXjBHyhYy2YuxEoDFkS6xoVzM7mafMFsyxkPirWMSm5i9l9PJWMOCvHIXZ5OLLf7MjFyBaW
5G24ohNnp9HCFx658CRIrXtMNfc0AoRwDwGwFk1xV1r0k+PcqFzM+eWvjWWZiIajp09KqWEjWgYH
rzsnB1aMLHXOR6v64YU8H67yjhaEqcFMGKvAfUY7qUdDJFUAKirTuGGhRKlLwp3HvcdVhs9c3oqi
YTkdUKDO5sLxGWSMs/SwD0ixnSRMHINI5pR1GtOBdUmj78fRN65jDS6vf21wycmejuvj7iOV+DZ2
QO8YgWChwXg0YgoOMcYHhYD4RYGV5fGNNK2tuMg5sesj4i15Tr9ed8BjBXiahJC28Jb2Www6r1Lb
uTdlXBS9ugtgF+iCWLZMgH89ODJrCS5E9RnYacsuznK1akU7ORgW5t2oMJt6CUCiHYdVKgFNPqHH
Wdy2HqrSIo48jRasu719c4Re2jkG2vFs/4ucOFgfVqiG0ZstvZAP25TIvvzy/ye1lPPr1nHdXrUF
WL984koT9NLuIdTeFM5P7RjWAhXhWprfqUP5tdEWIXB8fHE/5ijjG67AbX9TDyatULO4PgBnD0Zw
h/Ju2WaH1XQT5hLHoJ1iyK7Ds5IFN7EWeUd7HEsz6mVF8gcFFQuIaLgkG/bZMQeKdChsjtSviJEr
qD79eS8ySS/SIwH+21g9NwONP8jy0mXWxOt/hLG2ceBIlEa81Zrchj2hp+bQFrh0SgcyUHqcXHdw
ZSAeF1nSdjNJ1/l8e1SdEniyGBZDzbACDt0n7jRWdfwu5YY6ziNZq6Tv5EXNW7Atv90oocI9jX1G
Vc159B80p5+RfRMTsNAw67vTyoERP68KbWzXn4X2SWXCsyHLEFv9t4Ic7HDiNXjQmg9IZy2BQ/7x
sbxyohsxEFPivxNNJjmi4dKWm/LZ1OY5GdE3H3j9nbsbIBRIMdDTDfts2wdJAh05Rlk7wkE/VEkA
2Z1swWNQg4aUN3T1419HSTwF1ZicqBtQO7XN6C2isO3sykzhLtqt4d0f35Xho2IDLNL0oIvGl9jq
1Kd9mo39HgIkdhFFlAnWEfPrOP17fTSj3l8tUWVm3yRun8pw7FX5sDyk19IH/eqaXScV+wFIevqT
o+ckjYK6jd+8e6ir2rwbDWvt2IdSuNavA3Pm+RczLwIOO71TNFBZECNrtvG62ty2ulAsik86HKE8
CiPxUwp1tpgNN+HUyaukdUDoKa3KadSFdGcLndDAK4BztDp5s2ee4XYRbQaRQ2csQEHoTLil4I81
zASRHywfk7+4/CIvXGHqQ6Xk7/2QRw+0/6ZY2JWRp8iPALB9NvGtGe6T8xs40/NUykbKZGvYIB1J
QeKg0T5O1n/JXDZYe8MBlALMCV3hz5wuZuRYQZp93ULvC3arOQUypirqfJN2PZ2yEaSBeSXIEUTm
pSoMW/9sJccY2XNtt2YZNeq6ZB+NdWQBxQXF0wc5zLyuVkeP0JCpmDro8OF2zi+ejBH+l4cp67p1
3hHNQ6SR4iJ3ju2GA3cz2s+AAva6kfz5h8UqgDzrHsu55Dit4sEtRlM1HPJtKJKGh9f3T85U9lae
sOZ8Tw1SPDi4tQpkevXMFt8Z9UXOtjcKAD/HBCBHYrG4irDmkP+h2Pm/tGW8nD+WOd1XGallTYTh
5bDyP9KZTfTGSFANoU/yuatZuV6fVgE6jhBXNVfny4lym4G7Mk+22bs1jpTCqgTFT4pjvI4P1NeS
YUvAgNVv1PdTixUvE4IrRy4U33bNDRHI6oJ9JZpEl53njOrwsThCMkwyaVURHSIKBrzQygwjnqwq
hzitf+kVvxRaG6nyuxFFhv2nikwC9UB/ZlvYjixX5mOVgZQ8p3Ud74Rw/ywNrfa/VQfFCY4Sx3vb
QTwWtVpdJ6nXCzUxD914rsxNDOQCVmrm6SvA29CAsVht7FCJRYCr2KworTLSB28fH0wfQu+irix1
786pIBMtOQjWF6RM2YEi7DX4eccZ+vhn+iY6uw1hAi/xMvSttKIf2W9EpH7h2RlH9ftE+S+fXi+Y
FDjiGUvuB6EZvTiihxVpJaKDNNa4Fcucv/dHYpOF0wls01Bt7m6KdaiN9JlonpC86tmBbUU4v6cw
Jw4J5KWPS4ClzMKshgp00MHyC/7eKpOVoo++TVLq2w9evFoioCKIyHZwidXKqrnYCXfPMhIgohtw
+re9n/rxDR/1yAE+wFbLPLfZ/LnQk0HsPv0DVAYKk59M/vVnbBYetd5eZSl5pVpOt/jyiMGBLBCb
WUbDvcSk2VuvHAVldkZ/S58JaHcYdT4IsvZsWmcbWmzrZapJTBNQaNjmP1+3sFdSs0ToAXpdzJB5
hliTEUmVqUtDbxB6YyJJDRCs7uFOaooOs0Gzzxx/L+rMqvr3WWbaGo+WrOgfJpJNW7QIWhMp5Zk8
+tg9GHYauLJZOPbjR9hlcJqoF4bPNCHHWVUkBmL81h6n3ZfgYnNjAdAOIQ3c0ry2PR+qyvLMoeM4
DlWexjGUqr421klPsWiNXmhVKMw+XBIkKhELsGHH3R3NhdCnMOH5ypm6necM8ORXGzOdQmuAQaVo
3qX9Aqp2N2jZwGV1OxVgKzVILl+9ZgJWh+8Eugfl6Rdiovrc9Ee4EoNyh5p8Y0kOuIU/ynjiBOEe
azxjKe9t94wwwnRkqLbIFX54BUZ+7yIez8kaW9A9y+8JZ5vxK2CYk4ukKtd6a1HRxqKO6BYnIrCY
qo+n6gnqfNLffx3Rtou3DogYoysQ1LgAr3NGzKPrVRf2KDoy7oCufehvv9hvazhZvAvz77flWzoE
l1U8WQDgof8kkM1g10J9j62W5f1p8gW045/2PoRE8Kz9jgU5zqDQxVV90yZDf3EDcnt4ypp7d9lM
OPYCNiAEiMaQCCM9MHpcYYYKhER7QTr/7q0b3VRRczPxNik7p92xYDgaJYYFpVa73GFe4tZeD+z8
w/Q8CnwE8LkUAV4sF+I6JLtiye1hc8blUfCTLrvVtCzeSRfnvQ9VwcJYmcQnY16/OsCog7FGixNh
oOVQSXTZw5y13J/pPR3meKBd3sVfS/FjBg0fXL0Szz0AcAyzzCyKi2nVFPAJ3idP9jLF4EDmz/BI
dH7VMX97YMpzLQfgcXyXJNL9tN7/bPeDvFmlgKXdZeR1AWxJsKF7mwORYAZqqb1pE5qVssrhRrni
IuQD9O/yfNIwtJAmz8wuDbjgCdUyTSCGEqfvUAg34bXGc787kijbQu9xwfPD5wPkcNXke8nWzLwu
TsILjQdXWQQDKFdFDI0pgu9LeJNS1kUAqU7vJRUPT9cCiW2E1IPujVIO36vMZYbI4QrKTbAUV7cX
j5fL/nCRoCNJNxNKngdv1DoxvDZ79q7OR0QkaOpWzKD1llEBFb3loEIyxm5jyMbeZIr8ROAMVKhs
lfcJh0Q+lLpnoxfuDYVSWw8z3pxd5AX5JlqR5SnluKeutteP5waM/iB96Y/4wIgbhSTvsvDPvXyZ
Y9YLH4nkkawPH3qlCVaELVYA+jkgoqGuWt1JAm3djCvr0ACH16oK5Jr0/lsJ+fNt4qzkukSRNSFV
p3YqKhRWnqMD2DQUOQcwTfyGZJtc0Z5stVaoAUqBbeqMkSZSYiZnBbeOYg1U2GMFD1uRuU960LFH
U84akjBQB1+6u+vltpCePIs1IX1CtZsJovI09ry4J6ovrLqHEZWODXeqiVdbk3p8cWrR3ziPJ1Gq
c4KZIHORT+bYw1DMdcPhV2s6hP9jj1vRRnZs0v7mCdw0p9YSJar6VLyz6Va/q7dbrQCKGLorwNur
FSLWUa0XT7Czs+80YRHCDVv3eTr/RrFJs8gO0XgPo5CKlQjrJzftsbvPCjQ32g39BTlQHssyo+tm
VUw4Vn53QfpNpfcPItbOuzMfClAF72mbIKucywd8mQdVGFMxbQBkbFZSsOZ6pTl8xr/eItYSTLCX
mYnaX6ywb4zRG/JrMXKTELgUY+IeVGCdQG2dUbAiRsS+7bzhymniPKjd5olXQPI7C6GHcgmFscI1
lTDTOSciYzCzrzF8fzNbwFE9Ph/k52NXfzPWb5av+wHM6zzr5YfUl9SxJgNmuUirHzph2M2DdaTN
/dudumHZ5BTEd+Gc39zv9ojQ0ETGQJFDetIDePgwXK6ak8YxHHfvC03/MWcaJ20j9GiRilHEFAvH
HBMsBsDS0gNOIBD3d+/nD0z/A/qrmD0OCjZgCBDsi0P+clGx37+RGvzGVu5XJtrcS709mrl07m8d
h/ZTZlVzySMZzKLA1L/mLIMSZHCPzry5aRPAXtXOhQ0ivR1oO9HSuVdAMdNveOx5EPCmD/yMjUEb
NAGYb+X4/+5WmxRmOZ/hESOMnDpT0Xzeq2YvEN2CqDQhC/hx5JxaAwcfE/nBrbpITIujb7XM8Xti
dlZfZg26ON2DoeM4jrYKTo88M41YZVsemTItv0D3KF0MVAAEDw+ZjINPmkht4TSB8WcksUAdx8Oo
O/U1SHqs22+2sCpYFbRmEy2NNZbtI30VSzAi8Sh+PVArRhsCFITkn42vqIktByLa7z5XujXquoB6
+kCY476AckZY+lPs10sqv+EDrdRw9/xKcb17uFo+oage5c/NLUzeaL7l7ijEgldvHYxFYdOkSC32
0EmH6Ysy6OIDUnseUqzggBdJ3iuzgh5X5HI+BSXklMVAFWh1stbUHZQ51HZ4qEiZgtiPFeOOqhQh
XHC6pYUb7J8fz1Sse5IQVsSGZEvBwMyjuVu3JWq+W263Sc+BALsmlbECIbwQXVSp4JymBIEDlQKh
tvmnnHESUoBmuGNW7O9WFJz5TSpFj3tk0FPiKhxnQ9/gEDk7mjppPsQgkcwPmFjTEVl430PSShk4
upjSiH7UaFzYbsReQLhDul43K11cPAG/jtN0IcyFBYqUV/taN0y7HJiAsGDBaRgUl5N779/Ii6Uo
DfleJzDyD1kNCHRI4/m5zK2FbLwByd++lAn60I1DHK0xJR6piTdF6YerTflN60NYmnXMIbBa3SE1
DGuWraXHmHNO5HfkLkOypl4u+zS1mBgr87qZAbIiDFjqHNsOyPkHBxYKnCURVrkoeJzSpmrdF1JW
HKklzGO5i/+kuJbBorL16F9CHiNQuCW1dg1/8cxSuaM5utFanVGRmhDRhYFb9894/bDUP6N95F/6
5o3eRgQ6h7AHm43PzFuqdU19rdnEVQsKfMn2yB+MjYh21CVwZH8H/BvFa0DjVPGkPaXS0UYpkLAn
N/imOyK7VwJfFT+dPjjPQMcTSzP/M/A1ExRj8jdgjtSod0WuQMxmQK4Fw1jGIiyEMijrs+jPvfNa
uk95WUhRiD2pKLOtzvY1z3UdDGKfyCf3gmO31gNr6G/l2cetU1xs48UOuu5fL0pF1zoK5TIonqjg
0TfBNL3OFRax8UbXLOABdgYmDltg0rIuKVrQFr5tXrAgihXhVJjvk37aO5DZRNIdVBAYoXl+wc31
CMNdmDNkPL3uyWzrLncK2x50/UFDe91oXl6A/EOt13VO+YdeJn8rwYU+Xcw70EzCWDsbeoI0r7gd
OTTrZjmzkBaFkwkrLK3PBCCQ2mHrFnntM8oH4AboOfuMX8t8ffLHclmKXB7Fv13bzkoo8DBnesYK
vTJlq0Qis1IlWhmZvgYp6xPqaCrAhLkDMbvvaP/sLnZFw8a4p86mD4OfCYpgEe/apCpP3EzjhdoF
WAlyRBRnPQ3eXT1RNkglWaTA5aqbiwYlohodKWzbh46JBVIZ/Oara2Ix6ZRPuB0a0Le4UA5ZR3kv
RvjvFRACxIKeUm+cqXOC1tZqpeaJ1/psGxF2HrJEHM70fglhVXsok5zg3f1P1iu931zPb3W19TxQ
ANqI8PTxpY6uB9+pCIcwRkv61vZgLoJ2pe6K/cczP1RQwlXUiXHgX5fF8gcZ3irviLFpdCdZH8NK
mChe2/S4KApD7A8Y5tUAhpVEhXL0WZS/JcAYGLmB/vmgLcFF/32/ibHNumqjAm4fn1AIrs1RbGIq
czuUs034y4e5nYmB0Ab9bz4lL6I2AdIgqWC+mj+ZGslh+3lcrn1AgKml3bLlYY0ftRH1AroLINnB
cuksprQLysT+RNcGR/7aiHm32jGF3MAGJAAPXFLXgONw5AdTS38dbH2B7xxtsh+WsjdneuMsXoPE
+bpfImf9gZBZekt0/Haq+1nTUJZogsWJhzKJMfZWeqf0dHNdkzTSb1lKq3L35tIxUh7rEil1EqPJ
l4bUe0I52qxueE/P8CCPpfrcnkuqdWEA8+kvwrOiSaGY5CMwxRkemHp2GtceSTLNyw/QO4a+RPTU
5j9bqjwlbCvl4ulofKFnouaR6OAmo+Nigcz+xV5J7lJREot3Efnzgz9pbAgloSrQr3kVai32CNXw
GnxznDSWTF/Icw0kjajFJBicFG1zRMB7qXhO5niXvJ1sUibUJg9+JxwxbK4XcCBxqSomiSHgk2cl
PrMq/cM4R0uCxA3A4BQw8r1SpxGgFduqz3c6Qo2Fc5IQIStsslCPlKqStRCtschUibGldxbrRM1C
jaQstFk1TqkgLXxKIe1WaWEE8LeWLszu4qU12XGO/yd+bf5TWWzYjkYmpIJCcPfKUyeMk76LPE/N
s6aGKrrjLNOsAtk6qypENfWCBYoKIi1HyCIBxcMQCxTsnP1dJTf9YSKHO4KnDSmOryFf3N1aXyVo
6qJe1m4ccCnIRMdK6Cvq9tRecvkCTwageeAdt9uuzBalZEQexTQFkfl6RJd06RGezkRSpq1r8VGk
6Ix5l6egBTgk9gc8EFoy1TwN/xwXZXX7ZrsWT3hRXCwJpUkYZ5Dz8hkTexKk3tmbJCK10+JUTUD0
54ceReaoKqtDRLCCs3C5TDTn3BWRNZSYYA8w9Tx9+hfxKCpStehSt02JrypxYO94dt0LS7XmvfFR
N6umzDwAtVDpIFfWgZCtTF9fBXesDwQLUxcxQeYo4tTlLfSgbCN0eehWrYGJ+4HI/TbSwmcM5Izs
5IZr7mRG3yBBea8Q8BHVkeCo2ZkbwlrdPdtrpOrFKUjGM+9Hdr/Zt/MARP1jsAqvIZLSl/keOfgL
3cusGh1Du4CIhN1SU8QzYxDyccN0A6N7eZXVugRjwLfimnI4dR8tGJVLNGJx9drUZykyIfvCV6Sc
2ykUJPL+f0B2nJkl8k3oqmEudnir+ZuT2BtGoH+UmEgzKzx6KxSRm/Ik1+avpggEsQYz5R4vZFbq
k9RCtpKYQOxfqNd/oxMx5jM4sGOufS1ZR1W6c6GGunr5sTRG3H4hx5BHlMrL2zOPihEUmDIdxWt2
qU/2SwH5kIRoRq8hj79GZXMCDFII7tNnc9hTho3rAyZPpWdTnViT4xOiV9QQ43IQUmq4R7xiRvPR
o7wIBSbMVEVzRhndOcP6iAhN28KKqjdsUFa9Nj8VWqNv7ynzVsPe5k1yDY71g39ybqGEgCDtzRfH
iMdMc7OP794a1D/2wTUvjj30N/vyOV7hAqvE0wu/SmjMZKC8OC5jGlFqr20L/5f4oLFmUMude7I2
yCvrTfWDwTdezkjtH6g7bZ39ILHqOHI6bgvVreh1mpesLNBiBb8sLtAf6QrPjiaeuul/kD8TyhAH
e5MkkmAlyuZXRCg3buLpbLUDBKl+DB9BpovmMrV8VKSeNIIQV9fLhAJMzGPWCzGvVshIMEsgDTan
FQ9qovXWAACvPNnUm7JrQORfcIdzditQ/JaEmEFbldsdWo9Y4u9Z2cyV+ijLUqH+bFOnfYozksd4
6kPjNPQXR7KFefworKWsHwkh9KvPmWhJOP8wQwXmfEs4MyFEq1ssy9vhop54/W+BC/vkDv6Bd3Xm
WkYyKJhXEgkg2FjRzWWlWtqR2nEH6rS1giCkxAVmJQDRt56Lxq+q4WIMxK+dKf5/IQ6VqL5zacc4
TM9aNwNcVfaX7polfJphbBXASEG8cYIQU1lmffVGI06kzVaWJh5MWVpS89Fv+XUlV1aspTIkg0b4
2HyFThrSRQu5QAi0K2+S6tTtfxi8eCpqW4fzaIBPfxHMDHC/MSuzlokywBGIJrZp/pYrIHZAyLH2
lDg9vL7W1GTKBBWpokN4HrsKxoFtjpiG+w4NVpHd9ZGys9+W9MPXgt2hLq0dsY/FMoPlzh/flm1K
J1UE8yisNLYTnRP0OmxwW/e3rv4N5wPdP/nHpq9RX97pC4SBlusijOgGsd8NlSF+3YeMwedcBtNl
2pyFd0/CEZuYaZiv8NODc4OPAObPiak4g1Xqe1x3KjUB5PrRjLnbsM8ZUyij5WElfaquQOStiCOb
pUauCoayXMn/aCpSLBGVl1NdLVHa21/EYtKk5ICrdl4Nn35Dy1v1pbq2Z2wrV32/v2s5pojOf6Nn
4yzol3PrWKb9Yfs4Z2OHMEx5+IvExh9rq0+MBe5RfynTuQuNgvkUcf2z3tEnMIJW+vI/B9koHNrv
HsoreTWrmsUBRZxHBiKjK+y1ShtgCa1t14dgpcahiEMFijdJHxoNxInHIluiDLPY5WeN+NzLw/n2
7PIFWMJ4H8Wzbe9TWw9iggu0iErqWq0pMv4YpMhsPbCqIb1HLAr0JDP70wMgw6P+YqKvV8mSCIj4
QUcRLbWGjQEeYEpg9ZmeKaEKcJzuakRP8qU0wGudY2VUgMbYYnhE3vduKRagGxSPScX94laH6Lnl
oSOro97lzfHxzeW5J8/pVg1IgQNNB843eP4S0kOEFe3Ks9PhTO8RQv4RCh1Gn/1ML4+DdAy/seDc
8K8UlA2AN7io1ySACe/qHHXI0qVtk2IHvb2h7GKiSuD9BnsC6MKi98Rk2KDCM2KA0dAKUAvOcqsF
PJoIqsUUovGtHLdfyazx6L8iyuprI42l3NLP7l52HReu7UnTZKwXQf2IfGavqr/qclNCxGxtQZUC
GBf1ac7wPDckb/JMrzBctPm0roshk6wSjPCLF+VehItDxUisUh44radij0c9sgYlFtbmmQJXcKpg
/ZWJJ54RlllcJzibGbyqmmhS9N/JFxA9J8hYdqF7ktzbAATTVqwyU9G3Tl1LD9qI3fsu+HZnauvZ
2XfxpNznAIqBHroBu6SE42t4uvv8OQwY8YVLTpTPm6/TR8LsN3vwc1ajadkN05HRUJWSd8ePJb7t
/iNMhWMYSrgAlDOvSbEd/2rsmHZGT0xw4Z92wTmpLCsB2dhCzYjtNJObLTVYLWjZvsyisotgaiIV
mH0SXag6hOI/6ICK3EIdxFtGK/WcCbp/+qMg9Gwqv/ei4f0vUOEILrNKJnImmeBPUm8PrdGwCtYP
DxGE6J/Cmfr2Jm80VlpRnB+RD/TtB2sLv5jmPh/clEKtI9MK51Fpg0Zqyb4DMbZiY4ae5ysR4LBp
6SsyLtUjeJMHL3fwRQ+A6dy8BhkCEeSwErv1YSe1b8dnUfbFNs2ZeSS3fFARCX8el45R94utJhp3
HsckohCDJct2oApWNLB23No6m+XbJOwLsCuhCyg8qtUeUQV1B0zi/eXJ6IM+mCTXkijf9c1F7O1s
k64dA61jV8UyzPqgh+UqF/EqE7PlPgxKGd6Gaz7lAlSrJrIbBaduruNn3u1fsik7vhkrGB+Qy1kf
yzgTE6QaENxbix3X3L5p+hZj9YcXp1mJcMPlAaxeb5sskypWDt+jhitdfguqoMb5AO1oh6l2xPNn
UFLOfGnYOQGAk8dr0OVjc1OkrS3eJvE/XbHumSASaf9ikozRA2ACPhkhkMa0ftPxQv0mgiu4Uv2a
K8ah0syppTin9MXU9Y1Y/moMbCtYmQIEHsczF5SNfMzlgoA5nfZFwFB0RNImn3J78TjB4eEkEIbC
KcTpcTiEHR93mD7bKv1NJ8oGswnLqMu51J17k+VR4xID13uevHMDJwy07GbMbeYQWm6Tc0rXt9Mf
wWPUT5T3z7AIt4611GKft88TvXMuD+z6HcKXlflP5YkAMeJ3SlvRzdbg2WkVpFmfRkKQ8J99sY1y
5ikox7r/nUeFXdW2sTvfp/ysgQwQe/yoO04lq5xOMAdJt9pIYMyi+jMuKQMuyj36wYWQfwh+ysBx
uSqjgBgX975lYeihgPMXe0p7fKHevmMe5FuoRJLBpGKrbvtT6Vp1fW3/VY9NQjkvps63k5haltij
JMzkaR+awhaNZDxJakUdYzxprzFhIalHNLlc7TatKfZcLQVFeh0H2BrxRqjj7lPInlGb+BxXNHNx
qxG0ZlYVle0W59kJWyUnAasv3hu1Jv6Q7QMj0aJuePu5LGY9XZjrW8wESdR38RGaH6W7lk9yYNTU
KvNFrK/+QvO46reQfuk2VOFRNWQeLlhaZF0DADVGJ3G7Ky+lUZN+K3hyGqmnL0jtO5b8d8GkuJPy
k3x7KmUMFCKX0x+6MD7dKrNWg2pYznh7onMHdRl852KQNpYeItHeCZb8WF4VdNLEbAe+vOTDaROK
15uB9mG/VGpUdhDPnjxzWtRDE+odGawiV2OPeIZ3NN0hBcnLcAiqhvbPoYbUtAq30J+ZaPGxk/xG
Y8nBTQE5kKfbcj18NccdqBxZ9NAtr3kE/ah9TB49dbGqI0A3KFCNJt4oHheFFQqqS0mkVvVY+q5P
aYk/BS0ZT5Bu4n5N+ocSA05/0F321VhKQX2HFZvAjAPCLK0FNYFvHYjTKjYAh9blUToyQwqDKqSi
aR6z5fMZj/A2F+x80zufyKAAcAF0QRiKMEDtvI1WTuzmI058cnq6FOGu3kbJztFTPvLyHsX50NSS
Dxr4DlFj6FKqRvPoF6ZlxPO0Ss7gUUU63CvkmiKwIPuOrKywdewTstSvmb7AbACGRQ1KuZ10yVZC
5sE7sc5ncZTdDx5KNgrlQzAhk+ZiOfumUYiAUKLKD3d9EemMRMWqUozt3pI4mF1ixII0dJwdA04J
ooOUx3/LGSLYLJqoFjU5mjaScIvAKat1KEAKLFKbqZ0CuKPapWATRVjU2f6AYOMZBJvm3xTg4xz5
UzGMso5I0Du3v8g0ptN697KlHlKMSjLsCpaa77eotNA2QPFj9Vwc7Ow8NeujuvZEJX/Lh5bkU8US
5UeCxX78GbHzqP0xqDp47mSECIEGn2f3zM4sp3vDxwEfBLc6UyV0Fly2Mty5aiGF7ogZUqmAqAh6
awsUgXgoFtMRBpV1tvQD7Va5aeVV/bj15f4cS86gH6UcQ20Pt+1wUKhgWcsbLZvwlM8kJNnqwczB
LfGMq8bPq9/TvYA3PcXtiVRa4T5VuFpBHXpDt5hqfeEasnHdknDQIsfPAm/oDOY5ssOyfyS862SM
mBA4KemdSrvYifUocrCrDLM1p6dOLiitDfxFnv5qlOwI+ayNKw//Fhe49h+mudxen+z9zVudxSJ7
18Y9VM40ulf6BHGSaWfCc20SKsXZTgCpXtxwUJ0dyOWHEP52ZtGz8z1HWib25XZ/bdSwBNLWHVZ4
bjOqunmCQDXFLE3cTQm2DEaf9wKPBBEUeJfDmX7Tu0jSL6Hgu2nyHJxTsboezMNfb4tPzIHSA6l7
uEmHNVsZXkvmlo539KfSfgqy3gY/tHisLA2sB0aQvetEwmztEMq/6N9OgsBoxcf7mkw1vNvFgI13
0X72B7smyiUq9a85Oaz5jaQoYfV/52rXB+Gs1dapO2sZO1zNs6HIRprDSNCYZlW/DNDxbiLzmtut
YA7lVPFxVuQAIri7n5xzlfTCm9LPEQdHG85CQFriWlLkz0AqJ7caI+WL4WcGgg00FrxDDgN1mth7
FLmWZc24nSNMBWLmJx5MOS7WJGzs6q+RjXzs08wr5+APq9zuAMAI6qOnO52QOGf8nTpwdo2jBCZ9
114AJp9QE5NbU4zrtknlBEntFoM/zafcg2BnsgBcoiiM2eSJ6/ggyOx0XNhcsoNn28QPI2J9WAyJ
PeVrjYXaVvQtR/mScCmgIZto4jS5wirKXRrHDqN6fWEdvVMvWlusj0Q1N0P/k4lIjgBOlQZkCNin
bYMkKpX2ZDWc49a596aELNMfgwXBCyYE8Gq4gzJ4aJ0O2VwOXXNcaXEIB7DWH/qf1sluNAxiIBpP
iLLlmOOu+aHLoi64JgPasQo70GDk1a2Z2yXlCA/JgLsAWPirCRbK05VW1XGVOmIl3bRODFt5+rTK
oY2eGzJ47LupGEsSewb9pienV6YCkBwaMe6VORpK0p5lpz55r29lTbhValNOuoYy6aNZVzXrsHsF
/YXzq+Zz45gPD26A7HqYmL9Ugwt6x+tvZ14sPtWet2rTSvdqWwXQAkDqxTCBQdsUgnNmEvtfGrFV
ObHKyAJcDBmEQxHEyVJM/PNncoRfiqdNCxvtzDCDXh6bif5Rh7hZexEr7T4gQia2dfHGyDEAxSuq
9b/brpzEhFrZT/AGG+RvZnrF++Ck8uKeeMnUYtV1bRfILxE8x0z1AdMAtMjyZnT2Z/Ms3BF13LAs
8rjQH5KAPyyLe+XLtcDQVDGn0izyzxtvQ/2EMJJt03PPEg+cQkanl5CwUG4BwsxQvgr3e/qMd2IT
28pnfFxKH2yZXEOAcGShxO/WjE+oYgXLiywi4NuTTtR9dXBzs+M8irlP1M62kwYEV1m5j1vChbHY
gdAuzPgto2q1TGoqoBDSLrf4dvGx2Upk7VeLw0lgCsvzxq5IPLSbEuBQkEYT3ewPZ/XeEEQjy21c
D17BoDD94qIV+vFMsUDQ8/+B1sv4YpZQ6An2KxBtqbbh6i7CSV86AAYrCRteE1vdfUDGqE4FhomN
fyx4EB7ZZ0TRcEnYlyfry0PWUom8jZks+9eaxD4braRW0Yi5qs8m9WCJH7/4VPuKCODbL8EF2xmT
ZDpnLl/UJwy8yn2CUY/FjAufR2fwdHiAa5bwmGXZPTZf9PM7SsJ5KA3SB9GcwbL0hzdEUWWKQt/l
Oo1qjvWTKR25XJAu9QxkQCrZRSyz0IcDwDJPm2HvNwyZTlpj4SClm2zwSVXVNyD1NUI2ESK/kTu0
gwFZyhicSbgOVj4T3ODEv2Pj0M6BTAvhs6kgnNj1mVfnNIWpcmE5W7EB+F/XEx03xM0qhqogFPo6
czSIu9B3h6T3NALCN8Gz9aKUMesjIyEFwS/no0I1l+qorXufo1gUc1PgexhH4etva3I9ZNk1ISRh
abJpjRo15c7zhLQsPhZso2i9ue04KXywzTcI/2+YUYNXoCyoizmtXK2AgYMVsU1GK8r8568ZP/kY
yJFOTC+kx6PR5G6A8ZeU9ogsDMvY4RlfpkPs2GwetRFwenYjfXWc+qEyJd4lgIJkhi8ABbwFXfaj
K1mpldB4zgJEd3+M1oYmp5mZwlJF1OHrIQl/jIserHiytjg4jRszOrD5QLVT2v6D+VPCML/JIkV/
86f8IAQOmsRADz7qRQdGAGNxRXvF8ZXLrQp0S/UIH8+RA9Fm3YZC0XD94hyt+PITgzDUZuBuI0p2
hxvyhk0yrGprt+HAJ9gDRfZIESPx95vBjyA5b5q/OhlvmB/Asg/gTceRrfn+WEko8Eg01HFvmLXg
bIAYu7/xBtOGFi9+z9D7Z2GdBnB/8/f1iTnbNqtEqRZVFlQAKbiB4WCx7U7Jc7ntJPVMdipZz/Cs
qrWXzgxp28JtrnKkwQzyDQUzuFSfjEegNURf4AnM4Ugws6GARKzacbf856aKIBdiJb8y1bwOUR/+
rlRzk26R8RYr9EM/tPK4Q5uc0Xj6Tq1xo4dMQEdGVLYEdcnRcIYSiA54EKhoHwbdZ6soFt0b7Z1r
03AS5RmC1xuhbs9dNQqCVhON+zs+Mk0d5m3bMSSZ5to5OtsvZh3/x0h74rliMt3268QzVwVE086Q
Xmjc4e12DbIboJwLbAnU65K8iS/DBuuc2d3bKdxEc4G1SbgL56exd3MVVdNkFFNStVt1EPBh5ArC
pbdtEyO7a6PWP4RC4yvtV6H7UXyJvAXjoiYjykI4/9fRXdwmTKRDa97sNHwmBC32j5hukSaWLuAz
d8tzKCT0zpELcGDtaNphDnRcJW8P17c7ekpBoNc4vJqrah4DIlSqqQlZ7Oe6lTXzJrhwEVwKo3Vo
pISm2b8StYwXKOEinoUd6DO+t+9Syeg7cuRdmvIf3CaTUMzs6Kiq/QwvFo6o28m06zrLStTpFtso
rLQzd8g7NcUXV0owB5Y6Jr/4G/8nn30cEpIxhNHDZLHsrUZ0pK3/YlE9WULgzh8u3Pd01jRO/ZZK
lSpUt5Q+YKUWFmoHQ+oPOmB2f/ZQmsx77waVMcOnCL5XMX1xf9vdcvHJ8+/6Uxs5vWzao727mXhP
ltV+RNS5ngOnRkjWa2kMD8xMfpkWXBJVUUoVvOzXbMCtarpcWm4gJwZQzPwaFPdz/CWcYRiOp4iH
m4mYrz/KE2M5oY1J2J3edjThb/SLT051umCmmc1lAvaXF/FMW6Oc1KUQkY2PQQFvxjk4cbhdA4L7
e/5HU+FmP1QzNgX0L6hw2lGfYDGDz7uZee8cE4jy75IYtPZiugRqMF4wKFo7BtM1yUk5FUMLHmGi
bTOEBUgzb7HhxMk5O8t+qrPOC1kC3LChh+hNx9ZpUAd46B+JWSMmohhoXT4+0OK/5yMh55EcKxaT
FUS4liZlXrhYuZf8jeTq5QN2DS4FUuzN+gyTc93wrgEycSRbrO8fWRz8gM3GRtYUs3pI1eaU5pKw
LHPtHXJfm49b2n3Tx5kt4/bYIH+7lHqOrdj2O44GlfGuVlepWW75zcOI6nluNEb40pdiVympBPZE
YsZkghi+cz+OaDATfgzunZ3nmQVWMjYwvcqu4RGlV4FYZffTjlrFV1hn9ELL2IA8KoN6GRIgpzeP
eVoEuXlaNTUjulXFaD0uyjWH/+5H7W5J5BO20A2xZR+rlu6OBBzMt+AETrHUP9Aq2UBxFQx3a9Tv
qfcFHUgfksmnJ2apNniWYgFwNW0fX1ktsfYiv+QwoTAovnxCB5yYV2gwT8W1F9Jo6O/ArECafTnp
SShvHngru8GHv3R6Mq+lZj7UGk2vsyHkxytRy8UW1rbzpTfS45sy6+HJyZqhuC0gJ0BYPM97zMZi
pflFR4PewpgMYWqcN2rzPAAKehqH8QxRUcSiUZo3LQCgz97evP9+NeSRtyeYPxf+XM0kjLFSe+VF
0TGXVaQZxHf8OkyjgYjq+vDntwyPIehnObbNB356sLUiRiD0ezh0f8lW0bwRaoxXr4ZcIUP0X5Gr
ngc9awA/cLI5VAMVNrtYqwufMcBXUzTmnp9+3CgGHeuPq+lHoMUn4EwoV+RBeuQM4yWlNjg5djsi
t6vkVFSn30kpQ0k7a7WZlHti7AKDcNm0MP8YuKuj3zwqjV3fcrWNtsqfWmCJ7/rtVoQE3gmVAVdv
sM8nXTG2YlHWeiLfpocR2BjZ7dDhR+uiaPrKFKTHoS8N8PZIyjQmlGsEvVnqvxd5RpTWugmX5+e4
WYvmG4BFpf+FR2MZtyB/jddfT/qJtVhXdJ4MFVoO7vwydOFBHKB1j5n+AY8XG9/MX3gNLKinnhzO
OSo12pCv2xr1bheXMVsKG6Xq/fB7LLusap3e7IcQg0muhj3NDY5DQjt1+7PXb/bRTg97+cv9djuh
pa3e3rSJqkPR/9+h64rD6Z+2gl3JBt8TqNUrEvLQnstP1paxQv6fLi7FYipbQXXKTdKuzgd5NXSo
p2QV5rDpzrnxDsDUVk45NbO1dB/pbYhEKl6ZVFRTtNzoqLikV6aSoxAitY4JRlmx57nxoSe5T6l8
jgt5ao3OZ3qqpqTWsWrgEEMf9OEf8nkSi/qp/9oAtsV57tA3g8JNmRqs42njhojOryix8juzWAkP
6gMnO9q/3sk9cxj0VOZAcVbMviu1zWw8uqhScn4qn+X8oCJhndJqglQ36w0vSGuvcX1EYJegYyl2
CCvSD2sO3qrQGnGZ6KvmGZySjBklnTiOZRFhC9tknATwDL6z3zqxXkbJCGYkysW1tsCfc2DHB/Us
FUBNhxCOhamcBFore44jFF35p7Begmyl/1qVoYn7T0sJ9dcorxYnpil+49DMiSBIfXgINMQVzz8E
Dt4rusyx/don0pJfr4IlT5woWfz5XZDI5fd+g3Y9eX5V4UjRJp5p0DBmpWaTw0YwmpFcfg7D1iJp
mYThnG6Ix127SBtCh8ZnKLAmp9nRozYEZk3NDfY8Vq4zbxwEp1anjA0VjlA1AAHvHcxZYUEBtDMC
CcUGfIEbnPdNdiqUcsCt4GxjCD2l+wzZUeqnhq1us7rcK+7+21KhRgp5x7rjyh5tBNeggP7pImU+
5+izpDr54DZAMtDlSCb3VPt0SMRcjiviOQH4cvZcUEr5SaKjwXUamn60aKZKIv9aCYkYrSyT67Lm
FImE8+kLSmHhmGr5Wu4YoX5JLJ0eqFJOz76VtNKLapBihmV6QYYWua64ThG8m5Gw8SlaZrRlL1Is
5Gc6wa4m7orgQvzVX7BCSVDTrpL3FO+GKX7PeghykELd9ACKBUC/VjYOz7sEZbOTu4aiSEga3kQ2
XuCMPuK8OS1LjbQqrav67Okeu995t/Dc8deV9+f5kTxTkhhy+Gmkhxb4C0I+xGI9bi2gbSMOtkYz
3o3XHbLNmq5O9lH2YPTnQQfJiGJ73vOyvEus8NACXcLVqAbd8lrVnuU/MdOkyaFPgBlh7pHqKUdT
KDAxuEkW49vWPS8nwF9Bcv0QEo/2iRxT77QRoKGaLVLJAFCZAKHl9zGwfvNe47v66wYkdNhtzNnd
gxRrfIKP3z5nwWklBrv2ZCH3l/fSMvWbI+fxYZCgoHALyHn5gnqP7GeRqV5TRGgiHoupRUjaC/Oo
NCBdtRneEaHjUSmwTU2dAN7DfHTiLNCyWGLikgHGfdD2mgJtQNdyDxvBDb9OFLWd0q6KPXJ8ijbm
m7+epi/jXUzJAIl6RdMV6skaP2rfZ3WJ81ET4gLn7pl2gw2bDSopf1pD9nAHAzY2A3nTt7ef0m6g
PXBhBSXt4s0NPY8lwGrRi+/NAmNOBFKj06d+ox2UminrnanM3fSpej5mCb1b9bco5s7geh33Kry8
+A3PzCYLaREIUw5O0YFr4++pTpxdOnwoEqIQuehezZ33gAjJYA3Lz9Bx0zmv6xS0glTCCNDuQ424
KfrmZO6L7ZDg/yEPNbO3MPxWYBKErbeqlC4VnDSzi4NxiHxctkVIhoNbpILvUADA+WtghvqkgmxY
MAxEFAxv1ys4QXD6rpY7mIvmryLZRPzTaoChLKnVM2T46iUluyHcbqeWT9dj3jWLIUqx4h9Vfqnk
4+45KUJiJjNlMPdhKhc/N0r4wresuLfaWSOzNSvKVFa0esqkUK9//O0Dv2/UKxhzRx6FS8oZedjB
28GJyzHgFt6Obi/8OHCjdvAZ6i5N6yQo2t+phCgaXy8qmgd/rQYofggpXZm3z2CDYFjDtfcQso7S
vsiGW/QiAIeUcsOef83EhArUAzlXIkvqqv8+B+W/YYTXCHAf2ZIkFY2LQ/enNWZGfpRr2luA4zWh
JVCKinWo/GXBZjqf4zNiXTQnNx1wldX0c5kqQZQzttxViYg3hVOv9MlPjjaZ3vfFzexn5+o9AbY4
aM2oDfgX4jZnRQIM6pM8dLuatWOi8iFLZSSfuOdX6VSYV7hghSCYn5o3PZ2UjaOGcudUHqi3jDEp
yJeEiDj+NesBN8Ohd0ua58B4RRLYdnw+70kaoc5i4fEhPxo4RM3cPnvOuaNLwM0cmNYJI5AVQXJX
pMfHLNAfdWnAECWPhVf93Y8DDSR+Yd1BhGZssZNBnqno9lV5qs/avvHYBXs5tIkdujq1jf78FWU9
8+feDONczMEkexoCJdL6lZmJOQ+/mo5v8mUwoIlGQIRLTQwVRkob6fu7FPnugk1BybPOfKS8v8hW
uoEQU/Se/hjZWqoaIrw5ZXq8pL0SZKJLOZN8kRlRnIypHiE94fHRRK5sOF57dRzEDqIXcjAoO/OJ
1ig6k0jEiJKerzHhIbEOXyIgQvarZa1ZDIMlM9ciu3waUHegFN+x0g1Cs1H0tO27kx4ejAwXrnI9
GOi11L7N3+K924MfVssYZYX0aHJpfu6RKYGMrYbD6z1Bzrx/xevzd/3mZgbY/URrr0dfFw+cdZcU
K+sDXgoa9KtU04sbn8pzK0G0tdourn1mH6csaHw6qWaEYjxcWLgQ755xxmAdVMAOB4H27mJ/0iqv
CAPmiSz3KFvJYSf0vOpUmfmXmalhFK5eeOE7sU9zN6bUOrsgl+PhGpmEnn9bpNVHI1NaVCtJWLyG
hWDztw+Lrr8MK2Z6NWtC7Dlz4vW/e6IilF58oLYXrSm5QCmPdUrhiR8AO2kPgx9vGeuG9fN0GrJj
p40izalHnKjpNG30LQH/6ZAvLmWrQwlcy1bWhW1CK2+No4ejrzNEE+KM9cX9LsnAlZ5nrkzJyWsX
3QhlQdhXTSoksQ7pfxLy0nHBcTLFLtsnX/nT/DIFwuh2pX04LVsknD/8vETDHduciyRngmyH2SPk
3N4/pKEbM+I5PDhnF5d0XSsWfVUNC8za4gjJM5JeD5lUnZZzbFtweI3xdNLgN2QkjjpQCFInCTUe
Q6eUx63NIUMyu1Mo3kNUzbHx6cIWLpZEYg7H00pFd5w4ros71w8qI3mIE+xxPCbqYBURRA3lI7wY
Zq6zDcvFCdxPKnt6CGdZoSv60kxWTRTeo2U6Er/nqaqBJVwerBOslbcfm++VhRAC6weT1baYq5Jk
BEy8WrT42x+YoYb/NK/wNVGT3MA4FFjzZm6s+9Qe/sXL+YBQLWAfVaFD4e9ZUOCTLfwqO/39K54K
AfNMYIOdR7HpKbJbQ/0MrCwxgSFxynPjFkUzmyeLuLlL1lOLv58xJlTTD7Gg8eBJxNVxsd8rFSJb
bvOko9dSgvtEOYO5UENvPZt+QACD90aoe/HqXUffpdJH62AHiCaHHuegbmSiaDo10lL/LPY4A9W6
8zv1WzIOIa9doARXVVVaEJn/6m1/CvO7wrZ3xydR6Er2xTSLp0aBXMQOAgUr2qyhzd6IdFi1czVO
MXIxmw4Ncc6i/AxaPBkYlsqkq9vFm0LCsn5x5IWkmadYlW3MtPv2SkIvXsPjixU6+dT4AKwYq4uq
fJuAvcF5J9HMBgNVjWhhiHFSzC1XFPYbgM51Oz+a8U7d+NbxEh8smiuH3x2j+ZPnL7KmDXfowBuP
knIgpNHSn3F+5WepVhFyIB+2qTowxpgKuEXIOWgqUA9imh6K4bCZIfL6LC8skfntMhx8WQyxHLCb
7YLmiwz/47Qc0eDruF+My+9e15k9OSxShS3ealyjzNBDXtM21GUKoapeHh7G6ov6u/HP/vaFm9Yp
PPWGeljwKvfaEsNfDgY3PrznBPzhvCBkWfGe5d8B5GBm/zmsTs4sWSpjb/NzZYy5n9Nb83M2TqYb
ja02PBSFIGhnwSfYUX5fLPzOkgcvb8lk8fJkN6ZDo3u5MZWtvG33OTzf1mt/xSNrhJQNL/XWqEGu
t0v+ireYZCtdE5zKtiziJCPqyFlzZ7lcBdIDVTJERo3AZKeMjHdFRIgm6XjlfvbXoVVICWlshlxu
uQHsYd6admJVVMjSO5XJPTvBJCHT+l14LvqyKqd0HsBJoupWzmFGTUXj4rSXbYMAu/RoqcakNxKz
mJVoGoNsf6nAdVuJdaXgv86tBAuqgFMVSnB+hTPdehe3l0F4gsjEWFqqvYDssXJAC2WeBbpaoc4V
6R+Oam9hsJwtC+mx9zXvlG/9n31hk5n+w3I9nlVv3F0I04sRrsAUsNBBkojdDwv/JdIX3gQ7K451
REyJj49R8asz8nMzcjjVkjR4VzC4cSHg8TsZuw3lHPitocg+Z7kPovo3qiheCctr/8+n67re08rx
xJrAF9L9QWpugPdPidpdiWCo5d/r/ccMeKpPjVZzlDqoVFDF2bZaWHSBrSnUB6wFfUFbLBQHbLkI
HUF1M80Cm5BrF9piQe1cVLnTyZKnPgwLk8Iggh94cECWmfk53fMAAdyGUH6Lm0YRyslOkgqFJsyS
70/Zb6yj/67DsZDBZYv38oJRZuJgC40tF2P1FJHGsjIF4LasCHv3wVQk9sMyS0wzX9QsD2KkHfDD
NOy2WmevvF7cMq+j/OKtpCqxCzJSTYC7LsKv7Tdt1lkTg7EixRF03Xoh+isvxOSW+7q0c7DyOxBS
igdC6hp7JcOgfsZViBAS2yM+gA6ewcxFsGme5YpRVdPTbNAsnVWtvYcjD/Byuzyh5R6GnM9CbtR/
N9E3kRslSWgLNNi9VQo87uSzsgJv8I8gN0gl7V/NOcx/3XmPTUA+1FxOtk8phzBitR7S8Fh9ils5
jBxtP8xYAvblSNGnVqAUZ1tG//PJdi1llBB+zIJyoJnuptvAPl3g8ajQZeGJuskQVMp/eDxutpOW
OKNoin+ZKXFJwdi1aiS1CPgPfSP/2T8cbcUejAi2lzGu61iEkYIm6sz/ha9hEekwjvm15BAQiCNr
7rkFN3jxd3S5YL7oQogdeYy1MoTrwBsf4AR1URRAvd6l1bxg0ZB2/X7UZCwLzQ69J4qUy1y0S3TC
9rlFt4teanyIKIqHlaIdbksgcUghvkq0KyRE0LHn9t3S1dGXqu6uSRsoAgyF0gJj2VnhPMS0eCyZ
D7X5R8L4NJgC5YZYPQyAwSN0zXprakVNnWpEmaovMQmZpfPI80AO525vnsjCIiVenCINKEHFzk2l
5yLcJqWzAayqbeqbgU1qzhkjLO4IRCDBmyUAmTaNqKn0A/0X3+KWWpdBiR3nP0P7CzRlvzaVR8r9
dAISIiLi0NFqSsY9RIg0yNHHaf+7dV1SZcJzWqxoQk8qbrDA/3rfVH9gcdf5MEuC28cmDtAru20H
l+LSLRS088jG6r8XkUUBYaB1tI5LazX+CPe9Srh70rSVJNciaETRaxGTppLSXl9qc9OUNexBa49G
Zx7rcGb9teEZvm6HNpaDhb3PKJ3b1ZOp0Pl+cUtlSUU86/TC79KYiqm/arY6ccqEzZGWTkcLGE14
YCjkGp7rRw71jGSIf/njojKaDLnJJI3LlqIBUqQlMFeeVCUS2KBIHoNpNU+S2ZN5b4dIhbSk0hB0
KNhIoJzaljX/HU8ZLDUd/HWLVkYpn85+5lDsNyEnFtMwy/8PwAYyTFXSe9aL/VNdL6CtAnJwmK7F
MJEnTD45MTIlOTsRYtPPCE25evX7tv1Z0rTwqeaxoS8tt5tEdoPYOIbcF3QQggo4i0kSuafR/Snk
H2PxNiJAzF5w+rG2XJPfvC1woKmH58UrmYiQTa9p4USwGS1RT5BCw1JsLO8eQ53k8HfZPQT8B0h5
GnA+6PYxxtiRy1Q4ZXRLTvgtS+dUsyXyJSUip/J9kEnLGxiUfUJVP9WjrzCD8u3dGuFKHDbyd5oH
s2D7YA/u4uLw8kJdmdbo52tgm+cOKIbRQ85WLfsL2VB9ozCNN5vSDGemnCVgGeQXqxDQzuqI13YX
qfoxLxQ0s5kebG+51C24XHKyrWW9ztIVtyhbXdctJx853monkvpJvCyxN7A3ItNwD85xqRmB0a4m
TI4XPbRGwItyAYXW5B9ndyDiLhQuut9dNHMRNizAjjR4PPrbeopZqWVPxYs2aBbrERPr2BizP1Oa
Y2zl8L4MAgKW0h/HtgUpvVjPfUBga6EW0xzHlmqJjrwM5jCZwsR0SvUcHaBpuCFuvMwIkDKN+XOs
LMwT87FIMPaSCtFPwwer/J+c894KjrcfLuFDxaVnY8aBrIoJMQq2Vg/NjAvNqVh1Kq0RsMk2m6rR
Hlh1qbYEOaLIihwjfGGF1cysDBsQXTMZgrWMsmgGKr/rGCbORjuAETm5w0Bq4Lbr+9cZBzL034Xk
2aoTOVbpLmF/+wc+Nh9UJ+3F+LCBmeF+LSbSW52V9HLXYABkt3QTlDETNZrvuivUgkRguAYZUb+Z
1i5n9+eq31I9Ao/DEE9syqwq1Lok2Zn4LGtMoEVyvzCXJKp62nFIQA24vBbO6fFYMKZRF8JzfJvP
+wdwPl3+b0+tMST7s+FKtdX3Y1MSOtyfy1aSk69pwNq/FIros2qiz/VqBOMrSOiFH0wZqZWzn+6K
zg+zo71OUvvu6nKYhbsYyL46CRWYcdcXuNGmaouNcf5cRCX/LXMiGwIGz2NKqtByGcnNxa63J3j7
qyW1PZKSHb92g///6MwUl44tzMvzPVV2KOk0l3p0sin/RSD9EzzCbf1tHitJGcF4snY8Yyysloe6
VzGkWMDDXcmyQ1P2tCDE8+4HQGTEEdk4zg6hlVksyI2cLw+Dti3S8+ufyTFw4gwqeQNfe/ISXF07
XM3QXcqbmSk2P9eQUrR7ny3kaD8LSILCvd6FdxZETujhudANoiR+QVSX4W1lj4TnrQSGTs7bH/po
OK7GBSyeqnbP/oyl/2LQRLy6t2M496NnFGz5MV3sJ+pvdzBMEU+EhNgsitQvuK1FCirEIqxojz3H
CoOrmyGjyGAJopVg5+J+oiXZeYuOKgs1aCErtQwjUztcJtS+0EpaIm/HourzHPKaA0yZ7lsRsb32
LrkAAVZNTprGRvkTjcBSq6muzvP7g6injmpI4zSxdVbrZhHqrrrI5rYKX4jfIv194eGtfz56oTnJ
UzbaJPJydmYkt91qXl4in78Y7Qs1cuxjYtwJNpfqzqFa4QVSHtQD063ZmhH+ImXN7W2Hz/OzGrLd
4aHEYbSv7MQaH0UoNgZew0+yJ46diGedNoUICweIahzJs8NbaONVGOWmiRUxOyK1Cw2yxlrW+HXu
LltEQ5KwYkSBKhuRSA5xmywBrB7AoGk/BZmtYh8E2xeK+B0xeE7VtUIqhPvElgiS+P5GkmbJj69q
iZtBoE8sjCKlvSVnwYyjGH1lg2FkkA9acBTjpgPRKhhnVKDDhaDlqKVrPwXTepMuvFx+jVl0/Wha
Fb8n6K8IfXWmmW/FY6lGN57ag5Pv+wxHiuv9vyrdFIKQfSNm3hY7WZ229si7EEmPsRx0NbaRvR/2
wX8ODOgvdZLs497pKNhq2Xsi3gcSNrD/8xqZ0KN8MnjBGHgsfBeFIMNxqXCiJgT0HAk6jZHaeQx+
wwQj1iWUqRsGd29BkqPlZyWRs6CLL6LqXfzWNTca3qL9UDiB1Woe6bm6u3Dtp21/2REDfgOQw6P7
Yd4hWsYoc5+FzkhzCBmDvajgFOSRP/y8fA61YGjpUuc5E9E0iEjWl1tl4iUacQ7AE5F7UC0LInzo
M2H1jTfD2tJoZrjWox0h913Xf6C5r4kNvwbpDWZ36uXHRGfhBReFbnGe4CEbvRPQlH85g8HgA6OS
/blfD+pXdYFZuDTYNLD7EyTbhwb4OTKuzp16maXAsfHT/fW432/Ofs5+Ff9dYR4eI4W+6agXrBbO
aCvGZW6jYNORdSX6iZtCGfuWC77x2krWnckTMGwAFLgK3KbyTAzeeo1a2cKYRzKXwmzdEpFQeDo0
Kpjemu3ILcNrNBLVKHssvnlj6L1IDbYTfaXg+9UQyfNu316cZ8OAFsMol5Vnk4L4X7w08NM5fatY
tbf5mWE0p/+bjIL13oWVOvCiE5QQ7iolnx3Zkq272KcaCDajIsyxTfXmK7qwDDaz3fUrFbP0qiN8
+QyjjsvNDQjLl/oiJii9u10OD/bIr1uLnb0FqbwDfFgR+ZvO986YEona2DyZgOjdlLjNrpqBM9Dt
B7BdB5YYa1ywoNUduAsEIJRcyLQhpZT9pZFNUYLzUjHixKRoWWeEAkcxMnYcAfjlPvEUrYz5pmjX
3JX9pJbGP+ziqL883F+NTY+BevpjlwE6gOaR2NApHPz9hnU1hsyxpCV4uDq5GQs+pbR/jteqEREN
rQ7uGd0qhy2aOE2swzplhaEmphX4yDY7XC8Qy5pvYnU9oGERXahP/efUl8fG6xacY7YyFKxFEhtd
FgqaiDI6G38Xze/tluMPj37W6AQPeNkKGM8truLf/WqHfqMXtxc6Stu1//SPPSGGBx1+vnXZ4IrA
T9Q6LR9AIBjysg/Bnch1/PK0Yf3P4IjIhhAaLwObj6hNBq3/h4L3mvLpcyQ7mupvSkF5qv3HIXBT
4KnjxKZ4aWhw8zD5148Z3ol7BOympZbQicgQq3G5CyY0Z1VxXJ/61gXDnXBXtpVRE+feah9BDAL+
NCjcNGbQYfh46YGVLxdhRGJjyCWCBqnlA60jujT9RjnGGj+i1J/PXq7ff9rtIkUUVEDnYT0+PX//
jaNqFgSkBnK/SZ2Fc+hdQwcAfgG1lHUC0CtXJbq9onISosDe/Tx2/Gx6qoQa0PKaDutpIlr7vxzO
5W/KDnna76PBybemng/1NMBdr54KBCvLHahIX3ib9dqvuEpCSnQMCnSbuGgunB6vOtvBO4cUW9ud
bTUU3y9osXHFN8ejFt/bHi/9UKPnr2Kyu1XklwN6Lg5S1DYKmqqCPI/GnIxBj+xvFRapu96HODtC
ykjJVjn0YebcHJILIaBfaBYPwI/ROTL2TeX9P06dndFozAhmsSbCmvJLzDjlE8sOi4tCp4+3SFWC
6zOjLSOAxTseb04Tk4365qZQ6dHLuD1j7A6q7zxTmK7/gNAmGL93vdjucaHGt0/l3qIBI8DKNo7s
TaEFaVw3/XfRw+DeHUrbaBwXlvooSHpP670XS6C7PB9Ml2hc2W+Dhx/YyBKibs4nlfcWikxr7T+D
DF84sZQOrfRBvRXl8uUy7bWxhoCxhYUamIJiBzp81bJoaFtJjzx+F9jl65bTDypLrKUHozCPq1L9
g9Xh0TR3y/ccgMG/xAwX/EiNloNY3L0xpsCxv5iESzh2U0VsTVn4qafIlT3LJdPgLZhDUyOCkmHG
MDSk/GsBlF8FPbH3sfuRX2l3bsQHcWz5Fg8oakW/jzijoRCqD+wcT1bQR1/cYVVUCuBVPI0NlV2/
1VJrO0QKj9SOA1c2JAWf2ByFUsraGBWtzlJJ1qdOlYKV1xLQ3s9rY47FKvn0p2OaAs+XFBuNSBCu
VFWIy6M3iSgcpjnClxKprq+H/m9quKz3XHL8DpoBwelBQwSPpNXZQwr0KvDjpiXVtaMd4b5eKP6O
9oz9LVYZ4daYzhx3OnNlMZd9S+mJzHds0NN8d5NkGvShjbXj2e9sjjz1B27uJIzKdee/Se9EZ+KR
DEC2PAtHf1G6Yp2VhyO4h11um1FyzJMg3lkh/c3EI6dyw4r1gnuBTcVRSYARNJ7AcYnhGHuTb4Om
K6j4WNxSlULinquajOpBTPOu2rpKxohtvYdBLcBOebI1BacH6Y6tctxz5+qHOlMJ4YvdI2JuIol8
2g3ACMYoTs/CDf+a94YZsN3VsPTL9x+KDX/J6xYT4iPShyBMaojmaKShX2gSHt3kO6MpJNPXxlYe
monS6VBtY0I4o+qE+cRbv3RRWJ82TvdxOx3iapbHAMnJwbHsjZepP/dtZP96+FAa/2kXsgQ+KXNF
2seS0uSAQwdk4EMWDy00ZExD+fs+hQ6jlzkrPYLrYJZ4wZfRJ5gbZaTA/4j6j67Bzcr1m3/oHmoV
Rod/xCi8B1G0mdN3ACPLkaiHfztW0xYeNaUWZOJhAYQnzvG6a7+PJe/vdX7vZN4gDbWJB6iFnj06
QFujnJYralcpTjT5hO/tKbxRG2PJn4/tP07ltgXYC0+v7lZ3pYriHC11DGP9JpnG4hHyVf0MF3eG
wSNh01L9fN+GVAoWRSzuuMnhvmS6jeCc0QdlNm3/fcDJC4YFFaYk5kUGoLsrKiHkH6dkMsufmCm7
xAe+eIpKkKmd4Ypmo4nSTw6FBjOSopmSu3XFWJE8qBHFPrg3DBbt6JfBKO2veiZk9FQXq8DwHsiu
Pm54uhVvLbnzEicWVNrkx1pgOHb2CF+jJX5ci161YHCFBSEXQeK3qQwpdIKJOVZ+qoflEjRH1QJt
sxaSDxGox/5yVZ0/154inu7YvBI/v4EakfvtiXTgpxQkt8nPA/2tSwoihaHSKQInyfM7Wt/VOjOI
LIbU362t3yUKEcNTpxp0aoQFA26VPbubyycgSVN4GTISCDmmnInBYtc4C5E+jtayLJHS4pYkyxwZ
6zZiiH5nUHOmoxn7JcSvl0p/FgCk3NOA+itlh18wjS2BQnejKrHdiDGfFyrPxX0K9CAvdBb5TWux
ShlXGymzD+3MhD72TGnntwAW4G+APk8rNMAUIgjyqS6dXyKBB2Yz4r+S7N7ijhOihw64u0WrDGq6
GWNu5/d7322+ARAYSOJNQOaQvxC0BJXkSBLuGNYJYbUq5NRgQMQV4a+q0R+Z4Ko57xWK1yIPwEAy
wfiouO+xm5A3UqCRj8tYcvTYj6OvlF7jq+2FeEwUIfrjqReJUD5tRAIFbVhcvE3tOK+K3+0USy7D
L4X7Wr3v/92wQBSTWKu3WHs5f6AzzyrjcJCZJvw9Bcs1fKLAC506Rb3aSXQuKurnEnRnQt3X1ydT
evr/Ys2N3U2loUmq1nFrjAxN3GuqvFMbLvj0kYm1H1ShI/hlH+HH0dJHGA9B2y+TrPEErPG+bBbC
7EF7mv/UhV1KvVtDilazqBQLvumjtdd5Kce3xATYmWGEWBaShdcDT1ny5vFMq3U22OD1CSU1Z3h2
Nsd7tEM7y3/m8cZ/FnYViyYpVc6V65yTxyN37wfF5ZID45RX4WMeCpNLLOWu4ws/Gtczqx7Z0VGQ
XJF3wDGxt5l2CobWkM/gTts2mP0a2hxOPCL5vJ5m+iIVhlVqx1N/BFBmEsIEqcepY9BedA/Sjy18
rE9VJuE3/AT5EguP8Vx94+dooblUCRge7aSaava+il2Uu/6LT6vlmWAwuGPW7I1cpZfUOin0wWOe
z68ag8EUYsDSkFPtOGwZOrby3jv4zxmsgF2mfBy3m4q1H0+pn6xdDnmJcobmb7ODJ33h5mY3ojT3
NcQsLpLVtHxVctncai0duLvUcdmk+QVytjG9dWuBUxQZe4BIzuEW1ONZ7oOuWdKnS7KhQfc3FNdm
kev00gQxeocIp418AIK8psAbLTpuIttrV9Ayo4RIETN5/tkcmmVymK8acAHpEFkmzjwwNlSG1WIl
ZQTcJgYsIbCo7XJOLiuHscPcwLWvDZGlJRPfoMNAT5jR4UkdhS9bZ6gz3A8qd5ntprvwGLuemqnJ
Lx1fU7trvhoJB7SCMTBF54ImJYOGPoZlGdlaY+/nWbOls40iOgRbYHeZVGyVK7Ao01aursxgs5pU
V3wBFNgaP34GhF246VDWSsssrlLqHi9YbwlICO7Zep8cnkX/efZlsvnmxyVkQr8das3MCOSrzntv
dE3zdSrNZnCBWSSaPiEfH/8nq5cp7SAaLPO2qudgz5aVuYO1Iqjj5l4vZUtcMbXVrpbBv2BrXW0C
cv25mZ/5gBswpIq019WxfmGPWX2/QzFLAdbQXJvabPBVW148CIC7hvnnBIfdyugAbwdXUlpDqsOp
7pSivSa2QOz5xitlezO33xZSN+JcntcmAJNXeUhUmsRm4mauzeRDAWhM7hohrYwE+FaH4G1FRL9y
BjNVoS5loirtBmOyHQHn65KZefEzVh3PFVF/7MWfZYaRfu9s/uHsw9qJjSS+urqQ2+fs5XQd8Hiw
/pssjHRlMpNbC/u5+4XD5P+RzBdXQhKXrNCryPf6Kb4kpBzEBhe9rhysxK93UbV/E55kZOsxlN4G
7OtMF4eSDp7es9Kik4je3xHfD8QcVbZa07zk03wwfNI/mUmtjGy0DMumccQeNg6jkEjRyDayw66E
CWXi055ry/pZN8T4Z6oHRk9/eRMlbBjD+4NLjrLPaHjxSSlLcvAO3xRmNH830p8ilTOGeJ1PmTkL
5zWJ+mejr89UCYDst5VVIE6rXgglVPxAHDJ2Ssd8n93ZYgrF/hTib/qhh64YcbvZsfMbSS0/VbjO
+7Kbc8D4QXaMf3QAL1k15aO0Dsg/Z08nmpdTfXl3qNU19cDe/44A9DrKbemDLiFqgc/k/pHirZHB
9c5Ky/rt5rUf5E8e5/o3qTyVWRoGGFD0cZBKURlRE97YOM56C6bpgyB/FH/MkJ40/mPTh6tGR048
cFYARbAMm2AmzWF4eXVto+PTLd20m+D4fRSSAKPjDnOC0ZsD7/RimfJn3aTPFCJAUj+mPz0kyzdY
VVBNW89OMkXmr3ywiRgtmawuuo0LLMtDhUt7C7A/jmI/AGXfxlFxbCnLIP8WMiQte5jBrFh5DoiG
OHuTn0Le04QED9GZwwy686u3V732KdU77KwvH9k1IxuRUyhU32mM1kM9p0tPgZ7mXhDpYJqRXqW9
Ap8hG50eGM/psKX8ZF5J++GpYjNdhAWPijSMICvCIJzT/Jq9yeL67LShdLKav6MvoZb8ZCIp+bnY
ZWhPVWG6t0W1dkbkw/XlB4I0HaHUq7NGjNzV7faGyuuI/ZO6rf1jG88DiAV53ZqMixrPqRuygLW2
zO4XSyJdfNb6OzaUl0ku3OiIIxfhQH1ltEttN9M4SnFLVE0k5/tvQaYclsbRdG81qylPS+YnGrIB
d7Wc1sG3WAy5diGvFp7RxXYSBLEueQQNVSnObTU3YS8BLLxZx89nlv1CXQhrQCyEuVeahvdq//s1
HhGYFLCm9FPcqDI4tFHBb3Q53c61tEEFWf/sR4owYIV3LCj7gYUP5YLamiL/PIWZGQN5Z2lbAw2j
d35nlwr2/z6dByIcmaZXRQDMOpe/cshRomXI6ZHGt1av8SfZdPctVYUO1JMO5OTJN+gUN3t5VWw9
GszE82H3XH+jS0un+G6HFoljdNCX8UaED+yp0uU5znDvauZrWr5+EhrYk/g5nfqx/OYph8yKDqzq
YiyvVG5/c3ZfOVOJAdKeo1sq4RsLfBqWDUZwz7HJ+NmivSq832xw70/eA0tjHtQMw/3vjYcNHWHD
PX7NWmzsbg9QK3Fyt9bGd2ZbL1AEAfl19XszK46rIBusonEHTEJlccCL45fCAQ2hsYCHMknSGE8g
tKmnP0wBUiXoooOe5uHMGgOVLs7Vm4TUwRlWt66Tyv26rE2kqD2cCozIhKQ7lh568yArBCkU+v0q
AZqhK49/mWuPmK4ypJBBcze1KGd6UqI50inwSeIR0knyvRW/TAxl/hSVCdtffnRZyDNOXuOt9vuh
z0faj4Ec1urPpw0U6xq0EqsR55O6Btuzo+npBqE+7aeuX7w5Y2i7LU0WwfJcsF6KIlnG3H5RcRAS
Kjz2H379BHERYzZdttd+FXWe79CHSnuu/16E1DVV9W7mJkBphlSRV7UG6A6O+vuBs7wzlhd3i96K
nYYlAAA5oSt03FNgDesvugdzGOwBN2QvDB7+sOyO6+ierDS4P1qYcUnCkipSZuAOXa6eYRHgVHB5
sy8SfF5d6rENoeHwTxoSMRuZt0y/ttDO5EGbgxAGcsURY0nymK8tYaLaXWG9Ogfy2zZzgRkDhmiF
AK23LramFz3RWTBkd76nVYO3cLosWccxfb673V7F22dIRCEXnbOEkf7313z9VrPOL1Kl9/5iw/Zf
4xEG5ghOMA+m4/kWi28XvvBv6R36dhnnqMmVMvkKTlDLJ19DboPoKWJBh3XMbV5F5HEQ72igGoGr
xqNwonmaLkKMiF/DxRBlOsX/n2pl26edfwgTRudiGdICPTLMMYs7Z95XK/1yHJ/64ONwoGBTOBW0
LYEXzp3e+kET1OfuvyC4tOeER/qtR7pdWRfQnKU6CtfWumkA4tvCDC7VFZ5DTe1jPmCG8IPGtqR0
DFg91CZFDxbgSp4ZRoPIAgUX+ejzaCRt5y34d4XTtWrdvtmWT/8fGp6apvVOzttxcPkF0xDSvqPL
CeLoe3EERyWvsByQ0AHiL+eyyGVEKs7VJ3GKJYtYWLjdofB840lf9Q5IAMJt4P/YNtfpuTjSePLR
SU7xquSePnKg44dr8/amy620JJTf+egqR/JTGu11w2Je+jmbY8ISCPe8vXZE1dpphd9Z7ekVCJDf
HSBzxkYre2mK3+teG7z7zcPlWe722v9kJAceYVmh8/ior0NdqU1I2VbpH04PndQlk91Q3yqpZiUf
PVbyElan/Ga0O3lzmRHJjA2smWUp9N8A1MVMFi27hnzkCriVYmVm5oBDDqFSXPvpvZr3RkldwRvb
P0DRqvQjpIODODN9EqdgWTkVwpL2GjNT0e5v/CfSHZwl/0cJxOva8YtV7e3XRg2x2M4nae0bYfqA
4EpCdtBq1GoOsHZAff/Ou7QMlk6OClWk6Tqap5m9YFueDbUUy2QF0gCcbP2b9BsZtQ7T4GP4Q+5q
hkQ/6+0M3Be3aS+AuTnhJVY2dqm3GHWcTTtBEEYrvvEEdS5P9FQ3pH8VwmJSTzhPifls4B4dj0v1
glApI6p8PzigKYOaWGFC00SU2URhjus29WTcT0S1TyOX9lEVSXnEAbeYK9LKnePMFUyNZVjxIHfm
kGYycKixvQnF5e5qasOOGckbxzFldl5en7ZofbEoYJK1UFPyPXdyBDYq7WStBD5ic57GogiT1lBm
b1WADSVsi4LNFM4ADG6LNHp6VgN+IRVM/jmKeETvUVHgVHFvG3wxl3/wbVXHddNeYM010iJXDZNz
+L3oh/LLdG/htMxPxlr4XFmx8PyTGnFfAOEiTl5nGmbBhwExrSsd/OqF5huAvuhutBj/Zf9C3w1X
TR954/f86YGs4QzEFxJBRTIpPCbGQ0j4TTFQ2b7gtgxWVgX1GnZsM2opbRkCH2tkm/f0xEqllUEA
FtQwSWIdU+2/efz2lk1WaP8SwbaBAy3oReAV3zLzgp/xVGEpdzd3NplOCY3XKAE/pT6/Y4ZUwZwp
mHg/Jtoe53D0ZW/mELn3PRiWkMHj0QELwhHoF1/N8ZkenMPwCv0jdHy4tW4BYnHcL2u2B3hshNdW
x1LcJ2aEoM59KBkXGyD3URqImSqxqyNcUDx7XmVIlpwzm+aFW+/MXzUY5gEKSmUJbcsHZtg9aBRU
JIOjMS42dL8qN7aHk6Mq7bnbQJe7CM8T3Xm3YoztROQcQZG8WdX+09gKfYli3G88KlM3xD/r6eiR
pgaYIoOicijFCtUAOFXo86iKaQEXIhYbff5mF8k/5zJjmHORbA/t4/PxgSiYao2WiwBcosihCLlH
2fjbz0CNHRqVRujlwZo8hX+GEkzY4W1rKSkpFIiYNvSH8Flfia4ZYui+2lfpyQ/THbtGKUcJnu1T
TVrXpJ93l/oBqrdnGAFj+R0uNZHgpJkb2wzqBfgh6zBGDc1LkZanA1li9YKJsnIuVAyzxKs1yYDk
Oiqf9z7J7H6p7yHjDz881OgtUMuFqbktW6vIFpQGV3/0QolUEEhUXGqWL4A0ZiEJoxq9SyQvDFqv
7pAAp+Ancaq2XXjg9t5l4D3kPZrwYCXdlA5jDf0wm8bz+HPWChPw5hUKLw+6ss4rPVHNyHFOxc7F
IrTiLATRb6TkDAqc7VaqM7uCzLab24B/PT27OSnL9sOQzXfk1HZX9cWhLzd78Gr6Hg1hR2R7GKTp
V71DTV4gprQJtVz9Pjl7Q40cDQNTWW5oCDfch3NXxuzjU1W7EkRkA46QWF13w5VAhCYUUMnP0atK
n7Nhq+FuMb/UoioLiihiYHirPTYUbS25yvaJpXmtvxvsQqGUt41W8eY3svxBi2fG/MzT0RW/lAhz
/wkZfLZ4kEpA+qmc5gyDwSorvblrQQYkVcA0AF/uU7mEn1GlYsPmseAbBMKhoXDuJKPNNFJjTsBr
r5JAvj+41Y8TbJ17oKVKsYWL+aFHDx2zzVBW8TWDN41F6WbtXpzD2AiqdCacC+B1sEmgG9BXAlTW
4IyShW5AwAh4SeS+vw/dmJxXhKKbZWlaj6vhAzZN7td27duy4oTu8gsMr+vAYyRZNelFuRbhpbV5
D3f0L6+BHlyTp5V6tDUDUPqX8uUsw408Vn9CfyaP093h4xHKuX/DDIcXo/EG8e1i6JYn1yfzOnTJ
LwP0eIhqZ5zn3niaEdhqtteqXbyje4ztgXzocRrEHm53I7HxSfAxo9+aCzO+9oF+8l4HpEyO6ESs
Y6zLjIwplMlqXK/z8PpVqkualGKfQwwUt0qtZJwBAlOtCCj32FK/9Sc02geTX4ZU9qGuTZEXZQ1j
havXZwtiYc4duRR3vz32pADIIKPD2cTQ1a4jm93v2AGlrx9UdjcrlvOvRF21rOwcivYS8FMh0ZI0
iVi1W+OVxWh8IXUQbnL/sW/LnUPE4JLRs0OJ9FfsrOWRoykZldzxX8aVZisWrd/ugcLIwD+y8oM5
omxB+QkLQV8i7QlvT22SrR6hpzfoWINNfVYdS4PtKlANA0QMCRB1rGDlvY9M9XLHyLLRaxvjXy0f
zng7MyD7xbGuhgaKoZ0SPlNe9ed7iNh+Cqm9bE8im7PIb7KWcg8M9iO4XzmpD/XhMfzcwZ29vCWQ
upL48QArFbb6CQ3ZHf7tUeaLUj2FipOMeTdIUjTbxv6lbs5bjg2+GYei2W9raA9Rr32g/PtWGQIp
r+ugH6VixOzVt9ODXZYgbJPY+Kfe8GorKhVcYxsHXPVK4q9or68eNGNsl5K+ie3hs1ryfxJBruxG
ED7LN4kWZ9upCZkqaTGjk1szvtVXmzx8zheOkVjvUoiJOS0dx8QyePWyTFHO85cT/EX6ZGkHvvzZ
yYSZX+tc1WoZuakLsyuz8naX9ndnHJ4oJOvoVu+UNdP0cN5M/j6PNmW3QoGKmiWtsq7r+SwehI+D
2Xd4vYQ+o9cloRm5qYS6mDZ2bZwQSa7qNgbeqwn4fpcxdADIDsSuxvAOC7Ewxp/AmbnvJtxSPx3F
6GECF9z3dg7V+knHRc4yYaOSWwzxnMnNdt3t4Tb0R3mVrG1QqHHnCXxdMheIDGrFdhNRKKTSJF/+
aaldl8rufy7eIsmbDmpqWXGfBcFKce1jbuN+vzT8fhsAH9kK69AiwZNc4S7C3RKZGhwUD2fcu5wl
/T3HlP/mhIHfSUNdpxMyicStBrB+RQ+1rxwcSJDpBli11DHX4x2gC+XKMTxkmGDQLvmRDJgkcXWJ
8UV3YZCNybt8k895LGgSJvsi+TGL7CRUPC7SchpGtaJnMLDnb2zqe7Muc+psFot+OG6rNj2JXX7i
BmIMAYdi6WDCwQVuOET9kkRET1igc0FcVyPvwv1iEJHhYjD3nZasymyhMl/ULqGlkTLBe0mDZ6VY
AgvH70yFNVe2gyU4nTlQOuFgIsXPZgFryoXIFZiTaSY9r2MVgUI0j2GGSRKsrWeiz2w+XiYRn3tz
C+XBI2R/4apHuVXg6Pyq21w5CSxbZGe4MQYshbUvM3JP4QA5gkEupZ+mQ1ZnCaHVrx4NvMb58KOG
Df9ZojW7knTNAxdqAgvCgjKIdK/aasBw991RInrlT/twnc6jPi7mjdvq6cJQ9f5HUHNiP1IK+6ku
SUfrKilor6gODdJ9mAiQW5ww+SRVRJOec99AJINgQc3zYCnQB5Jft+ajrNBHatTKqEl7KSLMKIoW
YBZR0RZdtLzS3DuBLdmnG4NP7kgdQqUhMVcB4k7pi7z+TAtusm879L9hFEQN4Tof2+LD1SRTf/hl
nfHnDCfe86RvzVHMjiPDSS5cQLwV8apIQkUSk/Lfm3mOwS+rLNyG/9qOAlX49dVowB54NrO+74ez
cnMrp5HEOiQSR8W3GXSocWhd+8tQGQw4aROviNG/OrOnXC8UzCC0lEyvDuoZdhrffHbJSQNGGEnd
tF1KLAHFs3pCs10Y7u1RvBHJFxh49hOOwIGashh/rArvxTJp/anGjE06EBDKe5aM3iDaM4eUJ/L4
U98mjos/tYklXZFwdeU7StxEyIDiWx86uMp/l1nhVj/whStRRPBijAy7o/IJoOKt8Uzf/NHkdg63
LKaxdqi1Uej71LvigEDK7YGMfM6uZssU5+H/gWeAdy2fRuEGkzmQOEKV7YOyMtM1kIpFA8RNZIZg
ynvnu8+myrHc5H+oYUncpQ2nIMCVEPmDO2RC6ne6D86bxG2H005C6HLFXKCR/HylZTpxXNOoa39M
H35P5HFIEBUuj6YwEGv1qpB0HY/x8qJz0+7mTXfjYc0voItQnurj3BuBbnEAO9Z6CsdfE5pvz7mu
gp2451+1wNn9QOD40Vcg0lF532t2hZJk9VyntaysDlTfyN5Jep0A4sHW4zWuSXjU+KL8M8Xu8w19
M0QEloVGhP2eERDnf6wuwnzCzk4Yjqzet7ZYUxOO3i2XL3gWQwC5r7IJcXz/ESLP0FCOyBAfoWs2
gmXUM+TCSNhj8/gfCYsyc18CCczdPUMIHam/U3iNzi9Ajky6+M3AS9/ctT/QpU0Ubckz+EZtETAN
xLX2My1GCFsdJgizZcr53RnNLI8yM5ybC72PCpDuGpLqj9o/DH7qhzSqOv23rPY0lSTzofI2plgN
0Tte3C9+lQYie0aGDE/i6M7Br5lploNT+F3M4JgZJaX7W9gwKCVvcrtxbpLlMbrsiPog+hnh39t3
5CfkL1mFUk7omPrPBGSVRTSZVeBfm5nrepzvOjp8Y1W3SuK9VLCGd7VrOyHhp+JETImTwRMqj7bO
XQlMTYOjEX2AAFWWfoXwW2hdPRYC6A9mcCQpCW1PaEKBMybA6P75Y5CVfMVOpSC4M5mmjuTBCFcH
Rgc4zbLO3dtMikSmJBB3MqL7jkXkj4ynH5LRTDpEBIAGSuJVFoO8wWluVqJJm6pMQj4trYSbxMkc
7E0Kf5Y8gvyZ8mIbxrFd3XDvvil2HOSZ+ZZfG5+Qsi2knXHs4yaV4+FkhElp3EFWQ4hbAqJbX3mk
zWmXxl/qAYJpJxxufxIKrjGXsxrgmHhgHk3gpjtffkjaWTwrU+Q6Gb0V1niCGIlwDewHXkRtedzK
vmwd4t9qnT8Zp2irIYHNX4KFcdgZnPMg44Xvb/CsPpIb2nHKH47VeuWPgXol+3aR7zNVk1JGkoXk
WMKnqyzpY+bXxmivvfFtKjVvtQWGA1iusmbhD+PFR4MJnuY9I5V2UMWHb5ULr+dHdDDHVTNK81zv
tFtx/YECXtu82jOMcqtR5vt2siF3iu0PmWxEPn1QeZl70BMknWbQ73ysuFzNst6Z2oiyiqhYnMy7
TI+Bygrfu4Ri6oiNqF2AKkJ9Zq4ZrCtZRED/0Dv3wMKFZCaaNg5ljclzCqX1QY9lcuLjMeDAYI9f
h/zP25UEtBYnXHXNersmFF4BT8/CI/6WtjBacZNQqcSLwRXrfPOp4w60QCUal7nNoYN9ez4u53+U
AoYxgfREhQfcLCdTb8tqVFDxHnr4xlz13zgyHFiA7mVMuHhOhi1E/+/yWNHKANFX4bbeCR7ZnKwP
fncCwoIcClenavtnKWrFYgxt4AnIw+vmoByRdOR4xp4Z0auhZTFEp2HG+YF0OTUCzThhGNKyrpgy
zowrdkNhS/P1WznGlH/E/+AooxWVkHkeoZI+LoMmcHeILHw6HpWAvm0qoRURB+yOnnQOVAkp9bSm
aikYIPO4GLoIpNnGK/eXmAIwXhA7dBNErruDYufyLMhUyTU/T+THsl+9oVK/cizmZybp3N3j77jN
xnFiiwPTURmu7eNsAUYzpeQ10zLtnEtfXN116fhjQbAxymH6D4kyVYyS8Kmk6SQF37ZibgmSNaTt
SJQf74ZDRKZINlmEir269FRHeK9ktBxNy/4TMy+qvoiMwLnl0aRfrQW/s3jiYR2ra3B30sYW9oC4
WXa2V1H0fcXDBQDLzlmsxFe/Nw7IrVwg+jq818z4lHW6G8Tez3pxMWJ73mef2EYBuHI/uIoEE7iP
YFthzQAksTGi0uFDsAc2nxRQM+2GQW1JFE7Ei5uFPgHPXDBdgHPPUrB4IdEdBnDl7gxsrHyPaNQm
k3p7akRn2ZO3O2r5X/siG2EHB4uJtMLCwhGi0T5c4u0L9h5cLrDn6B357LGDiKB4lby0ssZwa86m
/4y88ZrWeCE4Io9mDIwqJmCgY15VsDoMpP+EHGh/6fEJdU1v+EqqJKbx5367NrlC1QQpZTzXpNQf
D0F8N/w86p3SFTk1gt9CEetOk6mBWn/yt9YjH4XjjYE/wzd9hOzxdBuC3PD3tYflSCoRKeWeb9GR
i0ztPA23/5hnlgj25OsZHQA9ROX4K2BERrntSqrmPt26yn3kWfgcPrgQDELKiFuQSLAvTZQqsZLs
M51HOJbFhNN1JeU8dRZy/Q0E+ly7bPV7xmNC3lIkOetUqfHwwFwB5MxTssVgp33LOODOEZlaILv3
xUKwH/9dsKK+MriyZhJ1XoE4JMsikxvzFYmaNwQDsLT+oEGC1mkhkw29qjzFXh9BEIALF/EDWR1l
L8DC7GbjKM5+n4F96wWErIqK7p2txQWq/U+dp1iMCz0TOLmbmfutDp3YRkhf0PSxgKi08RBABDEe
WKcxVmTfE5prWvM0ZOzbwnXw8LUK16KG2pq2F0LrVTLjv75YkP0a0nrz30GBSOKS+SUmsif5ldU7
6bGYjgSgwZpBAeq+3azgmUtcq+LX8eZcj4LzeJ79TBoeLUo/hd0QIg6bIryhPCIaaIpp2wQ5WGJw
44vI1MaOFPPgs504gYiccIquWws/FwdQmWPe6dhxMyColhvAWwgKOILdBAc4jxbyl9Zf9wpFYIFy
Vy52KM5w11sKRGpbdqu5TMLe15/ZeF6qlqTzRnUCLxfwGyEysHBEkAa37aKOFZYx0tGlZT5usHi7
53Rogsa56ebQ/Mz3rAU5glc+Wylx1GAV/qPGpqmfqy3apyR9QBvtdNWv6sC7vR7sdYEmf/aVJEEL
dHkhtUVPLZ1YzFUQhXvGS+uU0lRZKq1rjy/0wGuQgbVV8JGqSpXV2bQ2RidHC5dCjzWj6yun5wEq
XrDIvKu+1m51TJAZZn2nZSGLhZDqU6qQMHipyl/wqbn2DiYxbWn5Y17wVCKleJz80N6cZtYB8GT/
8s5EnLDYE7cNr9SXCPqQEPOvqkk8R57bv9YLsHTYIz/PUzkR87z61rwVN1+LtuJCqo7WZFkHM4sk
7nzlnNygmoC8CvZMrLQynNLfmTcLFr/aj52CZPU2Uf47sLB0dw2UyeNuvy8pYg71rtyfTH2Ps2hO
ohqPedyDhBLu5JWE+sGNzfCsSqT8Wx4FyINYLXPPK27VZwhQk+psnIGO9IPVJ6UufwtHr7TunRds
U1VTAe5IoWU0hAl4X5dt7c3KW+rypAOE5VpeByaPk4oI9QhSfbpYWqtfWNgDfHg/jiw2pJRm4GeV
JV1iA7h6wa/EeljJmgbKOI2tXGQYdgKoTW5Dc+I2GQdsxnLkM26c9G9cokbsUuRrhtPxskik8h3N
FESo2ZpVBVsfDuPYGXzfaLE+kLVrtJwKNZiKN42xYGPp2euYDiAsjF7dxeGalhLO7nH1jvUX1ldP
+dEzrU/M8IrUwt8sTz+MbuKXMjGxUH9yoOizyHHFZmNwD+ruckHXeqzRC7aV3JBY43YWDbEJsINK
jORc6LSfxdRSoRTv6b3Jq4f8RGuseEzJc6g6IW3HmkHA3Ls1PZ0uOhqCFPrbDphwW9BWFa8JlVFa
NT/z/5xx0CbWxym2jwlhV9Cp7rIp1Gt3VxTHTXde7XJ28Dq9gwJ4Z5PROznUfY18pwhvp4v+w7aX
wBdijmuqh0IsT21huH8hqNqIswb/8Tgi5B5fnJEala+9TAMhQxXPMY+GADX7oIryU6KW2bl7oxKi
V13be/bWdGP34e577OmoAl7kOISypuzckGUbY0Ql/VmUQmpelk9ye8xgQvXpEapVXNilhuTJorTL
owcP5e/QwwVOXjMh0FOJgsjmj/vxrL//mLr0Hmcj9WADgHWpan/vX20SKRx6dn2EGCgU/z5SWuMm
jaFn+x4aAX/pTpoL1xbLBh/iV8U3vIe9VBPlq5aFuSlUDhHt7Vpy2MrCs9erqJ39vuLiAA/kp9e5
kbPmsSrVG7G811QVE+osm0Npa61MWyPESpMHDu4aeZP0uaJEwF/66aVPVPpzTA9fosmjUlibKuJ/
dYMZe7yc0dvyfMf1dHdONImhlpk7lsWdBMDRQUIHbUehxnYRJUNZ52aIb3pLk6w5MB4/Ku8xdOqp
R5kCPRtzeHc81/SLN6L9TMhWu9I5lwaSTjMM+7reTPFSpi0X+zO95b5VE4F7+7WfF1EiRseNI+wx
wVDuyqtH7UvwVWN5FAe2cG9gMRlxiq6xKGQfkD40XjP1Q3CBkFmUNVm2rPsr76dwWLB39v0EQMpi
IW0VCqH+C+52dM3SBmiqeVQQG1loT13u/d+MDobUkFahSgEYFT3SmKc2xddXEOQ37mvQKNXJ+9Rk
Ws5nUUM9xufSk6djRkDxz43bt8B/LGfG9srN1sOb2KnbrG1ykzrZjMaBt1WxMhXH1fmECmG1uRxM
5fQyyroCt3wUHDWBr7mb00GY2XnxQI7oRvAoHQ/0ey/Lb2kJDmzuOMXBkCxawMIHP+uRirPOhUNC
DxQan5W+bWCGgd5BQ4aq25bn7E/kupRnP5jOCxRm0I/yyDq/U/3ghUP4SHNOXKl9EVDz7gFZ7TQB
rVUYrp1ohAxrTgB/vBV33oHvFAvYxyPC+OHbsctmXG3Bf3xn49JZOtYuzT2amumrJ690kELpvUNs
YkuElpxuWG7rXx7S+uyn7pXHOmZq75ygLZi0/DgsJjiI/pycPcN6DIollj3kEUwKTItJ1uA5ztzb
sYO47w8XPf2V/VyBknRe05G3lMqNK5cZOYVaIdzMpjh2VL8iFGy9S3+kX501pcRGoRFlcZquat9K
e2ybyQDoHcfLwwr1RBnvvibE8fXXY0JnSKDX3yUBwSu4APkZ0U9tNV7DKAqVa2Ahghm348FYo2he
SLOTeB7pVeqRLvhlJ+NJnOf6RG9aHIawU6dMVZlY8SYlWxa1l8y7KhZ/SS3C9w4Q356LngIWRsbY
7/fZHmdoKtH6hfsoh+E50Djue4vgekwcxpVDeWCJui/wsI7r5cK0vY3YRhZpXAU/GUkQmmwMcbYr
sFvgwLxHbxH55g0ldYEOPj98kDGTbFCvJC9h3/5SFeO985snrOsVzPaxxDdpy19heb62HKUVrNF2
9uGkLADBzrJS3E4YTl8fNgiLO0G280y54dWTiNPCGxaue0MzpVuRf6cwzp82akoNBvUctOquKBrY
UgPSGJ/RJae4jr+r2jyUYhHmcFoVbeI8J8notERzP+pt96TgGyvj2TTQzQwSUF390Fwd0flrdrpN
s1jFxFJEJG6AFRjYygJZh9h4x/dgUQe0Wdfq3J+Q+KS7Jobu6JzUsTJUL8KXyDkHPaK+OlFUSYz8
nNpbt1B1UDUUlh6I+VPUQy3y4CyH76yvNSXvv0X7V5VF8D+xFCTliQva1P81vQLlNP0WcL0y9JO0
hYSOXBEtm7IGUp/RBZSQvncEFMuyrijijOy7qsqwjhnPVazBb76dispmoKcWJnoe+1UQhe67Qp6+
RkslCYjOeGmHoH4GhIzLRm3ZYHYK9HlxZkh428CCtD3R25OS/CyEnuSFHwR4WDRxNIq7FZYWZV75
EMwsfcsGxCkl0Ur65pAT9TLRY3rVohR8ebgm0nAmivjssmc2k6dlZ4AftYOKpCDWIPjgXQHDFzxX
6ZUBQoxF0slCjP6uWO53xBohFiN8/KJU7QqgiOFc/Q6pzlMVVOhahJ6uPJawAB2dBUz+HPWLwcR/
5aCeyjnrP7fqFS9OsCJrQY4ukZT/CwJZ66wbtXqAY9Siiux7qiEoht/khEQCuo1n8J3t8bz4ew4Y
misCXke0AWjQO3uvnxSG2uCWAfGmAKKbztBEbgVll0ljlAVmQIxQ/xFf+99bnEM31ZMLhCYXgG9t
8k6Y9HRS0PygXPjyTk+OLFrFmv4TX7IObm19etchm99gRCyJloHCoPYNVWsMk7nI2tiOxi2VaOaJ
/cDvhBvYI8tPBHU/gRXljvWP/w+30xO2ETmkrfaNYQ/6pkxSs64b6rSjpAdcbxrEYUdaVTYgfSg0
cM0YjhGV5DjfHcnibIAmpY30cqjtpNwLip17lgvyTfPmPK92AudU96tHMBIQ9cEdC7T0oPad33jg
XP7x3NhIgKOw8a5RBWUAaJPxpN6cuFmOOQHNU+VNl+w5BR/bEbnInPYu8QTxzEF0Iw//I2rw9g/E
2nsUgjPkkGdo6wmnJ9VnTL77QpTECnvrRUAqIgn601dSAoYBqU/BXAntqeE4QFSallapFZAo5ij/
kardVWwEYfPpF7usFdRB55vqYSOlOrurK8nd/stRv1lCiXbUX05c0+yNLtB/1HRWxxpPeiQyaosX
OFWJuKBd2uctJUOt/wDGYs4qNgjkQjyl+IU5bXr1aJCGLVHuzLrkYyhoi6H5OMrQx1oBYA4JLdt7
DouCVRsn11ggnY2Kb5AkCGMYRbVg0fQ5NRFY5UlOTXAco+oUwIVpge8n+9hD1APxpplvXNdcg62p
psISwW2DUnjO2DgOI7gS0gfO6YW4hs2fEkSTU4YKtgtWjHJF5AVnnVrh4Q5ziCGNNCHTbbZ6dkDR
jaBnOOYfAd/wCFNXCrk9R1mG5tivUL2IJ7afde9jD3fofAGovXEsktGNpPyQkJ9BM1+nDY7az1D2
nZ3+ZRmLIc+srFxVhVsOlvSHAGc12xbaxe/4UCQmHJuDNz0JDTB79i0ecKxNfd0uO8CHp6yJG5vS
/wIxDpD6qD6Tj4XA1PRNcxWQCCIRyT3MCwawkKr82dggz+NxyPOvIMCZGwZcyFUT0rTzqcl5xXzn
y4SiadqQTqDziaVm/tgxPsZyflKUkJFd67bM6hHej7gdhJer+JvTMRke5bGYG5/Qt8GuZTWSAgdX
ndC+DQcdJPfWOWPIrsXveiefgBTbWiL+/po4P0N6Beg2DhmeQEvYAMRIw4TgpoBghS0GTD4exd/V
gzygztEO6ovEv+botU9TU9Dk7pyODDNK01Uuk+aaGsW49BBchwFFxPKAnjjTKU9PUwBZTe4hhCXN
nHuXkrIHnvaR44B8g5ydNfQrVyi2AuVXHayAaobr9NlfhW+oU9K2wFalkggh0s/NUyhw20ZIXisQ
RSz7RiHNxxUy7bI7+5ZLJLrJBXLca34NYzrqNj97sUjejIeBtu8w5sYyhoMefRLsSq/2wazHgtom
FtuQefzgAzr5E8VEI7Cb6qf81JwJpWaoWO6FtpiQhotLPqhgkGP0rj4tNsY9Y955Zds8YyHo2/FR
Q6CoRKIhUC0NI6kWjEHzTCTSK21CPmRpg4Y3uRU6dKcKp27K11uLm7fxyoWwbXaf6SbVdtmQ1cD9
oHxZ3UiEcxT0pqi6KiazRg5aqQSEHzA3mlZ9X2sJ94WXsqBqF+pBbO2SfU6ZLpW8sk3mdsjghDST
Nd/XA/GGViF01jYpK7DY7mCRXf0DbpqtNne1NBR3V+w0lzHfbKXsKZ55lnsrZj24EXWMz0Gt3wwy
8Jd5hTKP+YsXEV0GRvR8T7V5KV+aSmIOH9HYiBI+kbZKIF4/A2s1ulCKrmxNo1Ly9RjzFUJVdhk7
opcwFV6ag7AVOzg+GmiCFnWlmdt/Bd80KJerCYcsrOV9LzA3KWqJH9nIniAn0wXT8Ud1rpbsA79f
WP6eeNbwEuI3S7eeMbCabIAXwXEutKbZmeVoPJOb9q0I6BmBBn1s3esNWz4H/k+w5ii/f4FoCPbE
sbVSgUZrOV3BOY8pbRvUZ++3tAImqhy1B0Ff0C5sPEotxm1i5fWVPO2Q3+jN0crXmmL1KWaFWMLP
Bh37IJK/H2MwUT0PRCrwdsnTOkzjTWhiCXCO5ZIoo2rbmeV7rYgFGnz9mXNxWjeO76LXcSfrj9VA
J71/UerAaNYkXRhjBO62waxKNsJhz4pMYpm+GOnGniq9djcMmVO1IUKkwcCT2ePKP1gQrW0tIcmR
4fpN9qRdrJtqW6yIjHRTfUozDDtyMPuB6LD2SfAfn6hTgKotrwJ0sFhNAnLptVZQGLikt/ssUtGo
bqP+dPtjOzO5jo/6ik91H0zs5lJiaC66BOUwwv46Xq76hUhjFqq6Bxn0nf9CajoUiOMBCfoEp0Y/
7Vjf2rGK8pWyriFX9mf8M+P6h0lMDgIuqbu3Z0BDUtfKMamSbQro1ifXcLwIEkdIivcBiZA6WW57
c0cy6EI8rasoRBbkiD1/JOJMAj4OXOo/JlSb5wrHG5D7vEIXY0Y6nE3x5x8g3c3k+6axX678A32i
3meAp+xYG57uP+nmL0Msd6RvLkiuiECPjWtE2VyqyYXwFBYdAS6Ji1O0WnAeSdXA5hfHf4N1EUJ4
hPfyeamtmZ9jTEDvmDW99AmjDPygJsq5LVvGa9HpkjT1FhKjsL17RzELXCYhiEIQq3j3gcWy2jok
/vorR/oWhAYoJl76BV+88caHvvYjxwkgePuB7hXvzIKyFJfzWajYoWA96wUWL7TAChi7YKIeDK7S
fHhXrbReE7sc/m7+G6U9bAIBDV6BVs0123kd28GR4U60uJDytkN0m7zx1ghj9mCdlzMFCL1owsPf
IrEwQgqYlvCAbHDIq13pjwPv4Xd5meu0w/78Og9B18/rlBLsTK0J/2nfRwozAfFV4u9q88+lTcKA
VPKPvYuGWbFYdF6ckkMSia1mDPz/yJb6WYj9joYyfHQG5opsdhiCKx9Fua48wInfLOcMpLFeRrx/
LcVi0YtSgCY53YqT3BjkoiP6dUs1DO3Y/tFc3dXhv6N1LObjnLsOQ1ZLeE2vslEsdh5UB9cM1X52
LFx9CpYDq9GRlnyv9XxV5V6+OwLZo2WNtguLQ6Adp6AjWLZWEVPQkfzs0v97nmbesdN51AFmqCS+
J+pNW1a6MeGhu4PhI/Hx//c14Jkzf/6D/Mghz4+WNEKypBPvP2RhenLD6Hrr0qIYR4AtnOw6b/U6
e6RNoLZmprvr8TSbOe7klhuzyhkwxn+1wxaWdGKpAlhz7uZgnVJhpo/VOYHSwnHobuBceEJIUnhx
jO0OzKxepAV0X+TyXO/rrg4Vc9f7Kiwcppn21o2TiY3ELccjdtg13OVoaOWmNuFXIETU/fkhXyXZ
yfv+dYUOBC9N7Ps9yoCvPnNiXTATF8u4CuPW0H+GA797qfekZyva0YOZtHe1ca+WVI7aBh9mzGEF
DnE5S4YldqKsjiOMuUW5hIVrQkEqbEs5SIkTSn18PUtqY5ZISFOeESRr5Jyq9R+pKesoD3BgF1eW
VdjudV4aFTbKo69436yXDDiVcacGw9y1rh3AsHKXHybk/xCodVuzmSgFfRgsR648i7/EjkwMnsT5
3hz6sOd8Tbw+DyfFpPFGSe6HRBIxA7bpGZMh0/fQqmcL6XquXmd1ti0LjUMbAr868ch4l7VUDTTM
iFZs/dr+v8GAUCNY8lfH+Cdr3RZUPx98VOvcQvw0B5zc2LO79ZuQYaiGn9Fa89JCUtDje+Efbdq1
PYBeErcF+iMZA16hGYMx0Ij44wPurxWzm1JvA0txphOBWJwGhs/TWbJ3o/oxvpgtdwWqCCb9EzZQ
0Uq5GwUea/1Fpag22FBnPEtkiKYUcAmCO362H3eZjFeaC2MSndCEpHGIgdNRXWBDii5HXC9y738I
6zIq8IDLDcvRvh/ACHouneZ8giG/ci2av49huHF/3qgxk9G2XakKqy0vTkoSPJrA8lrvucEHT2JU
FeM9EDDpa7eGXsqAPgzNnhTck1Oac1lq6tyRa+wAeGalr8HjfrjvDciCuMoOxFLRy6xjJ2KA3Vjf
mnKp3OosG/TFH8ICCsxNYv8NvctECyAh5uqgIfh7KCkBao+MenH5B3UaIeMZA/Xx8yTiYVZICgwq
c9rIWKyCahjerQvmz5Py/4e2w1Xca/xzrwDfpgsnskSlv/SCN69FDA8kdKGKSbiXC6kmrFDYaBT1
A8p5Z98+kzvfXXrBIhBWv8GjuSPHtECDXU110TjebCxsVetW4bKFAk4eKTqVDN+BbG3quW+/1UtY
BQHvXakpVADSNUAIDyBiMumm6f1HcTApnjVaAr7PXCuPPL7UEM2xwfqqcfs5tuPmudD0KrkYnhjQ
pp6ixUARhQmG1/8vu5KgFymOdqS0fIv1NVszb35NRE7A9LlrkJ/7+TZK6SorEm/03Bw4EeuZ86Ng
s1h9dpCix5nel+N2I8p1buy0ABZYDt6OVs8qphJwFPhwKwnh8sqd/6by+xo41BYdQc/OZdlEMpJt
cUk7/iqirsTnTekZLY/gmOke23Ovhb8GruUoQcJjL2TLdAB69YpuHrkeTzmwYF5OT2aotmmeNzQ+
A0WDZ0oLmVr9XZsW7Dq60gy9ke1oo9giT/+PcvyjshyaoQ7LISQ8/oPzIbhDlXKp/LUZoPF01IOm
fqgriWvaq0bxOfx5ksJIGocZZfY9cmIHXfN0heGUu35ig6FcwtDaFFwgoxZdfXgx/04YV5chrzIz
z6oYAgBNnjvHOKTW6mTqlIBY9HqiBv0ai2Sr3scB3p2nOWiTP1FfNiNqfVBhxcTkBygcqGEajEFz
Pqj1zDgWVQTf/CiHyniutg0XMPj8w2sNR/CEIWq0/XDlkztfHLWuoMgJ+qKzOIzzdmXcy3emRBJO
dHeB7sFigDCOzFdI17IJ8oFX9dsDw8BI+qDbIuwOPQxL+4s0v2Q0p/u39yXr5cfNzm0vCpxf57rL
jIIBSr0j98y4fP7HeEg20NCHlFzddEZhZYQaWAJ6h4yuYHAgGoZWUrazaflQne66xCLQKND+Gn/d
zUjQmS+SlEIka2mpP6C0QgAJu8enQ094dIX9uma8PIp9D4oMd7BLs1U+wrNfVjPpkUPa9QGaznVJ
fCd6gOV2zjXKIEE7ocO2PE1YG2TXCyw1AiSHnPZ+1b2bZANd5Qe3GSejMQEooFRjGFZphSs8LZ+0
G30/qPNOCR0uoS9YQLdchIaEPK8r/5U8e/UQZKmNCpdDyRCUVJkgYXJj1Qb9MzG54gLDWCsyaF1/
ToMX4W/t2X4WMyzXkEKeBidWpLghtNRgq3X9wnEQ6SlB9qud8z0oLOGVKCo3UeJZWG7vrvymkz2m
BLJ8lxtvBQ16q1q/Ldmn1UuOIPETYvZH/LN6DqjYmCbDScosRtdzxJ2VTqJvKbhZVDJz0XAlbZCj
wfMcipd8luHYvG8hzGqNaaL6hxCsoHEqotTz5MQQshDhPFRfV3sS1N7/7x4cmDqmz3ZB0KGRRQID
813nQV1e1kD0Qwv3Ur9wb3wAC08dO3iMCvf7QQrSKZ2vf9iMv6uqOQoEvvlBVPhu164sl9H8iQMj
cWzGxGK8WPqR4zqwiEjx6pkQhiXvMGbARR/nZXaEzosocWp8VnPu8lGyBDG2Iu9yH39lo9fRqBoz
DzA2gnmUh54m475FMB6wL1P0S8GxqZsQkVWToXM7I9BxKF1B1cep1xHwTnLm1qfneTu4FzDblwnS
pg7OMexDwVOBbRYzqJdclgo/mC9CAxYWdrq95ock2FCFdKt7oP9HXLkKvzy4YaH0hm6Ygo8uu+W7
yJ0wVU/PYqS5ym3bZ1ejmkmm70dHkPB9QTlJVSCfRxStDaZl85R/dynsikAepbVmKG2duE5/kb3F
3QVKS93FfDa1PEKpWtO3ARa0LfXmAZydVrB1dAjFQSGksDqRK3wHGuV/iskF6rufDbxcceM8Wv3b
05QR6EjfLA7kcfdyQQjQpq7TwUgehE/XzdhPqZ5R3S/lNH61HGl4g4ofxhoo7WQQI2b8LInyP7mu
YZQy2eKa5l9JIQmua9NaFbv8iQMWEoiyqYuOAiHJ+u7V8Kn3RUKH+UoyO8y0+eKEDWIyX3Xw/UUj
yZrQvJJmwVVqcCpdQn6RNKgLZSG9EhJqZsiXzOeEwr4XPl2hlU+pZVsfYXuXyB/aY1ImvKh4QHxA
N+V2OWDm1lxC9gEWQRQ2cY4P8AY3KupnQfXR1/PzmGz/5XeFfvUUb7a7sVLMDmOVBGpKknmYGKBR
zSvopQ9U3sXO7tlD75PGX4ECMuyHpl0bClkR9nYzpMG0CsjKv3RoaQ4/ML4VAlG55ycaJl1hNRMa
TUzKhC/51TLnRDLHzsvz1kDVTEXagS53CT7kmPNEGOCmk2awIIDNvcJrIHdu33Jnyw9pZPmFicOP
FopfaEnlGBIKPFMmpPa9Tb2WsYopcABdrohPkEM9b4OqQSPc47VJsJRx2mSfEn/qaR09GMACxnd5
tNhubwCzZi/CU0g9dvP8cwIj9zN5CNe4ktg8z6xln4Roxj6CGY9lJqYuc+JSWlGL/JA/ylkbvG8R
RDZQ2wLxMQ9dEAcE9Cv+lRPq0oVQ0XzgJ5Pcbi6fW8cYRV2/Adgf6g+Qn7lQD1/17X0OmYnS11K2
Jkvvy0/Uy/+RraedeFOzg2Q7H09/jQX4j2KHdQM9uV5FlcP3n5qEI4CigbjBqTZmeXrOFWcn3Euh
fq5ozpdCZRokrAVRqhSw52o0IDRO155gDx7icmGQZfcw/c//PU9P97RSfu381ETyyuJ0D28vuhrq
5ayJHNDkRGn5W0SyYXG4/B9yqZxyfiI7pmmX9dS78hv69/6ckmZ1hZCruLmj/Zy9Qd4in5g/xMxP
WcdGEnBSYuxOqe9QOa0kFvIFKk9tjohPVbuU524i+hZQo0DZhy2ITk5ElKknMKtgISSkhYlcf29G
/2vigVpFwtkL3RwbB9x+3j+Udejm+tRGGrdQ2nW+8aOC7yEKs0MoPjnSy2PefdxQQpO1tp5wFJye
ssSE82f1OPqGYGTJOZ5e2SqyPAWILPURg7he8QFW4HuNYgnid2RFdC+JC58I7GuCuSqNHI1DxFju
2jffXfvheg4o7my7FUoXUZ8mqJcA7uGB9t4OQCPkFs1YK0WXW5m99PKRwPvBO6qptkfhhqUiwBEA
/AJUdxhIb64sbE6Y/buNRa7YyyxKRPHYH0uym+jyCBXCfBGPONoEK0qYsKRmuO2qg1wXNk8BzmXb
UqNDWhyR4EF01pmbZYIZT6YAn1pLQBDncO/o/dBWFBf1cjoeVfdoAiIN5mUSOdsXkbQOvLj8i1y7
5IFwTmRoo4H42i7lrnDJ+772HrT99o0qDNEVLlBYcPPfmukqGVlcKPAg+tcuaBom2RlHjzl0NAAD
GIKYXaX8+e+qx2E9pTcSjsYv+XV6hiMkkHVZiTCLp7NCpPZJI/osjoPwYUO9X7QSKLaGvQx72G1z
HRQvrdW0f8HX9eWJo8zpsamI0KwCU6kc7tcDbsE24ZhFHIK1tU6Hy9RmulGcp/tTNJcqV9kDzjql
q1B1hbMK/b92QSr7y5RX9O9GvD6l+Xuiwaa3l3g+orO1tTJHucc/SIbZH51Auz0YfHSfAxQFWeJ4
xei/aP8ZnDcQoL31UBZ6etKZIelKg/4y8Hrs+sv2F2t6CpNxacIq43U6lRsqqYPn6831qvJO+UeR
HlcsB60pd+H+gKSNzE6DvVXfmmWLJehzOy2DrK2nI9alCZdqdGYHJI6x5lPoQAu55AWzDZxEpnXL
ubNRUq+aC/7UykbXyqPQD8JmLZPJp4CjFEhll/cEcJAkdGMbHj0FaV+obISG9XCiHuVJoIk8x8GJ
92t+5oTjqqs7TVmo1h7MZTT4EEF1Vn7rrSNw09kOiMOgb1P0TeFz9wpWRLtX3cA+LqyeG1sGO7IU
d+npEcgsQfHo8nvS0AQBRCFo/yANcsBcjuD52Vc9WdsASvHzhQNLoSs0pIi6Sya5G6sKxql6uYhV
zju9ZIoh+gVo9Z5hfjNAYyyMT0bhBzTd8mC/bXJNWGGabShO3acO8GGILvJazc2FVZ8sGa3D0r8/
6PzoA3m0qgBzaa4b9hFTDzTBhpTkxoNfkQrWR1qbda1eZewGPPbCOzQgdUQeTmW4c8HSQGIo5hUO
URc/adDTHZpISNhH6DWpP5YdUizEMJ36p6+u0J0orgkLTdZB/N5sLJ5XEsGqTgxB2z1dqDbKIF6m
TGGtKhDvumYl2zbE/vySfvFotX9r7RhjbidsmxavBP40ydAGQqlEShTwa7USmumMmJRk3XJESsDz
ceEa1BfEfs8A/7Ax/A4Rohom8Xp8UelB1GfuJrX+74wVy0lOfoWRQ1iWJ63v9gsYcB6xJAQSs41U
tpmbEADkAwA5J6xRs8ycBYwRZ2fL+kxCJiwnw3ljzkQxxKmSZgdiOy5HNmSHJNfn9xS8mRBi2wVy
jYL7c4WA6FfUYdkhDivVARz1iE+oYrxt9Vk6gvBjBbiaYUVvq4jJHf5cU70iXBJtnXaws35lE3VK
hj9cKmv6lGByon3tFoENQ4TJB9zEVCtgcbUjdqbkn3JmWlwSCOz9ieBxiaQC2NB2hDDcFYLs0h/J
uSnMWK2HrEY3lK1pJUsAhxrzlnxZ/EwgeHU8+KKQVkbo6lFsUS1fPATVyMTvbGcu5n5cYgB2qW44
KisZ3cy3oVLPMoQhQcDd7EI4rpMluFx6rFcgVZgZk19eUm/g9A304d7YsJfQ6Ki8hwccLIffEAtv
ctbaZUJ9I+7st3I0g5Qkrm4Xi7TnhyTR0ASJEyBFcpykHsX2GpJkERyfhyfCYzFLnEVy+d3O8Z1P
onFdjSYmgGQsj6jB+AXDma7xBp97R4ZZbyOgMFc4S/S3WLMT4ZeUwaYN0e7Sn9qEIxOLRn3ADiin
juz0aYlmC91AJ4f4FSzXRPctMyi8P3yZO1iwVuhBZtpqGFPtY38+ttWen2dCTvU0l6hnNwN5BiWG
N8FXvdDDT23JTT5Qo+K21/6X0D53b8TpIW5zazAHiSAA49hpUxdjsSBc5JAbm6wPOJzzliD3GYWL
+zUYaJvrc4jtf/yzG51/AFRlOXGV21Sfw8Yc3CBGYvdN09xfAZ75FxwFwYaTOhXoftkYftFtrKFU
ievLSXdL9iyyiupJFj+5m21XKFR+Dfiz5x426Lp4bpTCVsIEJ6EZI+53kObjl64hDYqt0xbPXdQY
ROPmQLEsxs+Th979ioTgE6I+LOMotKcBSffNT1We0fWdBR6zfNj1AoIRvv2su1Zs5Rg8ROWouqs0
yXXPoMaCce1u3km90f8yBEp7xbCmEBiALQrwVR3GaWQRfQguqIVb6JCQy0JicGaFN86YBzJVc4In
D4d5277EKqUO8TYI2s7hQmXjfajuJatGvjxwEs6DrRB47hIZs3XD5wD5bPrqrWE9/BDTPxGqTl67
JAv+KUsfL0uJL/clC1X5A6nib5aLevf+1FwOCnHhyV6IWnBqVpT/YjGUdrHD6foyRXnI9G3vaUJ/
td4M17U2fJmGANK5BjM8DbCm0JT7fd2lyYfOgTeuk5FQ7xhgpOYc2Rg7AW8obvZuvNYUoDq4EyjW
kFGUu5sCYZ2SB2ywSoXjPo6GTDzlD7wmvr+YAPqf4SNg8biHPDSXP/yE6zbNRHER0v92cq4XaY/m
y1trZhlaqoTu4zBwNXM0OxecdpulXLfBtFPk+48vRLLtwlvTr8oNrC/W8rxxmJF/M1UxWULcp3gZ
kIYbK5cIWaUFq62uCYuwJ2IDFpxfUJta6/YUgNaP2pcWtv/bD+BBEb9E4HXRxex5UCf+4XQkAng6
KI19qoXjrKWTmMtBCKZkRCA1ONdI4YU32Isdw3TZB6zOenasnr7K/++tw2m3Iif7fpv0Pzu0s75H
EhH5BXeHt+XdU2r5G2wj4E0DjR8rrr4Ud8SzQACM5cNycOYBwD7QUph5vPlhh7Qo4tF9yAHl1vXS
70ug7leyZUvHiTo5FDKvk6QZgdxBc4hf7WrOt1C0+Zi500OriG5gEiVRIQ5dWTIo1V7qvPloFExY
Gv93H12LS7FPf30dGmmcP//Xf518wHFZIObhqgqZrQu044rKq+FxKg/pereiIkzyb+CqcndU63X8
ALCc4Kvb4LGo/tkZYAI/m84BlvRMEE9f2xMj80gbHwKMB5wpmAgv5Y7heiYv20sjXBD9DbGHky+Y
GS2iEugX051G8VvWtllKRWuurCzy6MC/+WbfhFA24RBPhC/BOFyMDGuJ6WVW6aw4BXB6iYOWZPLb
KSuTv2RcGFamsgP2BlLiF4KUSwFSSviGt+yP03sia1KZeahWaIfCpuTkcm3ST09truCqyUCZmjro
rB7Ka3yf4wLFNAXHF0cbbPmtR73Sm3fri+lr+pBxd5QWPXZ6npd6NhWCG7XReT8N1IGfY/DqVKmz
qlAeDmeB5wwHAfdQGlKZkr6Jx3sTCm78zCW5E1/QrPnh3LA2DdduUEYURDrNbSQAgQHi3hKkLOu0
TL1u/9MurhVpvaOvR6eAoRr+t8ValGJC6fdJvYKhwWfTQMb4tFhe4JBoTjd7VccQwJB2QWNiISzz
h77+rXPr57rmTLWq+MbT2MVZi6Z3alZ54k8OwxBSsSyybdjXZs0Wm6EOvXZSXkeGM5Iy1Qt62z5T
qOzBs7olzEjbESv0VM4WMORoC9KKHtJqrFFFzOS+8IBn8wylpRPwbxztOPdUZO4WsugUATmP8wt/
Up1KBPj41zx2R/W/zkqpHR7eY+y5cfcikZVhrBFda643wi2Rqg5mCd3Dj1CW6OkorAQB8tScz1Tc
4Kbr/qbo938g83y//s/dkCAtfvM10G4wrf+WGkQLd0cjpfJh/T+DM5vP4Oj+CHWrZixLOKL8RVLF
q/fPV+UwaKtelxS7kw10YE7hoGOpeUKOaMB8Zzk5JJS+A2WbACdDUlmrrzsT/mFr7YMinMH7RBko
bfsuDIb+3XrSvGAnzvMPQ7LlJx+jwjl8S6PLuP4osRFxzy/Gp9AB/S422cgHqg4w0X8B/jhd4zun
JQ2h24k2F44y6TFa6qMRk/mh4FRpxeASf2pgyQtippV66ZmRUSI8nLXFc3yFljpELtLGWLrA6YMc
ZaYpLwnC3GenRPwkfXPl26/HiFtpIAle9Y0FB8VjWfbrkkN3/HEBanRqQnLnZNSwAwPCPqzZlhSO
Tyy+ifr0BMRQkmCbTMbjO+9BDZrR3aMIxRca2wkELAvZf2trnOgDtwp5poWd1IRz519QMGgJ/Hyb
BE5C+COFlElS8VUNqxFJlbqGb91fiBLBkpP0mzLjf+bmmLntll6A02sF30f4tdkjSOB7P7Tzo20k
MEoTuqrhTYHsJGwCX7xY2E4V+1gCIqS5K6QrbV48yZDDwUizsxBV6235ESFlUZh0KAvbr3iRRuhq
PhHe2LgRjrDA0XgzIr+R3uNzMg3AIRLoqVTfm5jNafN/ldmCA+dbGJX6oGrRYfOw+xAwbhxYxhVU
cCrPvbUeeOxzmixIx2Jh5wBkHMVAXuBcELxfyZwyfKHs765iZT7m44Dh7nYdj4Nc++HnEu8I4cAb
ZcC9sEqkYKzT5wTNWSVhV7/gMKQ7G4NtmjiRdzMBI011waH/Vg1Byj22WGe79ZW9e9oeB01JqwBK
H5Ah/bXw10aMh9w7EyzM6jkyvP/O9pF6WIEypsCZqARnNfnQmVlDa1DtV0xsBo9thnMQiPt4S1O0
o2poSZ94N9fEB8nvjgxuC20/8TFaJHHFNZNr7kpN7X3q2Q5+Y//lZ9rOJiDQM4s0kZkZ2dPjdTJP
TBHjjekg2tJrU49JF/Y+SHXJACrLJpKsN2gFkfCTPaCWvlJRDZCZGiuFwGo+s/SYval35lFWQH0g
Khrpmu3r+C0zlY3Z/FVcPLZuSzguuqXm2KArguoCEQ3nzrFwkjEaMsW3GRnQsMdjk4ua/cas37JM
NKhuXmo2cv7zTF21zda+ykAVG2BLCtzIlqKHcVcM5PMWd/vJs7EJPDvU6/TFMGUeyGwazhFLImJq
zbDr0PcDpVnpwovQOZ8fV4SfgiCaRjlB0Nh4RX0hEhfnCk0LJ5a4giIPDO23Q8pWaGuPWGG9e6p8
GiWYL2wnU6irfXcmhOQuMsnTVH3nkxNTTBdig/aZgKCDnupc8ZYKVRl4bDPoPHXIyD6xFJvJPRUA
JjrHXCCDk0q/5HZ/03VAQS/jiUfnwkIukkqzsVEOjyRfUVAKKIIZJS530eHNeZ1fLbcQGIHAHbAm
kbiPVdnlVnFbiB1fKgJYCUbWkRf0W3NWToOMQ9//IMAZelbICb0Vj9zn3Nt5lfEp5na3KyzQa9mp
Hn8cTLw0WgmhGBFuL4/W4NIcsoRDNUmEfSGv4+GUfsKmKQxL4pqc+X5peO6XWZMC83GNWMjo8j/2
t274w/4CK/i4v+rMXFpdAMBTa+VP+a8C9aJA5qrFDqDBTvhCPh5KWXu+5IUVO+T/La1fW7nn4Pcu
Fc+UXO7Fa6UVVOhfMGusDOW+0LLodbPJex70hxc2RYjuu9gUbf9nqvp3NCzdi1yU/Rbr27ena4RS
0QfhZeId8sr/iRtfgfJyKEs5XN4s2a0GTJHPD8SyAmfF5f2aB+h1LwAsBezKFnk7I/o/jCLPfbmL
uO8Mc/iQJNkYKZLEoYC1LFdIb3lyMTLfcgkzcuodSIpOB7Im/Oi+0FwlTq4P3vRloubdlVMqxj8m
0ffc51zNMxwCWyqsTguJE9udrLQc1EyoveK/xe+XdqoK0CPdY2mpX97o++fkxhyVzCQgrDOT3cbH
ejI8RUzR+IoQzA2GLrEA91Tdg97tyJjFRI/0LO89GJmf2YN4qC6fH+najDt8h9yzC+tT82/ozNaK
T4ZmFL7o7nFEum+iQnJnxnky9dwfFJ2igGOO0d0RyvTRj+vz0yxsqBHqd9svvKgMA/iqzccc8Bhb
DtHVUWgJygx/arvaHBlIxznKrcG2ERlNze7Vy7K+9eWxb+gKLjyn/eqByPk44DtKsFIWY/ZvL79i
wdNVf5nZx2FFDu7NpyCXvyutu5aYdskXal2DZ30wuJwfr/2SC8/Fu8sZKR740iAEYiPUr1XrECOV
tmAsjdSW/WmuLhd/4CV/MvJlGuJnspTyJJi1EDQ662cZfD4kNDtoDY2rPbIw1aAwdwy+BxnRRax/
rfjaUZj++UhXXNlJybe9lIS+t5GpsQgEYBf+WJyhGarPwnk9zSOn2E/UIhoO/1cIxyEM8LgXEWrX
zbyTiIe5uLT3RuMuFRVvBCJ/ofl5hEG7Zh3i5fxWhW6FUH8KwEf1gbAbPJhzdJNCGEwCIe6nbce1
13OO4gQyKlSTjLxDumloQKsO9pKT1a6EwKFL2PnxF17WiDoQi2YNvyXi4ehhPTkQ24qS1z8Oz63B
kCR4OqSCasdVRnZ4lx4xHCgrzn/L1ePQbjsgYSg0E6B55GHuq3PuzCup4YU+pKYsUNfLl6nW8OYj
oFJxV9Y47i6/3yCZXfIITZz/4+zhgql1gTQQhNw8bzd2NKApMBCdl29OHZH62JMwRMg1xIFv9uPG
y6f1J3nmuw3zbejNYu8hcCsNgnSO+FJsSSqTilhqYaKJx6Fh7UzJtmSREZLvqMC61HZoPnUX3LUA
ehMT8p4P8KcR3fQAKBMBsXwqfYKqFZroWQHlmO2yRBs6DzgfxZXoJBt9LncD3D5aKqz3dNB+PyKt
N4xcMHl5G6E/LwLfS3oHO4X/epeoUINTLj+Q02L7j1PBkRibrUsf00MF8V2u82juQegtc1JeqISO
x0gd8c8XCn+otzQ50+jMeRnlofr7yTf5PPi0sSSaKHS+TYG9SsDW+K99Cqn7+VjRmSoJcRvNAe4k
Y8hH2k4WB6OlrlAHuJ65xOBt66jVxQgZQpMu8mIR06uEqr4HMFGitIVg3s5q9f7f4E3Nz6PU0UdX
0KLSbOXR/zn4WBQovX2A/JEmh2KJTwkr5+GwCkvAtPZQh3QueQMn73I94IyTJHN3A9dWB1CJvgy/
IQjwTDcLycyzby4kg7BPYsIivpeSRygSWGNRkOKp+Wod3aqpkO936BCo/i/zIkuTk1Pcx4b6jqn3
Rti6GFgjMDySZXz8LT8iErkr1egM4Y335tN5dDDUxmk5N9ZzhNHVcp8fgpMaoXGzchKDaQVs9bO9
N0AGZiMGObltBcu7C8WANe1IYeqyRxi8E4KheKU4895RMlmST91IfM2vhf8dmWP4QOott5EqUTNf
VZUwGls9aNcGqduBDMUPRUN4Q+WbKYjGhWNkj8xR1ty1mLjieME+mhsQAa9Hg60+Ycp4KrZKz6WF
bzPzSLj51vhkftvGPNpT4g8WDya7pOcbT2MutzTX/w+CYcOLYWCplKYQvfTm5xFb9YM13bkVek0n
Dy4IjY7TC/ovfdFvgRpUgpN31v+pWn+XC4PCl/EaRpR9upIMjRPclSgbdxoDAyzzihpoXnzJ3yBI
yKr5SvrwCKvfPEVFhtht452/KKRzgZTiZHCPXYbnIuu8DXRm3R6wwQBRBCp3OO2mA6yaDjrRwEke
ZV1KVs+8EMriiOi8PwjBb1nij6ETD8vZOvnJoeYLy1lmLMGW/jd30wMY4B5j5hxgRHLBoHrkQBl9
JyFvrqoIdH+rYnmnmK/L5iHRPNZlMXajzSf2ec1nHr5DXcN0YXF9vWsaRjN6vSAkrjd9mOZuIi90
0/rXPrJ4dPVlGQhSki+SUQr3puYkLiS01h8rZPTGchVtjBPEE7sLCAgxnVPOVTBK8+02oQCaO7SD
ZvfKTLNoH03QTouJz/SdgC44fTLyUvJWJTl7RIbGYgh3VdypLysYP44lPv8Eh/gD3tC+eflGVEQk
EIhv7U/TtxS9Ga1hRLjh2bftM5+XLRdQzuXTPhQTzEir9FopCv6XR2r7IInhyQAPC9irvpPJu51I
vgM5+2lT+MMn7Ix13twvjVlCzQdPt34Vw2Ho5um+9tbnjY5DCh9Xo8wYfKGAERs3OLyBilFvUwW/
lG9+O7L8CqqZMDrw1GpbW6CJlgxliraqNcDD+jrFavncCqec5C19WgvVvsl8L4C50yeoSUz3zkBE
AV6yRce7UpY+2j+F6C7xnmV0fqmcFDHuZqEEjCziWuzlbxAbkrMhBMlb7K9h+3Hk4sdkFnVFQImH
8pOJS4e2n8SzRyfDphOw1nlP9sx3K3QdmYYDRnFzShS2AhhLzERZYqldiditOFiA0wsRJ8+WQ7F7
x34/SKrF8kUijYMhc0o21jAqYutkZeUYzta7AgYrobENKKaP/mifsvlVBwBYmgXf3BHZWZV0RZY2
sbP9uAxjv4g9Krp0Z9pCO7Z+SYV7/vjito7et4cyTJWlycqvCQ1qlq4NJeEyzrJzgj3nrg3vyXBh
isjtCB9jeLHp1uzA7xyx6e+9klZ8gClV+UI/2XymsddvHXa1+SMnsV6hYuA9wtlH00YeFfPL7uNJ
y417Jj8aWvwegOSRVLhrXFAlTi9STjm1/UaoMCrs4902lR8SArsF3kthuOmJkgxrAb9VdRuY6EiA
SjDjqC9ac/3tbZbvsZX1Q8LUJkMGgyFxzwf9CDwlEXe5n5GsaQqGG0Ij+fDl8WwOssHl4r2sQTne
K6Pn80i1bQ6K9rVO49lAf2gh/nkhFA7R7umWpDB8JgKrQFxVTw8cVI1JKjUOkF02o/lM0IIQG8yC
2sLYSRdtVwdpWNRX5BVmrEI5eDsm01MVFbgxLhXxDZfhPpYBdiss6lPd9pSTKIR6FKId/uyv4NTi
xf1wbpvXxtRNVwiRjWF2exCqU/V0sQ7cGYkv/RjjR2bDfDU2JKXP7IWyI2fU2dqPFTQctM/igFH8
idScFZpgno6SY0H4s+GNkpeYk4KttBCSRPIgsxKiwT/1OpWz24ytDh7L4DF6fkNkDM5hkIU63cjP
WzObdHgsz2KTKCuaLqr5fyhNeIoZ+AHCMioyYHChnxnIi7zoYWKH97P/R7t55XmbJTvMDhFML/CT
sPdave1RPVdghL4BeiqCYFu+ZjXZK5zu7+xtRn+pqGU8XK0h3sqO5yHuB9lbbHkaIVWbkLYfymVg
SbogXSCbAAn966C2trFctrMTdWJ7b3gpj4HG2wR+hk2EtDS0KyzmhZUG/+7FkbCMDjbxdXNDh+ih
JA7ud5JkxnxXMDZZd+msCGCOK0t23OE3j7RHmMzE7S+scIIEulBYtWJzX62cRzdK8AkQAMGOSk33
d1np5H/6upl2P2bRkVpxFNhtBNpv7jp0wi2GkmqkoDZph44UIQcvFbSND8UsJb8WV7bGirjP+CrW
y2yILOS/2vXViauEPyCCHtNruQwihMYwKjhQCrnW2/qOahXi2AbPTHLjlnEXnQO0L55VDccSbZOu
JGS0/KD1ZUNTK08EWvoK97GOSxE6R24Q+fi2D/A/dQtUTI149g76ehXY3DK88DYp4VvkiiRZX/1f
Q0GWqLvnmi+6BrWgLtm84qvOmoxRhJNv92cP2tYXCAdkaZKINwmhuKi+Dl3CS2as43+dnMCV8qN2
X4/oMuVm3o7dVCApUPupTgu6AkQyWSK6Tn1ixq/KaRD8o+4GZgGoGh5/03YSNbLqnlPhbGcOftJy
GjCB5nPzC3Y8baV4ZITL2x32MbUmu4aDTKjjQzAat/wfE2nZi1zujhYrqXykdJxyhQpj9jFXgIMN
1itguJdyNsNejz7D5hDjVh+QiMqeviRTzYGbSuN0msgArNK5s94BaGN2KdW6RhtCM84CK3mpm5w6
4AWy0kY1fH9Ae5FeMFBgf3QlXEgftORD2HWH5voDH8WXHJc3AmWNUI0lIckc146xOui2fMe5LYNG
8L4ES9HDS5/egYVyuI+WzG7Rg9ZvSrZuVN/juRBFw2y0HlvhXXvHyIGYn6tyiz6j1nRia7ADK7Dq
awn0KjNvjrwgQ4NBzT8xp/a6gint+vHZcozSqbytdxHVdA0c3mw3hZk6WG6HEJe8sJESGV4ZeRpu
O224sG5XuDmFu779dZ+IJcHRAdO6o4zL0w2NKzCfnNSanCZgTvMasbDv8i2i3MsPJcetaB9lopP6
nKWqiIoJ2SuPGj7/J2/+el8JLVMt4Qpw5SmLScGra93uVvB9Q1cv2HgnrQXiy4c40Y5zGZVeLFOK
2RqTwM/i2y/5QakN7Sli0JAx63/s2k9r7g6/6YSxQ+fel1ItElkbfXXc2ROW+2cc0/y+8snBJdE7
LZiPSmW29BWAnVRXUYtGyyy4psHXuBWmWQTPuBDFZbbEuaqNbKNA4pDPEQ8T1/BGSYdBxnxzFKtf
j2reLNbPjKJ+TbqlyyBZcl5T2lQ/3nwQXFP7B/PmmAt19QvrsjBa8I7vxuu+Arvr++B4GjtSHmTA
sGTazTYJYmnKjAZHEh2BpoS6/zSPGCMoquSlddkqddfG/htDZNYfA541eaIt9LnKbf/OAfrMzf5H
txp/q9bCjRmdAyG1ThNRD3VIw2TYzNooyKKHo3loWNuxVm6M78oo9iL9EkOnWMRJ0+Lf2iogoifd
iiZWpjhhtYD03k+zOluLaZoNGfXgqP1S0ghTyHuHozUmtsJyMsTYncE96HVwWl/L8f0tXZC/+OrM
u32LkaZEUQdPZILZILf/mlWxEzSdPmyPFkTcJ7QI18SppuxEeDHvEltwkH5l0n8pdQR8DJZvN82l
yk25/FFM12RCS1taBUspeh+F1Be4GeTTwsQxsNH8JBHh0kiPbHiwIrcoL8BLAXuy6htx4HGIHWzN
ixROvP/+QTMfpWTbDemG6vXBkQzUqWIcUCGbYFSk0k96xwMvtwXUhdgU6ohCb2fFLkjKw1qlScv2
UVtYd22qfUth+mtrEk/c+JWbJgt5FGJSl0xhxRtPhhkr5nbjDUy6uPN/+4//wsXPHKSWS7lMnJFO
tcHHmqu9vGYX8rXJ9uKB/mz7HmfOC5zXuOpABnxoKCYmDuEcxtba5MfBNPbc9F2EXhjdL7+tfZLV
lS/s/EF6ZMJlIAnHsdnzVOVFbSLZELt9ExpEFZIWuq2yLp3scUlcJgdqbuo9mm/vS2y3DpYGFp3s
Y48bzM42Yq99mizEsKVlRV07PrrWGu7tTcUkSCLC9KNfPQ7yHa//ipPkzciw+yN1GRt5h88vp2xJ
IJyr0stxjOy9RhhNgFGJPL8Jsv8/j7o5XxtC90mweQlOPMw9sn1l18CwhAoeI0T01B2Vwy/MJ5/x
5FMJa78BtGBPfxrX7U1W83+dQ1lFVD2507Xcf/3BJESoHGAfIu97CKJWO8KH2hjReGlH5F1OT9A9
cu/LZWfV4FUaxko+ePzUUSuKSRVxlSmlNmwy5g1Q4AoQebHTVGvXyB9/8S6W7nyiMTUq1TTpHhgP
RuBCH/s8sJign7GXyEpuD8ObNqvppf6ORjkYctcC/ruVWQUE0rjhN+7yKpSfYiyTiCh7AGRw3E2k
MQHDfREsOTaiRZIyBk26myJRhnwFXdyBf81bd4vRI/QuVYHCBNqwcI/pELy3c/S8LAdLazt+wV0n
bWweRLDSDlnakVspmNaMilYC5s/Wf8218s+xNdIQOrg5wHG12V/lB5jo6qMYZ3QrDHMLGoUrVke1
G472h4F/g4OVJM8Gdz27yBNQQZ5O5W3fwl6rUVotCeVH1smDgzL4Qwcb4/PMJftpCkDJlOlkvoM2
fCC9bIQc4yL6NOZYsLlEYJ72s7mQzXNp345tbjZ25N9616ojSeQ+sULHduia693Csxx/3W2NWqEI
V8mzt1HLu4QrQiBxoUn5DNW58DFR/b/5DRrmksRks5gmffY6DIV29fe1rJgkIhPf6GCkYEaKnNwx
8CCJNvqvodn77K/TNJ4MEXVxqA5BAx77yFawRdvpPRCdxZa+R6nQYM+2R9R6hQBK4N6+t96UJ3eZ
SQsq8G3wv5ib3rXVHaBWqYk1nucSI22bt9cbzaooU0XEN5er+agnuSbl4KtsK/X4T/x5EPCxEaWm
yFIAKFjBlZ6P8CIXxo795oVgXapiI+oFSBphPjNHTuh1DeAZ5RILUt87DDcZL+68f4s0NUCcPDqs
HKO7jk58+F+4npJLBdhImTS89S/MZrYduQHhKMK+KrV+lYF+w/AfoX9aWzuT2X1jrX+FhiduVKO1
uWMYn3Ha+UmkiF9Ub8zLu4vIYL3n/1n+hOZqTOOJrrlv4bJbBDZJV+ap8HPRDFKxGre5pv8H7YP8
gr1SoBDoXvNjsJVX4Kq6G02vGSbzs2SSeJi4D8abqcgtB7BCASHmdqdxitj+t7CMWZE2ZY6IIMqb
GtINCKYxYxzcmsQdu4u64+i0qoNp+DJX+go6TuQB38ehuOorYKAC6s9getezVBPfj1F+Or6Dnug5
8tIdHOKCvvPczCgQ52xTF+BSjD7EQeHN3pKPVRd1TJEBMRjt1opiBS6MeRbGbJxdPdMysVPWvhb3
aWu3vVEAmKUTQID2zjDRfciTBBb3BAGT1jW+EIk0Ozc4opRT5/k7P7uV10tXg4VhbxdwavpHuc8w
CPqaDnO7oTKfcHBnHrDGW+xgZFw5Oqf9FXo4BdiYHXf+LSbY0B1KvbG3umR0WvqGi0C4kRXLQCNN
6g64Rxk2DZd3wV7MjnVEgcafFz8DGGdYsXaMDnG6ojl8ItpktFXKmJdgfbAOwq3ePnRSO/duG+TM
2upvtglkoueo4lVwugpWHcGGc/pt4kqtOmgBSaBd46IZROTZw4Ve3ngCKgNiaKkHHODUsBkYCwOF
by3RAVa2aAFn+UZ2b/3LN98FcdYidQ/W5G1svG5coif8LUnS9J6ebsZxo1S4U6QPeZzCJjIkD1C3
0qbO7zASs6I2jItG1h8+WDc1Hz3woPmf4w448QBqImtq8gn5nKOGWIGAT7DgYhhmr/n23WWusEMN
tNKdVls4OJriu193FhK3gg4/lL6PLnCE2Jomxv3Kt+15FamIyHjEcU9LgC3TfPxeeZ3icdm8Q4XF
ppGfzDKgW2qHU9w7LUnkypA9Md5JMJATy0aJtJ5zC3tXPQ+sptq3ce5SHvhTjnMg8+U6Ark9dQ9Z
Maschk0CCjte4DpQwxd68PsB8YbVwmMN4P7+ZfmNjWW8BGViyEm7TLOX0P2VM125ETDbHx+EHZJD
9HO1pRgexpa7633Bxj8iXomdRbqIpeRBGL/l+sojRi+mFE2Jry+SOI3qIyrAVRoyFrHTHMmrBR6q
Q3H7T6xgh/sZPaHcMbHCg8Wu/rHRkiwvIub65tGP4V8qzl8rV6XD9XuSvtYqlI2I8oyGb7ja7MXJ
Gx9NtTx5Aou6dU87frP+gPkRwARW0uMz6MwNw6FCAWp1Bwv8fsFM0Z83mjy0tpH28PYsc03gJm7t
6YcT9JVQsOsYVS3i6QkZrJKnunGJCb16rKD9vPq0ZWIycYu+x16x2do++W6TwO4zM9VLZhsGOYau
z/KycFj6ajN+ycXOWeiZFX2Xkk8Lz7T10hTV8va+aGTxc0MZUKW8+yohuoOMiMxL5BPETwMVJ9ky
7VS0XS6sWU+NxBw6wOXUnHnCIh0OJZYFY7UrMgC8wT5OoXgZcwN7iERkQr/NYjgLZFPiFxYLbdwq
emFpbZEu/Xz2MGklifj6yNGLTESBSHuiX22e3j6Xy2HAWXF11bxZZkZ6i1BrHGYyYPEpCkHYLIds
QZJ69J/7gaQc2nLKyvHFluqzmowpH5HZDXiP4b9NDbR98H5iVRqtWBcWJ74sVoSaUpoWp/iMIdNE
X02jcN+avrJZ/57uUPTos/e1G4RNOMBhbmwnSIfeGuowDNl5dP7d0CkUVZ8LQT4MfkOnDwBW4scH
7GyzPl8PmFyjlkczpMAwTdXEp+fA6IH1/C0Ok33MLcEn9wJyDpqK6XuExSatl5WYL7Y4mf/oqGEY
ZukZkMILVMmuYCpVCtW6xE5St4nuUnBrpnwFhGTHvG4OvRHfP5mvxRG+5YWBGKp49VJvagwNPw5C
GOlx4Huyj2d5X7/+S7OZi41dy6Ow3ev1jLoLDPnNFodB3by5lnEN9QnxZmZmadzEBfx1F0xxi0WF
rtDH/1vVp1zCVKyO7VCSvzst9mtW/SiFlcobCBDb2lYDwO5R3c5x94TNJFmyeLEZj2NIIReXz16d
aVXH3Hu/5rcJu2Vw4Rs6df4O0C/sotAh/EjMicvWf13ArCwKxulFNKDbymi2sG7FzJKANgw8qieM
OzVagtwjVXTNc2zMpGChVvKH14MhhuxEitoIOVo/hrEPBG7FIxoaC3L1ARxro5RsSrVgUBvAKbKn
LN7Rm/JgS7B9Exp4Kz15N6B2WfGq4S5i+7GStQecmOrQyLMSjA1Xe47jIcpLRsllxPnU6u9g2cPk
1caKoOp9x+cVk55nI/vAE2NGVv0Uxb0GA7pR+9CbYZ90P7oaK+AeduNJZo18X0vQRb58obOgr0nF
Yd0dEQEJsLMHGzMA9C4KHO3U7c+26P+A7AeTnRjNd9J+NTlY5oOViyrL4VtVaGD2znS5gvtdUuqq
L9kCUqUAaV52kjVRj6jKM2blmXXrpp/CP2BLdb4Zaye8A9/Fh5lHlaNVzERT5f19moXCbE+H7EKV
qlKsUDy64dHdvrZLQQMV6j9Kw+A31sOl7CFqEN6Sav8/YU5xCTKASwXmRsrKEzHBw5SIbwL5Wpcq
e5dgM1r8WUwl1VAqUwS1g5YoTyrhJmTUYYSjMciLgC/uF6OaiNRxrKVphfeOlW3K/odX7fvR8Ura
l3BORw8TjAw3arLrUH6HZaE8Ksl0121cbbLB3EQaXhQY0Ci6zD7RtuuVgakZIrWZcWj6x0E5B64/
nxr+efh3+kqxb9GxHmne9pTURnip5207HR9ItnEqBPDbkNGt3QLPBSOGsGVzS5Db/5r0C45au71H
3VGsmwlbaZK1SJoGK5TRJALMj0nK+mdMFYxWdZRtvsjwRwTPUWqy4qcvEXP29Shyyw8jaCK43cHY
C7CC5zToceuxBEJyEcpNvsfYzXPfUfw8z6EXfCkFSYC1rnMfKhTCRLC+/YnHkh5JkT6ZH9EasL9N
+766HKcEAmKsjl8OFRunRTcOuXm5aw2K4w35X4cuPZXmhYr0MIIkjdogmjrE2IZjLoA0l1Fhal7z
qduIQLQh6WxlyE2LXUIQDeblIeG7VUmpIUwsVnIGjw0goRA7ZJM2Tk+pKZNUqTHlehQAxGfCnO5+
tWS4wB6gh/IW7d2aIB1DTQXPrgXMKiOvDhhfnsOjtTskp7FqOozqJkrkNMjIBtB0bqsKqD1QdUem
sADJQGIOfNyWCSYmGOc+MyNnJcThpxyIA7xumVOHlnyrHhZtpXFYdf125PZcEHQ5CNSdm0glScVC
q38ArcPL9Xx2/g3nyUSmGkWMhqh0f9BcnBIQrfsP5OvsePmMXHaM2Pqpvq/nW5dXUpwHFoRSkQrd
F9ocCRhKPdHnrc6GxmRT2vZwNUEU/w83jtp/cs6kQPA4drcbuWBJ9+SVOnkYsXuBvJQL4OMS3Ice
qGEuIhKxt+U7o3dPcWX+P1Wks6Cd4pIWam7+OHKgNumXCGknOQ32YS4rv5Bdj2myzt1cCXEDIzpy
1Zd2HSa5xs+O9Vqp3kHpSFAV6Ro5EfaefbYJic90qvRPzCIqPtV15lPyO2GpCvBXx3+UJFBIZTXV
we0kgQAuDJIvtR6XlxixNt0Rl9at7pfITTT4TuuXPM1XkT5+IrZl8tAVRYWv/0pZl/X467ES2SE4
cI0xzK0KRKNpIstaB+osnLAnzpH8lRC3NeMRs7ACm/axBjJcEXUrbhJUt5Y3u70jhd/sZa0AduwQ
1jskgKw/KuDWuI/+9PhI0rN74zFDX2Ta2pMvxcWyw1n+e/jrA3Y4aF59NquBnyIqsplLmyPtleyv
m3RZoPNzL4O+muH2QBw/pg/tw+MDc6mgvdkJ4R7XujEdnMCaQ/k058eOm5Dq3WQ5XjIK3D7ANpDa
lBXMeegBxIiFKxUI/BMWeC4M+ELpTLB8i4FK6bQ+TYRmdKyoSiOhom4IJ1hPQb8GDvQRSLumOQjD
ed1EkrD6eKeo6Ptjh/gUfBaCZiEaKiXSfOzdHLbq+GxglpFL0hOIyIEaLHXlbERxh5MFle0gdonZ
TZgTJRVKJtbRQQRJNuKh0CTJs8dczDLTIUOM+cTou4fh2FgeJTzNrP23zRoh0jImTQqcEm0c+h+a
AnRPPoK9DawfN5l0Wwch/XEGPb7QAcvksQOS8C61a2Z3t+l3bB65Mq3Adta92wKJxOQa5Eitqy2U
WkkCJM9PuY9PtU57JVMfXoSzkZMkNFYg43Q9wzbATjeWDsiroRmkRXLc9q90d0eBevKZIVy1zEEN
ZWKsyfRVe4vXNUdgyZfuzN/5CppkdRVrS+T5zcIsGyyajO9C/1hZPDMAkjIlJRbIGtN6GcHp6Lfj
ok4CkHWD6alGrxhIH7W/HzqyvKC4k1Uv1Y3uKtvxQ2KDkz4jX/yaUcbDclq7FbJYUYtkvst+w5AF
dJax9k7NVzTPWzWymOe9mHl8ZaXSO5MKhDb9xP1BYpe+0NtDvVS299QxFgTOnWIYgAif1jgMatiD
HRAJrgXqgB0TAmsMI9cNjYHcejm65UnyjRGw/lnfUZDdfQKFx2AgDW1FgEZvWG1mtmyPAfgBbFQs
1X7s8kbcJ+LNM/MZwkxLTL/feCyTkoOVgO3p34KXXPYH5A7O0TpDPTzgZoXjnCfg9jD2MjhazE0A
hUq9lVp/g/U6M0ELDP8LPhxmYMDHKW/RxRVdO5B4SMgNpO/XklByoPUwY/14PQ09vohoAqYXu2k4
YSZKOvi0K1AAn+rPI9r/PbM4BQwct6wXyhUm7SPHZ4ByzlHMODhqscmVTtCi5nAX8be57lKGyklL
9ohGihlExLORim/TEKUJyv2hMDWR4MIsp02S/fXdYwKpThvW/FiE3y4LeGbe7vT6J9SmnIF5zqZM
Ofde8KwzmZSKTNFWhJWszRflV4l6GgYL/bwQKrQzX8b/rxYrfmfbUPhUO2+8FP2EABQmoBOe3X3h
PF3DAYlub8J1WORJEuard90TPnSdG1sypHiMFw+qWPLDhLBuRa67O9cnQn+b1e7ceE6x246xcqMi
8k5mL0wvHUuBixV+n0YOid+GFBeaXX3g24MOk8koij3jmc21By5jjf8xJ9Nm3EtEDCm3A2iBLwCq
0voMWb2s/JDaekDrfDOhGg3XPxaHQ7UDFuhQmo9uW0EkaJBEQ2txoOoaYYDSbsO/3/wZkKwGkyoU
2KnFBVdRckN0XDCd/xxsmNLcosBMg1aJKKEvzyyHjvBy3wEAicDWgjGw8zpf/rGgnnxSO1Y8cHMN
/fQrVAD5mOAnx4OOJwWn1prr+dw+/zlWh4+9skHVv7uPe4HhDFD682lwvGvw3lqlGvee6X9Dq7P9
BkztBwz8PTvHAD01N0Y4fvoZTIaCanbIKF6TXRjPpSmlqo+mbzz9hr5kNJqEy8j2AOIIfE3eBfXf
c+3jEvbanYUTajMTNUzN2AUoF834teVlyVkl/vL4LJ7z+OUn6BSsjlmSFdxxwhzry2Kcywmg5RsC
PQ8973z22lbZxc2KSsQomqYVg1xwz/77NDktveQv7B4u/jiKJSZnZCKMoimllSGGsIQiQPaAEjWz
tVw3op9BaltvcNFi5NGHszCERRWup537C9601EK8o6LuxKviodW8LHJY7fVtnV4TvCZ795h/2K0W
mBXKJu/k6zzXXTrkWE0Z5YvBkMMfaV4PsSoYm2WVuhi0TquoJEsZnC5VkXA7WMRYeOdRywoQXXe5
Q2Ke9eDm3/XCHG+INtBAffSixpH+xheIpeHBgz6XQrPiTygryjHGsifig9sbZK6881yMzHSFjvBG
GPL/bwUIHYn78JTKsfTPx4sQUUjxdreg5/8EemTERR4S02LWWtog8E8hFOS87tmEbWpMM4xaxr7C
WVUUGU1ZT/2MwkdkndnKmgEAGafrE6geZKfxkWzwq6e8i3oz594LZhnz68fFWG6Ua+JJveERFdwT
hVrZaj4t796yHmN0G9Luhdyn34BMz5f/clV8/3q8FqbmmPNSfxv8awejr5jpkQhgAO9jPodwNQRi
HgEmu82sFEZrG7O0GkB9xBZnJPyyi0/7rXm+AYPg2JUWGYLMFZcQP4dmKtIenIm8G1L77xp32iEe
x5ImKD/p9gyWKpd+j5awcjfOO6WtSujNKKulTfpHQuFtWyCMD9UCuo4cSNhqe7pGsZrGP7F6cBOs
v0z9e3c3KaCkNQLZmAijscw0D+uIseIfE817n50mrd0oqqTovn5OO1A5UWQmryG1SL5v3+SZc60P
URXYEDs7PttRaAAdFK1rRQ3AfYwbC4P+irQ9DlQPxNn941UNK0V5uSfB05t/akN5xv4Igm/cuR2C
IvzPpqvTZrx4mxebYxrE/NtFbTx0VG/j6sQev/AEmvgnhVrElhZCnlhWcAYTZk8P18SWoZZZKVJB
HfLetpxWytWk23rgifWID8DC/cnWaubsFv9pS3Pk6UC/Alr+kKBqh0IGGvNxIIsjpI2OUMney/Ln
cq9yJGDXPGk0ETXoTGbGPn5CnhG2BDndN7WN0tLKcXu0M0xAytGNgqtD/XKTVrB0nrQpB/ASaPXR
QQCjJy2OiGC4BBpDSwg5T+U80jZ/QjTEiuaX/FgHa1asNfnYd/Bnp51Z0CfeIrhKtlNl8RMSwDQk
3QM6A8Et9vqiLa4sR1Q9263e7xYS5POPH0FdCY8zgLFhssfVhSmZPIqu7z0TL6gpDuTaPiu2/tKN
7snNdWrCDxsXzQpcAAYJrOz5a+RIp15swGUWc1gyn43n+kADKOeYMZ9qirI88gqNsk6EoZ24+ipl
+6D3hYnuiXjOM/OgQlRGDZ4fHThRuNN2n3oV8l+EbOFYL5Ip6v4boxWDLUMVn70MA4WiwuJP1F+E
Xlrv8lQHTovQYGTt7OqWldTF8cSWteGiJBsislwscl8sgZvzi1L3rTDF5iEStyqkJUcTBlwYapR2
t6k2tkhGcmuALsD5TqKt8evZxalrgCWqq3trCg6J+NoTyrvovrjr3XSYCnYiJTcpkPwHCCu+FrlO
8frp9wnw9Ht/OmvktKTfkNGUiWwi+XzHNWz8/Ef8rKUqv3O9rOJBlGbN5jGewbfem0y6eqzyKrEV
XjPSRMql5LNSw8y1fRTQxCAS6aYhGXspdn2HKkODz8J6Wr3Gwvl+FLBfCbOECzWkywFMXJL++8Vv
5wJMU9cDWRZq8t7+Iv6gX4Df5yB9SeO0dum0qwEmR+R9TK44tvlR1as+pAa63VvlV0thp1SCXXT/
Nqs5o5+sWCKp86nxkpmI3jRCKkwBuSKk9WSF2hguq/d6kyoBrZCrArXpvKlguZhQXdpTqmvzlYDi
lH8X50LnMWOn9kmk8QvFQPagMc2r7x65phb5A1Old8n7iS0hH40xfL0IklxGLXBTsu+DP6BS/7O4
wFXaEPMw+fToSbopRE6XK6WlGeA7eC7oIBEPtfOBcQp4ePZ2aHmxQU3Pw7dFH3hMuDgJ2AAcO5ED
FzkC/tEh8Gpm89dv9NyyM3FQyW0yHlykwYsCOmYF98HeZv/xfs3S7irZARfOMwwOaoSZrB/aYyKo
5/GDtN/GvjdgD64TBbORnwiXGqLM6lJ3qObmeRGz3f00P6U+b2D3SRpXNXWenXavRxyPNiSWDAez
s6E5GIwKF7cEKNiXru4Fbi5c/os0w/myUevQEkjIgSqna4jFYVh4wopHXcdTeThlCUStP57oESPL
ZL1nENAZ7lIj478XZhjHHzmYF2GKVBwaAxIWJ4svSauGYxvvHTc5BgXj92Bq+PrO6gXi4waucUYU
f9BXjYsFIZabxUSYuRDd6zqxh7Q14CW+j5bjOkKZaMnPtdZA40BosOAWEcaUtvhuthWENjFiru3k
J+9Ws7etOB6N16rcpAaWHJ1OzZNsPOJWuxYkvw+9ejY9amLC9IE4BagkeUJPEfWs+W/C60fyQHnL
FAyE9aKWGXM23Zcx+E213VWn+hQ5e7bdHsk8W9h4blysKojXOW18hnA8mNyAU0sfUmP6wYft1iRQ
5uQ9ujbFYAIyV6SUNaXmrJfC4rAjz+x/wjetcaumJ2W5gvZv6NdAB2d5y98D8mcE4Tg8K7Wf1eTH
VLobZ0IC9E93wHmTU+Vs7UC36+/MvT041btfyx6TxMQixpsMJLjnGd6b1mFB+TQ50HTcUhWdore+
WuzHVne0PTN9O2IFRuGntetmvl7XwcUTSC6Ut5tJ1RWD0vvaCkX4WdCOF3jYBe15XtJcemKKUr9r
nH+L3GQOePJv2Gi+Cwg7tHE8xmCumnUVz3hxI98LckRWLkXXkpKcflE6MZBnxbzDYz1Sdhfr0akf
juDaoMZG3GdsIAuFEvKHNho8B4lGpQPAZx7a+vvJa+7T9Oa01XeR90rhnOmNMEj7i0bawPkvw5nH
3KNMzKeVIA3Mw505CeEY4eQZBwVhJ8AS7PsplveHAdqSRVWLEw5++i2PHUKxnUUkao/o73U55AGU
JaENqopf6Q2XWjmC3TTXJ5NdQ+l+E3FJoTDSEdSaYYnL2ixF9AoHS6W5r5ba7bm6E1m9NZDwyA0U
JIdJpj8BAhNaZNpKhmPzZCdUeUVkFOW6kJ5h0h2lZzNNV4+eMGQF7WvbwiXEVQsHA037sT3o+SNV
h9GYo34M6Dppo6bpyWiWg8gz+LkWyN2FXptQlKKmnm+MQhJNNrHlea0jm9R+kCaxh+qr37zS0KHC
IFXSwRmkVLDKQbFHavYKKWJPnX9TXgQoJcPH4WWwaYxhIG8wgYO+UyR506K/Kcs633tneypBvGmz
sdW6Of1RJSJooDGTIXdn+gZQwoH+/T/C5ox6oL6a5OjfSliCuwjRG3lxkKt7HLvGe7I2OKgbYq1j
0dh4ToYsv8kxCYynMy9L3oUBgHRTj7HKYxUnVa8wPtgrugtQh0qhTo/mK7kdnHY8NDx0pYgDYT+l
Faqfeae5gdS/CMwvtzKoGPoiAPrpdBVauSxzOQXCPog659/eZbr2/DbzzozLxFUKpXbSUY/tFa9K
jT4NDv+o2ODji6ydlL3glvJUwgZqTu5v7Offr1+8xuHMwvtiQaV10YFhIy1Yqi3lLBl0uwKaY2G/
EfSrgM8WMTwRrcTdWZmv1QfqTLnE7STrA5QmrOyPcJsj5sLsBt7toxfS9AWuXFByX1TH+ofKbSBs
vo64eDeM0x2AXT+JmlfnmfoasXNmBH0S4mx9VT5kRB9se9migcTbCXFlCnJm1lEJsekOSRhx8ARP
PTZyd6NNNy7gC8cn8VTEAApoOCszThzwjDy89TkW95OS0hUoOHvviMk8V8JBun8SX3+5scqQMjVP
R+ZykcA8M9EMqbhHkVeBbGx9lqMCPDGltinI9VjTN6GS6PIYrvsf9+iTJ0uUEJ6aVRIq6cCtLqkq
nmQeNon9lvTwgtt5e2jJ8kI4KA4kGUQVh6kRfZxQ6Z125IuGSy+xw2zMKuHQ3RoMF0yKd3RMqrrJ
LHZJl2Esqc7a5CzRrp5cwKY5kh93lhdxiANVKx8H5OceReykCnN3Br2Pl/QyAi90qz7QBLavGs4z
n8TvROT6y6M6rO/1IiluMa2xIsTQUxxsNz88GOn5FjcIBTDFux4T/a7jIIKxkA0KmxcVfc7lbcHV
JC7YSKczou8TR1ZlCndbeMoTPvsRvtpqwUESo4+gMV8WfZlYse9FgTpr5iIbqBljOphL3np5d6kK
kSsNiVE0tSGSPsAtCtkHn5yMTMXaOO8wy6xGMBh9w3xiK/QxI/huQwvSov5e1FI641oqHGMIFE6G
vbNAv2pGJyX2Su2xu+VmIVk20GNYR6c3dNKcDx0upKfWgc4RAW6t6lRN+0pEYuZx+8aBoMekF1aa
MUcIUHEAN7VLWiwo8UaapmRJroC0MpLx1blLYRNsTBbh0tAyErBJSQNhlc7C2qTB8Vap2xDojVQv
LPttMpxMKeS0kwxWZby2YTNYDpyB443SoZ755e9UmGsrB/QxI5LMSJJiGAXLnsDsfxG2o3G/PMhJ
ZJh1WMdB2fZJCei2KAYVx8182SRc9NEZEzCT4/JQenB9vvq5ZKdV+Qpj0sjiNT9NFd+l4xnw9lCH
ayo8WCElpmn9Om2fLcIGUpegF1O1ENS/ISq13+ERH0FFbqpBzdyJNURklEa/txTd53PAApSyYGPQ
y4s7irgbSwFCrDPxFqr+hE5q+hm02ZFGYIBhlHdKDSA9gEHFSwpznb+usSRoc86FTDz93W3Ui89d
bdpjWPrC4R0eIoFVXpqdEeTVA9FWIEa3UkLephHZ7CW3s70la8DqOhzVsPWwTi9qlBYoZ8PCrs/o
P3rnEjA17BrhlKzd30BLfSUYBs8lBw5zi7phYFI1uwKqFz9TMS0ZLPOna+uDUyRaetayQoO3ea60
Li2AAkeIOLyzbul9t09nWP7bCBxwNvevgoJ2I7RZdRieFohB1RrtcYd58HYFis6gQ3IZoSrvjR7m
gavlwqsvG+UwLMQ7C33kaOU67CqJYuEtMBh6Si946l2vohrxa48r2bP57TAidTQ2inqvj0ghZ3KM
89ak58D2yvq6dLLm0Xnaif8OXJqEbyaT5ZNeTN0itKWQ30s5IdG9e2zAFFhp+dpaI0zfPXxYXOuF
AF3mVXvbsB7+in0dx60ZY8kHK0ePeioRyjaGFnTvrwVExGZteUkD8A5X7klpqkftiE65/PF8YXs6
owRFqtiZYzdILctbGQOYHYy1oZ9wfkKpW/B9deXCMgElKRD0ZiKF4YnW7lQ7ZUN0nhPp9psSlH1n
6UrJOH3Vbv5clP7EBv+yCxy92/gB5EXdohYR5usrgWfa16kFXDWZcP7jBYU7kUn1BSgkDaGgqgIy
dSvkaGSnxLX138wIhKLsYtVAVOR8Rm0qtQqt4nUfEGnRhBphlpYRJ4wJMwtzOYXHzNMZsCisEche
mezBbePB9Pjo0t5B3/AivAIP4ex1Crq/QzHAymLM4zw/az5B8J9UV36wMtFDu/l4HAUPUSz3HUuU
ekiSvl1hEMSVMf1RVp8rC74Xb6vZNllM1RS/0GttUMkiS1DbYMR83BIl60M9Abd6HyW+fDAORe/y
mcjZ83mc6BwZ6y/2WBT51D7CYsmKrQ1T/fHGpQw6vZuVbRjOG0i1/7SDVaXfDzaUm4en5ON5YMOu
UXwG9nxkJ8daiG2xQRWsGy9KVpFc9Xqsh7AaNLef4CP6/7KWwpdd/D028o4SAaXEYyUAw+z8c+7D
eVsY9YxtCy/yPZLWbaDuFNL/Q69qZbDqkMofLAq46FupW7MmKHI967VGtGP9c1wwqYss4VeJQ0LV
3mmI3qDldIgJ0CoU3EnCGSd7HJfM5inGan7KksI+tiBcYZZ/HmNYit5/VMmBwRN1JvsR8AmKGeU6
XSmXMxmG9l4YWS1WTkxNHUE04gX+9OSVuHHu0e5ec1gmSB8f7A6xuegH+2b9zfFJplAv8BfwaxpV
6K29gifCV/xZErn1oIztmgLOnX0HtD0byvpfsasw41H4goCi7fFLRsKIJ9N/j77aFi27BY+DK/EI
AKZDRSLCPM+s4I2GU4v+xE4AX22HpAhmNCukmpolSRRNGzeZ+x88sFjYI6OM2YcS/QorOeqE2l8F
7x307XiGb5tuoiJqUKy7DcH1Wf01SWFOGYL1FWUuqr8uC25XM6wpbXaUYREG+Z2Ffze5UbfwUkFX
7a+3xdmoizQ/+78MKb3ZD1X6RTE8rxCC46i87Pk24OQSlDV23eEoJna3PF9ppBppls9Nr9zyCvbl
i2ke8KrfsZ3OUxHNvZ8HFY6d4I/OKbYK3Vjyf5quR7zkyTYLYSImIvjE31zpZPCihrVnQrix4z6Q
D3isbmN/+qxTm7fbtV2U4BLNdpKP6glijKQ/QnmmyadFwuem5lLI2/PR1B5H+Q289nT7wKB0qoVa
kbmc498qPxUOvukYkBkYppZb+FP2yhbHtCcbdgmrl1BmLrxxtwJwaEZw+P9NHzf4k8Wwnl+YGptH
FWtANJ9Jg/ZsVsROXGTSbBXIenwEJ47PFoIW06LUzBoKHzRrSzzauTIECvm9tjFE0/orIdg/sTWB
c5/Isu/XTWSFxMahIZlbrrYODVvjHewhG+lTLlhT86JEG+FpHEW2/xju+nUYLbwHD88YvmYB72FG
kEb4hr38ONvFBHRhrgxYWH2rShsUL3C8U9rBFB5NjNnZ3huMoxdeZ11CxOek/B0A66t3s/yIwY2y
pkY4Bq/AAOBe6QRw1vztdaEt/pl+kVtC+f91zs9MEPKgSmEyfNY8AxIafCXZkCJBjct2tk7FZPZA
l2OERsLiCxIenPDmrmLX3yk2MpE7inIzEdtDiQhD43nmsUMSwXvA1QGxyc/+uw/EAEV/MO6uqECY
O6c2ujymDoQuh2+4pBvfcd5NPIS8nPaisqgQj+FfMaFiMf39F3HllT7n+cYYMIlY+6+9tF2rxvPq
RLtQLZBgUhF8Cvg7o5xqkZ5iOLijspvhAP0g9sXGEhCmgpGEBc0k+P7MWHH8KsDaD7/f7GQ+/odJ
KcFiF//LvOO4E7XJk3YxoG/A+cPUQwtzXbUIK4sHzHW8FXfnCdKGJ9MYxGtVvZG8z9AaTWPHlaZA
dJ/94cwcDkBqJIl1gQ/1fAQHSbPQKSJybDumdHwC5uvI5+XAPZryKqgBU6Hu5/U+GtKsqTg0GZx5
fxHcDPWqgxVz3u9T1EFJKEiQaiRgwBsTqKktb9flYSUenWNXzEV5TFZ6ncKks/UcSL6JbTM1m/om
t58NG9ZIKuSEAR7vHMkzt47TGaMzJ1imhPRfzoD7+eNdlvVYeUITDz8unzKPMjuCyAZoQsrC1cme
bhicNWQ1Q3agAssWw+zExT2+ZfxOvPgZhxunf+iT04k2IIe46NzmRt/82aY3KfseR+pVCcCb66+D
XRIYKGrRr15RrCEpVML9z8GWCxqlyaWyHjlc7kTDe0SUbdYlkqro2FWykVL6KJwJRolGbVSrf+gE
MicfqHeuRq0dMgS6/7G7m9BpGIL7kw7GLrZZXEf1AFc0mLVcemrmCoWhBm81TgQLVon5QUgkKkD9
/zvv2kdSCQDlJDiIApPiWvmAN5KhNtR4bNNTDQcnhqMVbXx4wAyHucw1IC3WVVM8CDyQ5mPDWvd1
mpKtf1ctXP8MVJYMKXPJlsOg0Bmw7GjORYd/Qb2Un9vNXreISCZPGIFdvQOrdRKibQl97FgIzLeS
nD8m9T+hxNK7DA5ZvrGpUWiW0quj0Ttx0pqUh7SNeZhndhF1PqkJGxZIgAZ0kaaInP0XH56ff657
ljrL9ucdnJ3UvQWveepX03AYbL6SID40EbTOV6QHMO0hVGL5UK2aA32kSbv71S18s7iR0qcDASND
cuj1e24VfdTzYWJbVT3N+X9yoEXauYfaGZ41Z2tk85W/1RKOFRrTt7kHQaW62ZN6ubPCAPTlw2H9
gYoM/PysggBuWmRPP+Zip7iOfkxqFYw4Esw3x1oNeWIv/oYSlosTUCziY/W6ZmVUiMUWIFEEyQJt
SRGPmzuTbckisuxUhz+RDLBHpj6bB41rj9vtSpZZ5PDqfH0OkBqdVtqcul3PX/TmD+K2qQjEnk0+
QGDmPhE5a6aaQLfj9rwrIDOf9DQMIzacpoCuIG/ABMrDvQIP5Ete3w/bjLaA41QOgUJ4qqB6QNZI
M9Xnd+qk23ePK4oBrkulluA12zsr1NJBnOyVDyfGEZ0kHLqNTZVkI8aA/J4MI/DvMXkz82OaSFQJ
D6FRaOfeT0mMuoWwjDOPJqz9aPOwfmF5KpC1XOfma2icGnDtPq26fJlleXxj3+LWwxmu2gQYp670
zgKUzw1rQBpyRP5uRgggZHbEXRhb0ZAlfaVmhLw9QPbpEHxxNE2edyIwvKQRpaJnVwSEjnZWFbJL
WFXjA0boCj4CwMV+SUDqqzbopDo8fr0LN2R45pZmAZ8updgzUECNrcWM81IYsNMTyNx03GY4Ikzm
T5eiUZ0FqPK5dQwbTsYvm322+2qw5CDPOzz4TC5gnFnPBoAs9SkxDi/R6wSPBdsnPCOvbq0oDZKJ
SKqIxmX2UtH7iqdjMpFh88ZideQk+GpkN1CbKRXnqCWirtfprz7w/HbiyOOhCTfnP9HxP4qnexDW
1fNWtXdEQ4Ro+eWCLOc0H60Br10TG8rB5M1QEH91vAHo1fWrJzk2hI2RTWePWLXj0ouZoM2lZjWu
l52UqYrPwOsyz/Ujlq1r8aq1kDza9s07MwhZaI87oYJh+KfCM3UIRSW3xW3LdC3bMXBWCWNsJN/5
2TjN8ZkqyC9ruDqx5p/lXAvlI6qyW/oQN5PHvb5Tm8S6Ue/PYlm1UkMojsR9F+F9B0u99d26XFyv
7VphDCgri7lfIBKL9NFdafKLIw29vLyxjPYNg0seD3s9kRqcSJIy+YxjvUqaIXzEGX6vMUAaJjn8
8FhS6mbz9G00mQioaMTx6jWjmRFGYBJSW2DXxCW1iFcW95jLxU41w5DK0ptcLFPvbKEMNqTz0ggn
wfz0i++hg9irQBIEiPDtrYfxBYWYyzi8kQQv81r7Sw8osHjrWlf7oTOlNs6Zp3bb60LcRC3cLOv4
2JR2A+ZW26wPpQUkJx+KZbqSPmfftGEqAYjf8PCQjQ4IUOFb+JqXXrzz0FxW+qzdX+UyEN0SZjVR
/OQCG/u8D11ccVnzyAbXBdPQCciwYDCW19YswYVj/8XZ8yPICDkTypG2Gky1OibuZ2SM7/MAyR+b
8wq5SdUUfFX1enpoqfPi6Y27x4tTyzz2MhjDWEiaortV0FGNYGwgixUwIZoAx2LaKXE1uZvwn8y3
ORwQlJmYlzzT8rQH6aWHOQ4NGiumYOafZy39XdpEb/+0W3qzJPAt6SbPNALLqGMB4+Gvh+hlGFoO
nV0XRx2tPDiywxoM503Ia5U5NvGX+2OpRXTaawk4hRKm0bRV16ZiswpjcxxaVaH7QQU012lNvWgX
zeYEHOn04rZd/pduRuhugvmPh2yySBqic8VdhSYmnFiYpw22Nwrezc/+mrvE/r1bErRuIiaLILmZ
NdU+kIilWulNGBxWqZhIsMbzOWDc58vtt5B2aRczLDbpOD3vccVYade2VOyRlEEZExU0N1N6/4cQ
f12qYfazC2u4wqQyWomBKz9u3FTChyTP61Bam/PZ9mp2qvN7tLE10PeeS1DpXGS4Re/C7s3HiqAC
+qE9x6ndx20nByWrRqgvVBYOKGIZQ9W3E+ZJZ/W+cn3PndU/p0fO5B2msEz4ANrcW7WJ65Ga8Jpm
kM2IvUEWEMcb9Fttaz3+no39jWjMTh95rw7cex1HFIcRbWmQk+VIeDBsS8d+HBWCzSgcpyKOtwoF
OjDYZ7lvhna3DrmS9HtGTAKTAV4WdHK+ufXHURCoXpGPrMtAp2FHWcAVGM8N+RKwv7eT7f3SOdzN
2PVAslUhaXzxOhpWvQeFe0WOvee6TV1Umav2jH1ztORtn+vEqdrOccoj/URdzV9X9zl3R0m0kZ5B
LV6alpkx7cYcrFkXQILZwC/Y10ZrNS/kE+oab1zOltzd/OfxZKIgJoz+bVSSfggJYDODoc0DfIDE
DoFVv476UkfWUr2FqGP+GMPAPXbT4AnXL3DYalFKnSAwmDq2RUM6mddFFv9VfA4L7GI/Czp39l8j
jI9qI7UwF+MEtx/G7e3NHYmxJFf21Q+sLah3UIZLDMiWUxz33Hhv3ZMIFEahUzv4FOlpB3WWtL9E
q9HKtDM4+poiW2JJglepq6Vc151bHx30DzGNjypIyXt69lC152RTmSbF/GQtum4W/LgoXUsEg+fL
Okl+DTxW53toZZW9hOquT8lwzfwHbcIFQ4NPixE0cGb4MtpxiP/nQ/p5i5ypEp9RYdgUns0WRy8K
wQhIMGgfdGG1yXDsskhYNHYf/o+gjfjI3gSuHXH1julbs4QISPOJJK8ThSy/8AvypEu+Am4aeRwW
s70dBaYoJLw5KshCFQyJL31uwhmuuDmipv+/Jc0jAFExGQ4synbOM8xwdVdK6RiDilzvnTbVnqgI
/GBqQih2ptbfxflZhAb8M+JMY5MhRxvEslGkUgKh1LqcBUDDhccqcuMq75e/0STLANOYkZvJOIOJ
pYR7uLBoWGlhkuRGH9gHawHL0Oh3GD3BO+Uty0XUZr6uQZyctFM50gS3VdQw80c3Fnm4MsR7Ltov
3pCviDrpC7Zl+m6Aw9VyHka4mWJ5AQ5nqSgupxDdvjoSPCthrtcXHbMvMgdR8vvqERofNSk8kGZa
qU3eMOPw5S7qZan0u5F46KTW+p/FKk3mnyR6wI8GKIOhOtDzdD5DGUc4YCaeTmgENsigkosnODPF
cBZGTlKtEdrfVs0ZwmoRXQpescj8zHe45BqZMSTnfJWPj6WQ5K3DNTDdVgJw/hB59QsKcu+guUDw
IRyKog96Ma9GWo8zhltYdK+bCg9dcOkxc7ni99r3qLExQJxqiVkA9J6+q07GhH/uiYdIdPo2VEgm
pwLupPEV1VMpW5+ldw8WmME9UzwjJ7P0u0Wx8+VWNur9aFY1mKKN8R3zgfyjR3/vg5NKMD5nIkPL
aQF5YpVSQIj35VS9pYq9P9AkYZNjB3kwPmDdLCg8COqse2SU2yLcVel4nelKDsEl4z2N6pCPRYaJ
MhrsUaefctQ1PoC5ChlQM3K2bi5OeBWJzS6K9uacjAaBLjL4SWGrovW0Tk0CAgrGRMnDVdLUUrxx
ORTPBddtHxVznLNlxIk2E5T/v+JxwdqTExv4ZQvz+yUubrk5SvVarqgpyRJsiYr1g99QzLzSgqq+
NB9ITRLCuRiMtdLtejWMmDTWR4jbf6O0G4echVcj37Y/LwoQkuthQasW97gA5KKq86uYiBJnm2JI
5xUnCdYyxX3uQRxjNmFcXH2MfWMPw8TQ+HkhgnX7hnfSDpkqtk+ikh1O34MujvgbH129O4VcoOrH
+KybWtfs+d74Efxpn8Ox+tUYtqdBUb+fuJMiAw3TWB3ZbkaX782+2JwpbH3RjYkQqu+m3rBApJJK
KCrd3pIHZgqn2dL2c1KmjACztNipBEAWrfIVxKy8qcbKkou6Tbp9qCJDMnWAa9puSz6+VR0gdjRg
7GMJGbh7o5Q5poo7CyZFEuEkA6kug+e+eA79orVtl0vgplM88+mW6ACaFhB6zK0HZL9PDNM6u/ov
EzDnKaCJCdR2TuQ3h66gDA6DAQiO+H8vAJ36rvX9Sy2kCdXcmzmrr2Y3FJwTXx3M3ahQbDboyJuz
zHIQqpEUDkg8EUqUNyAjxzfOq2dYbImiGoxfhPcdIeTiLj4Sl9YBZ+94d2fXHb1yUy6y1tAFxOfc
pwwaPrWPpm+Xl5EHJZ/JT13yt2p22wqJMnAc/nKdJkDTUmPdaWOoQsTLHzN6DU1ElL6TEmQtCdSC
dcblEz3R8ngKJGeOLLMx721kqX879DB7GnMo5bdq3tCBEGTHW3RQWfSzWwl4wkAWKrcF/nQop/zr
7ysisEFOKH6AlzdJbL84g07xcwDUUqWX7FRvi543zeH8NBlVgE5aibihj9RCRKbrDIn3xvlKSjJR
woBYrqfXuje1SN08ojs397Ul6AqmuYR2A6HEyUbqCzV0/Jsin7tAiCMi9HiD6yqKQPdB4sC/gX23
fuR0W1prqSxMkLVKyUzGHAp8LWj6IfQ/8SU7GbV+Z42qm8x3kw4oQ/UaUfCq8a+oCv3jER7or4bk
7+Fms573U/yyX/dODqJwrHqjcWmHjMGveDEiprSEUHih7mGzBP1jWqW7yacUCY0Tw+otdNQ6qpx3
KmAdvePGsbW628HZOGqWRRHWpcyrxB8d/8xzjF7rqYWekjcJkisqgXiWMzfkV4G1BzwPE7jKMifT
KOGk22ZElG9pZS05UVJSaoH26pT2x8hJpbNAzzLK4lJD5aLzZgw1H8W7nCn2/rkIXushZHdYy1XO
CYIDOD0UJ6m5if+htOwhAiakmDURaEZ0in0b2gBlOYPIhnKJ4NaCcpaBZbMmveVQMY+34r1U4c6o
qoRHUlA0PzKY8umRNM6E6FPtSacbTo5sMdkUz3ltIOlyrZ9hzvMUD9EvP6oc7SCCpyqqmeb36YUc
GgCIQBM6ps8ZbFkVRpZEkrP/mojgAnEgnYryRx1KIg4gmdnupBKFIYZU/xZHkoz3GABbl5opti7W
R28hWLSIgqndB9aGleC+roVWg+lo4JSYo0WgU8+rLwElttRbpCWJFq/lN5ew1TtCCusYF1FHl1kt
9l0EAXU0ydp9GH+CM+haj4SIhk/8B906rSPz6sAEqnFPQPRZ0W5HaHwKVsswPflDMjq7ydH9YPki
AUz0m5PwBE9ta8wMIC1PXZtkQWRuZXQasafUjO5eh/hijdkubHaade3HE6T7m+MSSP1TX784CjQ/
r2MtUlUwywV2RZON83cfUwFWzLuXl8k6fHkI3O2ZSKZiFO1QEj6JzyA+birYQJztIxrdG3U1B/lC
cNVUo1PqZHJye0DaGwraca0WurU/spQgIXwmXXZ2Np42cePYSj7PkOGW1lYMQ++WT4/pxJK7ShpM
ZKqZNlbeobuppDqNCudl1VQQPkmDTCSdhgz4fCqcb6BJNPQH7g/3Q+oY0BHWjWH1MwplXg8c7ADQ
uxzaSZS600hTGi5VFDBNbcCEV1PL4ObO/9hTOqeX/EaiZGOIwVfHKSJz/bZrxu5lsq3n8xn/OjQ2
9QimPvJquto+saLVAAUUJq+d0x4DKYXuBcItpb2Q5zB9tZwPRBYubvOcRxrQehUKMd8FASuF6MxW
cKYPfTQeepzqKr/CETDWJ8qvfnvLVUUbAmeSXoWXNO7A4umCePBX7buWTj6fV83jMKdXmfmN8oWH
XaMKmilPr9plka1aqiSHmGvalkcn9ja1ZWN3583iw+hP4vaa0a/NhhuLpK9xPxNjclV3rfDGEULD
8gUAwjL45Lm5r4766QyPLHhB76mkVPtwYSwQNbliJ0o65sa96Ream+5c1Gr5ZqqvD4CxWVzgr7aJ
C0shKjz+w6EcmviYVK+bxy2EJLFgYY3H7XM0BjUguX1BIjVmQCzIsx/xdkj71dQyJuSVE6FeEy+E
u6NDc+8IMy4HcFEdcDZ131/6wp6IIKYWT1CEit0Ycjj6sfbCn2PvGif7R3J89evkb/ywC/zLM92a
ns0jNnx/94eSKfeBo8MB8t5WJLq5fd2PiLXYcjY36IMgOoYsh/4DCx9mpnqWRqhGghBOY9/lvM9f
dQZ3vqxZ51o5Kcn6zROimnPjbL1EC2tYVoI+1w5WM5gewzWrJQ5sy+g0hShGRLSdyCUGk679XiLt
mlntXDKDAGIA33kEtShNq4Pwmsi3qikao9V4uM5p4Zuzt0zd1qd8zgqF06uO/DvDbcF/I/KyF8s+
SzUlJ2T6v5xYoBOaILrbkcyoDj6hWMdj4W5ee7D56fwBSIVFaQyZUYZVF4RS9ZrWT+YMk2XFl0Pe
HUiWmOLA42KMkj2IuadGyao1PCvn3Amjx2INyVeIU0z7QPUyHXXPBuVu+5M8A5WI6sdc8pu9igSr
9CdWul0j0Qa56JgEBjnrbPMO2eaNIZae8pbSwGMRzPj0o6zlpy038Hv1us13gaSOFnVe7zfzZhXv
TVA9bxL34aKlDP8Ct9mfRvMlTrZjhpsA0vlbib9Wh5YTK5G381s3XV+vgO2wbGINRNfu1tdz69S6
PKZOfH6KQ2m2qd1AYO/PlulzukmtMyB4eCKPcuFQpZsX165eq/V6XpebV/E7XQukeHqGNM7ksE4x
QOf76lv1TxGRQSkjxpOKDx1iZgdWkT2WFNf4A0pOwHsd8A3Dag+tu1YxVlYc+hvF0TO/gXnxFsTN
gLbnS2y9kxcqbvF+UQmeQtogou+HwY6Kz7C5MNAy39vpb93fm+4WIRGiikYRMV3MQsHHboWyg/Pe
ZNNlABRBs4UDORdZuLRISciB3QWKN7sepxYAXQm4oNexHPhhB9lKYNqDtgxgE+oA6osw04YlWMHh
SXZFdPbg+H2Z2NGvbkp7uY9tkBJg0KeRVc5b0lA13AYoQGLWHTot7PTs4c6Dq6PXMx6z0XSjAi9I
E0hz/TBnn+WWFABv6fKOERAL3pJ78WIo6FoQ8eoObuBJTpyhXCSMBq1Hy/79NvUGsPFQJJi3H9xg
zKpMT4yGoYkz4IZCv82bjRzlzOSt7a+HH4HgEnzavG7SFbQgWideuCMm/wwVL0KCNpGYNxHMXgPq
o8j0WD4c1gV6aqTaaKwSB/QZ9UdkAUeOSpceEAyh7T6RxeZkG1A2+z8hCgbEOHalDcssh2WXoBhn
crxq03n1Nt3DBP7sRVB+O2C6WhqZlIicuXHnGjVh6cadmV0VgKuwzealJ5jyoH88Ljim3vKC6F+N
U5TPchCcJB/G8aGLKWtQ34sFY+mkxb3KWfPKfzaZezEL+1KpnhSBRl9JMnGJG0QTZXasZ8Z068NG
/1eXLAxyVnVPluy2TDmdZCCqkuvuEJZS7VP+OejSTUuFGhIApGle8yqsETA45g+dhM6g3mO43TOx
IW6BilscvzfFJeRit3oDOr0a+toAz4PR8SIxVJkUw8o6RXOhW0t+ix7DhkRirI/riZUHH025XQuO
zvG1JT1d0nD/+duURiWZxlg7ae4ILUnPcEg+mSB7i/RSylq2iJl20eCyTdN4MfNn6IOgGPDZhZDq
TffnaEgOk28udi0v2R+z5WPkTJQ6YS2+FvIbfbUhQERh7EuEoRxxDvP10gOZlppj5eQiNkH1m7PP
I/JpVJ/J1CIwQMmbPymEWaAnaKbxAuSaT4gHnhHkY9N23yw2dchhIlJuukIMB/+f+kXoX6hPeFrv
rFE/iHJ4Df2TeaTheX1N+L9u+491JSVNfviBpVUY+ICWW97dWpiJS57Cyds3+8jw6G2dg/q1v8Wb
YgP8SXbr9+f22j46aeCSyoWDWSBlP4ieY7pRYxJmSTdk3s0GV53FAd1VroskNgnHulVC6X11F+VT
JnJBOuzsoLBF1sFSjRluXYD0ckbGTmcTFj/4Q1Tc6iByU+enO2JPXtGHXFTU6O/OuMq+CJOdObEO
eDpqp3qnUI/r74phTywDAQFD4m9o9zyVYG62BT/XM7L3DZO1Ph69P2YPqPs3O+ZA/ai/+eypJdrx
fjaXUozvEaPtlu0KbXxbM8F68jQ+YjLCpP5kc9olBJv8Qav0UlOVno/ev4E2a+Cp3/4hLumsr4fC
dNUCZ6/nX8rSd31w4+yYYY/DhObxi98AbTqrEqhY5Pnu07dlS2HHC22yTxvqi7FcL9FRMhMYBUdF
eNL0wPSJvIfxI3v3VpL3Hp8XOn+Y8OLjLweLrUKfRX8CnSk5shj2gMnT2Fl69+tfacPGacJ87j1B
TiVKStuvl2jEfUWfFBy9YQOpIvrQ10hhJ0zEf9oJaQmLa+xbN8odwjHM4/sYD6cuLwop1liWP68D
zYjqDZ09WsypLGedpbMoKZwJxpuu9ygic8o0clOBlK0zUcfIzBfC6qtfmmMXrX3C0IIG/5mpTTtp
UUemY+2G7yOz8wL/b+6RuEx40LuD8lu0qXcCAkjVRyLnzx8sTj8q7loLTUf8cS4yuD7y92xKerhC
/t6ceJKP6dvOPATggsmeGmCbJ+PBC7dp8LnSLG06FmnSkH7FQ/7jep332qSSlLSZ0go5q2KA57uV
USSrbTID+S8OHJ65BiIDSNVopPtqhnvVxGWXrdbbYJ7t4z5i8Fq2c5wmlmsGwFeobGVVIt/+uRgd
W+K+pwMtglNa2lVYVWBbbwUm6TYos5ITDSwbJaA3apfTZn0nv3x4pQ1OBP5KBqenu8TNZx7zP7gN
0XKil7vT4uyn8jaXCVkiUCaxziMX56BgTWIFhej2ry2DgIXpGPVjruZZMoUWS/ifk6FJuElC3Wfl
hNv2bTACVuM/k5Ip+STzSo/OXibrcGWb/pTv1+qusYxy2q8wZGd2MpE9WiP8qUH1CGhN5TY7eZsI
xkwN7RT7TwYClr/hWq60JLLeCghrgITRYD+fuvTzA5wqDxgXjWVDw2rbZKiCZGfIVloUshII1xxY
sTQUFZj4ut3hkC3PSH8Ro5e80SesT9Exz48L/9kyb4q14cLa5WiFiiUXZtvWSpjvpy3kyFDsRynI
DXw1Hli/vtGCg4yG1UIaocd9D5r1AAGwYywwKFKT+ypNdxP7j82VsE0KCnaN72MUk0ytZh9HaT54
UpQSJHy6tnnwXxPJYZ1ous9F+rc6Xl35IWzurVWngYrQPkalNsTEBq/C0b2pvauF+dUt2+eS18TN
xKHetBWhWXkql/dQMVj+NEITROz4P98GLr0hV6XJca5YCnkrrL8vjDpu/q4MtdoNZyWfq4A3K/o5
ymieFLNNEUrssPEAzi74rGGzIdi+I95b+v8NjTOrfXT8t3GQwPgW7x+UANehl9VVoLNpNxiwS66E
uU8/aPL0z8yTjN4xFYYWgZKgaqrCq6C6n4oFzDGO20JPBeH0sgIKckZSAvPB63YvhSlxpgIPicLV
47y9WZh0F1ZvSiI9CY1QE899FH5dSEp/zvXAVTNSxKEhAYDbGd91R+sLeVmOXgtIzO9BkSTM9ofy
TsjhcZEyBESZCy9Nrcd52cwvAZp89LYnxWPAgEbY0FYV0H0LUXF5haSRMzHdp1xwrC9PIXkOD4xo
4CpUMZxdQbveYh81mK2uWlx/5RfeXCVUCCOoNQoH6tQXEzd27CAEmUtieEVSY2JzQlhNOhdqMouN
7KPTT24cTzRvDD+xiXuLBgTAWfPX3KRRGYFmR74W0w91BZBDJRdx+sfwbFWt2zbXr3jnu86ny0Oh
FkYBESnKAHkdtGY8nabCbNgaZDcuxX03jKPNimd7K/8CcM/AyCA8RzjhwfaXqOWbxSYvf0JG98cx
T4/PMYRkuF9dp0oUeoaYnjE88nxszsLznSaPU6Mr82ynK2ny+0n+cndKTzXC3PC2S3enGcSZvhEF
4yELlPNChG3ZGZdCSkm2Iyc8bxe8ug7HwqB9nPnPfC6e7A4WJYjHt45GqY9OZxWObTps0FtxdNfJ
h/RtR70iAUJjiHeJ9h3hiuWwzsaAKinOzAhLqTzpojjJ1Zra7YDqj2HToXYqYeOWlch5fIhKH8QU
SMO1RVgN8a+a/zHts7YsgIRsEKJg/JMcgVMjZkdCUd0/D1pDVDBP7lgOc7me2PRZlsrdw7Q7Onuc
mN3LelApLBIv/Lqj3Xjk73LwV+58zF6EZuCL8DkYZBQKrEeIKwYX8kCGerDjiE0Ad52X2pDsV82m
tVxMLkU5ZKbidC2x5PVjNeVk97qCQ7SFH8TV4gMSsqcjb9Xlu2LEqhh6kSWeZeWLGEw5KefUG2Lc
8VhtydxKJyWGetv5FAa6OX1rw2eqfAj9I7NAXzj7blkcjYP1IVbRxIdX+WI2LFNxA6A6q+Cl8opU
rl1xwoQoKwN5FxD352FwI0/C+wezC0pOT5/aoon13gMGKljXq4QU5Vaze5KluLpHoDrZ7lRbVXSr
p9rKfJYpodl6NbbgmBUGzt54L7/WXufz+rko2Xy1NSDVVifmk+u5gSapcQWH6ywLScD1/bAxEfg2
qnEK6Tp2rIvsPO3bp+u8R9Wz5xZcXL9781Yiuw1DaBAnJ0URDsH7p7ZeIFXnAFbQhVf7Zr+Vnhch
mx8QfQp4H+SrR70Ne8u4oz2uNz0UmXQiw+i7rooXCgOURLm0fiGnzwqAAK1DbgcBABwcvRaVEYPG
gUHhlwq5VX8DYab3d02uhlcN+NEqB9UJaOEOCj7bfSpA5fIt2fyaHHTAjJSWkaLSKn0pgWLav8Yv
lIGzjTgqcV3riv7ubVl6l0PC8W7ubgIjZiRHz1QIKVM1h1L6qg7SR0wROLF8qzyC4YVpwYr8mhzD
ENra6itiWBAAzFhjsNBYuePE0WKGKyQJDcgXWn85Q5WYg1gBgiNv/KExsq47RjL+5ZMJk5BfKV3q
GHZ+e7V//hRd6/4VJInRcrZ7oRCRgd1PFioWCz/tO1vivwskKkGLTtJ6gBrMvorx9URRX9dEcqgQ
Dm0R/syLl9xM44ObCZT+bNEmizz6C/X6TsW0cUErobWPIO0rRkeyg79fZyjyWvfCxIIFSdFJJDp6
n70XhC7vZoa6YFTCB+udx9kFNZxptJoR4LyA7R9ApWEcoMi1YLYwBPNwalKWzeQ71f5NfvlkuKOe
8XG4QwNzJ7LMZA/dm56hJN8GE01054f8i73Jk2mxn7PwnuFe4soLVabstT/lBO3hKZNzlcotROj0
6T2tjOYoL4vwQMEpZk+VpDePOhPCi/RMOt6/5XnVIPIXhruPxt79W+BOwNJExqVeNQgpgKnxh4uC
0LEX9tcECuP07ODbnM/OApZKDhBfaNMvZz57C8dsIN7mTdwAMR/9E1m7jJI6su6Um68mICjqAfiY
8db0MofuNa/ZHFrjnTBqK+zmdM5hh9aHn+zopZcpEbWz0zuZBZyvb/srzSup3BuO1Z4VisSb6BkA
WEwTVTEgfqRyYIPef2Q6/0JvkHZqK3jl7Q1A1m1UyncbH4sC22FBKo/ngiQ/F+VpZVmBCqBGefkw
GShYY8QbwlVvpWaunu8mbtnQicGm3Oo575m4EqbonJkYmB5WiV7fUM6AWO9cG//MuTvwSWCh26GP
knwV/2hvUE924bAIIZku1AiK83HrgtRtm/Z/yRqAJNRoTLiMSOFbwSl4fbocwOafWujmU07r/wRm
/l0jtar9qMInGqN49aYFXCky8bJHoZtLEvh0CblwrOosZln6XEmAn6rpP1wh6C3zq+Kct8R1L+vr
3vdZrBMBlgRhQd7ltC/kTEqU5c0LqZhzRJGsMktUDFAiqM/5aCONjlcxGPKF9OqD+udiTO86oViB
Ulk/l8oZfjPdVmSWTmpQHt9CuLZtGeQp/n+1rf3Eb7SBBi/JuVLSfM6JkprUN9QXy0JXK8oZkR5c
wJh/QJkATdHhqzqO2zUK3/IV0LIJJuyUqS4Cr7NJ4oiw2+GK59H5M+xjNuJiUM8H9Iu8P1I+f+rQ
FR0YGt5b+pi2TGX+KaXaWn2UKMVU+aDKuQvTUsG7YEal5vsrFnyXzQtWzt6ua9DTSHZjcONxb7c/
uiKnlpCNfXFJ5EepsZKRT+QL8lkkw5cX8kOPWVZmnICvk1FRYaUeRfz7cjKC4EoiMO4kvnssP1xF
jMJj6atG1xgNFgjb+HV1qZ8rk7b5P+dEoh307+zyAhutK7P7/sJsbyEJVsVzuVH0wb9hlrOcFwYG
O4ridvUW+Tq1KBOpvC9gaUpcZzrFNRmdHRXxwDH5lpUbzeiMO/3sP5xg1Yu8ahOpoo7IyjLfTKr1
n/QEyGtkS0fSyybTh/iuILpEuYkNd6UWgwCCyekhT6abkszi1NAAEktFOn9QiPOZvP4oU+o9BcWz
Tf6L0+SISI3RXWoJJQIAwZXwsxTXKX47FFfdBZE63NczHGAuVvEz6vw8PJH7PxSImmhVKQp3fI4q
wR/5H3fgXM0Bh57akI7bEPkwiEdsQHBzIdhwN5hWeyD75jsEasNTZsV0ILDANffGGVBsM2UQk8PJ
Ea6onvoA9/rKYu6UGPmQsdxfzQ+9DPy8NASuYUerbHDT7tHNU74WQGUVDtoQLyWw9PVA1VnodGD6
hMG+cWJt3+VWCEf42JHLghMUdVjhLjYOV7ch+X1En0futxBQdnUeXY8lP8E6GiQbB+R8nPJIi0hs
iUkdwZ3NhyFwOGS+ExxHEKku0UbwXcsimSfXn6yAy/Ymr3dHWWb6y/9dCxJPTwEeYcWmB6uUajqA
FNADYn59gMD+XAd1so6y+JMqAcrmfyDjzeK41Q+mQD6eLxRgHzdp57sc8e/r1uduJF2QFVYOZg58
g8l6WwPHN4dYBmxtH/SVewL+j+gGk6X+OKXUMvLMTUOAmIUHSv3ooqmCs8Qj9TCRQGpbm7L7AYqk
MjN1+sDg8iFd5n7xPRAw76+J3+CONanuzLDJk87VFBM4t6VPIgtorxpD5vVtgnW7Ejca0XgjDVhm
JQWxxm1fAhhfQiniGDqOHP7kdNeGha32cuW6CzJ8OS6WwrlvEtTybzCJRx1xT4XHr/vRo/2zg4q/
Kku3ThNi/lzkA92K+HL5ZhUg2+C3Hpuh9zM2HaSoshWOphelpGn2fAPwM4RgYOj/ePKEgnxY2tda
+wfM0AB+UebGFOchIoBDLfB2fTQG6qZG7RTcxss0i3lZXG832LcJrMFfzfqXbIc6YWJjbWi1Cg+S
kEbUemZQRH/kDRyyOtFahPrpsZGTmYQsZ1W7nY8ZxfRpNVMmZpTJP8HCe22Hqzf4tUz1dN2jMnR1
KBlQ67Jbhex3s2iLMLdHtXBZod4XSc/XPU56lx1DBMhsvT2BH+zVz328zfAO+i6RyOJKY5htvcsR
pxc5HVPWKs+ClBd8ThdlvR6wqPtQ4p8FyEFdvjkfyRnWQjw90LT4qUKGL76v0kNy7iIzcjHupFLl
TtUJduUY2koDiDPflkB35BkChV3OofSbwse3CKThke4YFEna5yY+2Ch9dX/pZeJQAQKJ3t5KApHH
wqAqCPS4i1uwmc3YhImoxQjTI/Uvn8ukYsbka+gjNLyaNf/urU0iyl6fI8gYTFnVdG85ycuI7NkK
Ih10upsZF2jSZB5+82Z/8gSWpBkmhs+lT8H+egys23/JiRW6t/B1WK4Tntq9XYhNZ3okAtgy3FGM
GmqPb2q+3tGs63Mgj7DxD7U9H0JF28GGe4CE3X2X8nRqEN84on8h5Ok22I1pUQDOlCk9A8FQh+Ux
V1eQysWhZ7/Yqu5vn4qI1gUtQzi4iWa3ZemPA/DqDlgtIBduc6uk43LvuRWkud9fbsXQ4p6JS//u
6GWKEHdecYIPvKnsyEqhjy/JtNA9ekap0CKmMtBYo/uQZsXnVczYHpYVNRVZarEhF9OgDishbM1S
t0uhKAFzgSHW8pYJipyCm4wsjxx+B5q/PuTKOFWcJLOwrmYtnuh0rmVRKLWCp0zuYPLkAFSgTp5H
4iUayLh0j6T1RBtPsabBQugvnZ+hRL9z+2p4c6CfN0jEYVhyquu47W25MVr1P3ANq84cdrC7I+N6
AxQx0rY+wXFu9sdpE7R3DYdD2gkTvgQv/LmsLikp684i++UBON+wrtjM39ZZwC8ct92jRgo0cGjf
w0m+61gfymbggKo0nnzk/qxThBPB/ig/oVj2dSByuVDOu+0VTtlA6yy7t7LKf1aDQflB8o2SDMP2
SUscx3bAhgtXeopJ+th5E4yzLeoFrV31Wby10qiVGvON3zr2UMTRq9nWQGo03KoDRmsRW4SbRftb
moWcYA6fxHDyMoORw6lqi+Nl66DOATxLmepp8v8L4i3dzrbc06uBOKVM6D+XWDd/v6EkWB2gu1zf
XMAG7IJDM5aMrr+aVWfsJ+HJqnXwmNJXZU7zb3hTY1/f8xUkJUIHK8ZKdIt9fPAFKG6+5a+FWXZC
JcGfR2Jv1wBAWrEwn38y2go7iXDNp33xpRuAXEBex8oC/4AbnjsdslUUj7eS3aIzGriI4iFBw89K
HaiXgi81jh5D39+kvs9GKtwU+ZhnjVXunXq3zCW+d7XSJ24EUdMBDPEyWbTVS2yz4eRUv+e0+zXU
ZTwwJkzLLNR6uXX4omUObwCF/yJf30rF5IL3nx9BwJJbI2rbJO71lLX33C60pM04O5X+shggl/vT
tHMN+gugksIgAOG3siniyvPbk5kZInaz+SekRB1GTwXrmcB/hdU9SwntQorNC6BYfpApslIjLvzZ
+8rIZZ33EdJG0iH3fLOh7u+cUovPofRVb9R4h3ey6KE2wv+7lHIy3NpSTxtEPz4yyoreMu7vGsDQ
1fKD5sQd8k+U+4HWFBuNc30Fqe1a6NWxD36d0h0cmlMKMI/+fDQl2OE5WpPSQ53kPMw3VmO+48db
//ATD8xa7k+ZSakRYB1UbkYQa5P6H3KDy+vpOjpJLrVZMEHL24DmYjBUFGRKkQC9/fYu0qobhwLe
rDboh+QMdpCnt79rGmodS85VoqeV9KRoVbqq0MlHF2ZE5xuKxQHVNzOBBevHJS375y+pthu69MLJ
/JfFbM3zJ7cZUkuEoexOsb9FnwWBGx/9HUTA9HDPcLS+B2yK2pogaM+hpxis5TPhJfdW8hA6d1ku
Cs4qCDngqdiHTkpWFYytLHtWXIWnn1pjbuv/9oHxglk2sn4pS3KV8qP+Cov3YtHiC0qgXENVb9cz
ggPOPjJIaufwJJZJBh5JDfyON3omxP9mN4cKAbUAQjCSJcOjPrtQYelcqmlgDh4S3qM4Z0YrBofD
lLO0uAkiR1WT2JyUuaz3aDDC9p60JsbzVRA0TZ2aqaHk34n/3TsLcpDiVpm/4d26BM7sQLWLNmhY
YmiYCxTtNE9qwBspyHA+oZoAhdV91oWIeY/jHljBCI5CXuGJSvbewHIZ8ElXI4nh+ysWieZy4C8z
0cFt1mMjXaAYWmZmCMJ6acg1s2yOo9zJqPZM1BRVnI3zr1NKjfX66anrSUCqSoFvQvaVxLVetCnv
lrI1YbWYlDrx8CnZumSwXEsfSh9HvMaGHKXgwP6KTXVzemrIJxjv0H3JnKdPmqm/YRz37/QhJbEv
U2nQGDHJoHTIbOcWpJx2RlulodwWjoWy7Ge5J8HE5aPyVoKMG0Bvm2/8jN6crR5DDLqVT6hQ+rUJ
8N724VdoFvjxZKkUdJo1QtXUteab/svcuZ2Q5kmf6OKLywjETMsybKnvRzRm5jvuW/TslLF+PoPm
6U961GgZbrenmWCVWjFKKU3RbA2eohySx7S6Yt4h4BBpPos+1Y/mpgYdBBz20pBb7s8A9X6ovQ+P
7ztuxENXp2GHjdCMV33iCJ2U7yAf9V6c9dO6H5TcOhHap4jPgvK7dCUxT8yECSTyXbCRmFV3sio3
CC9UpC3kBcQnx7+qbSGlNaokvYfGarar9F5/jFgeYo8FUeKfCsZwZIFdMOlAsIJV4A1a5c+HhJk1
fmWkTKfbwuAE4CXkjZ5nJ0M3V4DFgYYPXZMSCdWbQeOz1CfYUdbVxFVh5XvQjSRBM29m7qCtLoGX
ko4oUu5pApsfeWdf4TiDF4sSLkodr3HoYDSo/Dj+Phf/MHio4iDgEtyxYXixK1o/w8iY8NFV4Sw1
iH4yXp01mfqMZgZn+6y1aY0Qf+pRSIxPy58O9Y0ciG7zOACaUPy2n3nDaJ8wsaL066EiIoHgq9v5
1Ls9btyJ+1MI0XkDn7ezZ8Zg2GLJB6dZ8XEKyG/9TDnhn+hWaofK4rXB4gN134X9wWeHumrzYyhq
TXuxlN6vtDlGNZ9xk70y5LmutmEdrxr75KKqvAB77sSEgpmLacQF7CkJ7817FuZHS3wZR32Ra2fG
npsQFuMIfUqt26hGcnR3U05H6JGFsgaZ01VsKs8+HQoYq8p3xmHa1b1nW2Vb1d2+Uoi70UO4hZa2
2phI9N2jLCH9lb9XWAHaPkbkSeMJP1eUPnXkgDDBFZ26JhWfNxTYUaupV/r2dqcJ0r1RY/07101G
3B9zMxOMZm2Hhr/El7LToNqKW8ker0WnBpuL9ND5a8MkhKooU2+hGoHRIMy9EVbwnKl2MfjXe712
AmV+mDerX0gXui2tr4ZqmoXHR3f34vUY9vVKCCQJftRZ36ejYuslcfmt9Wh7nFy0ETTqZ+TxhdD+
cdHeFvisp6uYfu3ZRpCH3UZJZt0+vb8/L5kzFOaRVrlxPd5oftdxCMTLsWwMh983AThHFkFMFLdc
lqBs/XMAgmTt2jD1Zf2o33dBNtysgaCH4I1txXCHgiBOXk+krMPe6/trAlNj/UrBGpyPW4HMJKq9
aszyQdo4ReQRp2Ac8+yANXehT70+eAA1lkO7Ddk8pbRBWS6FQt1kRuleUa8mziwb5M1fQgFsTJIa
e10+1HkgLGgAAqNZ63y6vJLLBXogn6dvHUcLQUykLxnJDY5KH24qgPauWFfFtkQm+7yhHTrETxGl
G8/1HY6usYiIaWJBAvbcKXzh7vHQxhmuO0NMJgG0CGwNykrejlD6++YKOc/8RVLRD1dy4ZtKlKOV
YWT70gNkIonfoACNw6PW/VjQhJxTLDRVSxfirRxeugtZu+/nkD78SIfSECsjxL5tOejqtnVlGA84
EldG7y8Y0zd54oyYtg9QaPRxhchAlTYf6QOIr+CqxvmsxQWIcrfzu3bJ0WslX9vkQMxbEs4Sonni
HG5m3mSUYITygYilhaubGhLxrLFoCBT1HS7jSIphsWrrkseRt+Pn98JVm1lQFrW/QpLLqA6X+ENA
+EQHSuK+Yzq0eqm55hxxDBZChJd293zPvr1YBfkH6g67N0OjwbDJXBu70fgwlYh1FsnhzxZwioRB
7k4IsJ7+YijvxLvmQBuPODC2uwZVtmoXg6Wyg3dyKWf0DAn8TLlAxCOk7bcl8sHX/4dSWoCkpNJC
afiIQbrA7NJwldA6yAH+VX3fsO1ShHbwwrT76Aip8m5H9P0ars8BDlVXjWaqLe83bSR9Es3cM0jA
zNCmpqoEgVsKRxzg6Hm1E8Q6yDJZ8yBCJ9V7PkxKtXYsqDsizAbyoagEB4+ynQtSrzwOI8nu1KAK
S/60nhnNg+YJoYsU4L3TrjoeBrzNEaI81U4SsNpZBQcyU5EkV+5BnqR0PcieQUEmBucWIQxwY35l
c1o21B+wRjnxkhA49MZVnlaCYklj1LLsm1Y1nWhukD/BFU8PkaOReQYafGKdZ/wTwHCKd/gCFQkB
PWDS/GwzE043t/+Jwienjk3+EfF9edi4r1LNid6cdfAz1PRcGrM7lLmxWBvDUMhedMZBY3R7c2JS
qNcUTm0INQhkSEQSsxk0M9GempP38I2mJcrrX2QhYmGjtdISJvowrAeVefszyXY5f5uBoLPJ6aA9
Nsze01AP7XuIiQg4X2sXWj9CYLDGzSoQq+nZrnEAFc/okmzkxQCnDksBvD6zLy38ctL3LFb0k1C4
RigO+Vrj3s3xOmoOTVEAFHXxyhpbhHyCh1BeDkSNAJWwaghECuMJt/PKDnfG3A5dUgSd0lRaYkKo
vhVzL1RoxZd2Srg3IeKitXEHgK5hz6xhozT1SyDDOuaEKLBRNqLB1XrV5SDKeQyZRnDRQIVj77s+
vhytr3s26ZNqSycLChmG15OLBDMmXqs9UsZCAOApClXJFP9eAof4hY1bUdvo4UMyWFDEHKLvwJ0u
wcSU+7oMeHoCmGMhvTmW+a82BW4MvwBG5t92gTbFU1gOrl8g+LknxQvNe/+SJshvpdxvaGjqoVny
1SKsv8uxW32U6UBRqn2qiLrRsSP+2F95QrvhKGrEVtGYur96XEZ0utbkrmnG9/Mc3Bpx5lOFB1za
RZ7F4dgp+9ur1Zaf65/tpNsFRRndQ9MALObY+tdugmAwHj2mqHF+ee5aR3HptO0l6gmqMgIwPh1P
SNT/4RSpudN9D0qGcJV2p/7YrBfTHTNc9pb7DQ4mofxW/gRtEz6O23x0KbTRq9st8GXMiwUs4N4a
PcQFVuuNaJqabuLum2ndZdeNAYIibW9P6mFfRV8AP7RYmxRVE77I5Zk0MDqQLCRWNBXkuHk52eHg
33HNXYNhL+/Uw1jWZKB6T1VTMMhcL6RrzSxTieEvK3oqUTrRQJUt0h5Bve/gQSKN9HEYsc0XrEau
kLIS5a2IAS9lZDolzNpu9B46YL5Smr9qaENjpDC8Gu+uibDkZOO88nZJbW7PqfnFI1JoKgPDmCrL
iVP6QoEP8Ilg+r/XTVaRwjycnihpDzH5yX3WwfYGXVMgyTMJmZ05BmS2eCxsBeqW6U2m5desH/Eh
O2I0OxeqJMnwdctCG5b41Zm4eAQy43Fm9QSMTyrc/A+bWNQvL/uNLTb4nBy9IJXDkJqGPcj2UNxe
sDzPXWjI+ZEoZGPVKc7mmztsHPeTjxZeWg8ns9nZ4G8Y/I13IYrBQ/uIEqOrDH8kgy7k5RylCL3N
TbOslpqxaziFfSvJbqq5xC6Jgfldh1L4mJmL25AygV63A5vQpZdZfpN7jTSN0EJJUXiEoFzop1Zh
jWFwwmPEGJIu/NCqKGaXiaHsZBprlqOJqacdnx+nj5oNMSqbD6xl6NH0keRY+ZJBqcnf4gK8tBNJ
eeCW0aUmBTmWLHFX3CP6arPgNi7h35yrzskwEoaRKFEEjDX096+9zmMOT61bn11is8aQUeurJ8+n
J91j6s3jmLBG19APiuj4cV5h2qTXmb21cyx8Ve8x2KkCsFYK/naYS6yjh5nsTq1mgWa6Ioz7Tmuc
p43CuVYot2F+73k7sFWnVOL2AGZ4Qk6MAwQhcjIKO5unrOcp+CXTEF+NqGwtwnFfUb9ZlldDBV8Q
4FfNRs7bdoibHEEzE5v3Ia3NTHwOVyE6ddaUe1B211cISMhPxWfkJlouIpB6o71sB60s0d8PNJCV
ZS0bDQ9JezrSvhyvdjIyB8CqPABXrL7GoA1NyxC4GMWUSq9ZkRITALFQ3vVYud21qPbEZOVtOf+E
M4Df5o0UL9Is3SFutT1a0Nfy+Cc3dGVl3ORBVPWD39dS7u/HHYCxRrbpzZmvD59M/KoNEmFZf52X
sHFO/0+ij1HgVqE4ATdst+TccHotb0OPNiUeqhfc04a+mRYNVFY/C49AJm1EQd7mPLDF79XtPrkK
KuOGXqYHyO/1kCNTwWvzUaJ0+MRKfnny0QfFUIzFZtAhWhYOHFSNdi00/DQbgQUKkGUbs3M7ejxQ
UM+bkTOx0EPt87XeVi1dBCXYvjRZxV/kx4iZtjEpAwRGh8uluugRHaWqWRNJ0r9STP1bvG9cnka1
TU+36YQsHmVhInjR30cuEfbbvwsWxYOJL0SMPk7Pj4SbMk6s8E0SVb3MdViRFCc4T70yyLY5v7rY
ydgpBILSDUyFVM25KsMmsZz4s3pp+FBS2EXaczw/ONKBQsVmZiQKTI+I8IPLRduevnD8uVvj+F2t
OXgW1oNt6lTgSThiSSKAPJfMA/WsmR7fudW0IxcEiQKDTl5oapiDllPglyA481Y53ZjZMmzzbl3q
zXsy9UzEgby7F7B8BDI8IDpvGzLv+mCo6y+jybe8lVUQqc+uS6vQqRZkEJrzSXRRzf/y2nXVHoRk
+iz0rt9GdD5S4uLdzsTTr4LO8/BcA+SmrJB+F6VuPdrlMAYbTrf91eD5DdAaqDurB2fVK2/2qpAK
wmlwZMXSRVRHq+r2IgPGIxj87xwi/e4TcwuM31c0+XwZjekTbnY3BNdquZYMqtpVrn6GKEKDQTq3
L6vNxgcqK8+DoRNIiczLSQdqQ4E/ckO1VmT0NIzHBjCFuIt0s56GWqd7otOK3vF+Or6DTZLeLCzq
5A0e5VfXUe5qarejMxp66ScbzGL++b6ZfzFlTnQr0aB1OiTAJ831rKAVr1Ft9Xy7uC8cYM+g8wIM
/VPXC0fkJM9KOH80kxn2PyRi+OSazmNu4w+WLZADmgZIa6LmuSmaK3UK4NysgZTjMEWWtoQ97hLf
A+t4xDZuGpWS+2Sg1bWJ/bNpqrgdkpfQ7sPyXY2L9yWgUZ1U2eC6OobSLT3xGfn14K+m+S9GhTVE
eEgrBA1uTO4lzlNH0P308m1xYPgQv/Fbv8W/K6g6Ar0cLuqHtAf4vPNRJXQ4+IXmFSQszGem2YjU
u4WrPiXyPOFPRFPaq4JVFin9yBhVaHzjn/TbhfoAK2tQnaNe02Dfcfv6Xdf+LmDkHWfoBg2Xhfg6
jB9lCsliUzO32M0HVeFmY94TLinsL1IOPofj7WencsDCxpc8t7DlnVUfLps0q88YcDJzeO2o9vvv
kAnXOvMUKWfCpmxHNetbdByKNFSCn2Xt6LcarJceKfiYDtfVZBeU6MHx4hqJtE7cmwbAnRmJMhgm
aQZlZPURKRrgLNIJ0aewm3JYpbLu3RQFlxOSJlyzxVi7nbVbw8wzkXPvo/fkX4hXEVIbI/DfkhZa
FRk4MoqFcW+pvPFwJdqP1/pXdW2yBRMiht9LQrG8FsB3QV9ZhiqHOIKzpczM1/FFk+pFbD/WmcCh
aG/0v4TOgLmaIHPAgUPL9pSyiUx6hW6Kc68wFnJqAclpjRnH9FSF/628cGwn8XYM/QBDNL9AxHXE
eB0Og70gnqEetAfzVlB73bjQmw8Tld6OZl3Jd8fiFk701dQooE0fDsOa7F8L5uxNlL2BIosTPt1+
cLjdDXRzxfvF2lhp4tvtrt1Dw9koBtB9F+4Da6da9tA/RFYgffldC1Qx0DZjr0Re5NJGotspqlCj
f5yxGWzedEBWpMSluaBx+/RsXRHqjQi3Yxvk6yT+YwgSTzoFCCFzmHcXAUWTs2RCbYLRwdfn0F7m
sLNt9oypgmXfFr1QL+wThmisvJZg/nMvs/6y0fiC+ew/md9cEsJwQzagie+xMJBKKgd0GSqbzRXx
b2joOOkb+SJIigMLzzOVonoYa4MjfRYAlvKDnKA4IVpjW23x9I87JMV+pD/glrzdcIsJxA4Hdqgr
yy3LfSifP1zXIbM1WQ7x6GhgOX2MiF0tNJtlPwlfkJAuA3/lB50aE8r57Xx7tsNWU5Q6uK1sPGto
XkFTBZdGkTGnIal0L0HNC8pNwd9TYBVZl/WKxU6HysBD99jkqhTPNTVLPXPr73ptLPcAr3hk1ry+
52kQzT/hx8ehTmLi9+cd4zflkitD5zwpPOPn2Xyc4s9tpu4OR/efRTfqiODcjxhYDtbwUNKNvGJ4
j3jjLr2g4G6Og8QK0BW4eB+3QZsKPKlLML4wx4S4/okmFBZYAOZJ94UOEh6aKRGlusZWRXn156wp
PscsRHI2whA1rhlrcAKWMeQJEmDqpHUjqS2FkPGWc6rRHO6mX0C1zTiZb32nBZXvzcdMQmQ4VgZg
+VZ6xA59K+Ft7dPinRakFDVVuvtbaFphpfmC9ok/FxSyLJKeh16IarIGNag69h2L2AeJ8wYbBbJQ
RmPdP39QpbIJm2Pn5NmW2ZjfipQfs5hsN1qLPTbn95JWaclHDNPheiyRv7CKmnBEQYwz9Gq18qtJ
AWqg74JD+Cc814spvrcrFHA8HnjNcTzRHQesEGUMguX3Uv8SEHlHGcKuX6ZdTb8uK3ILW2Db9/y8
uW+dBu5pdVfuZ+rfuNuFI/fWsiPZTJZbY21fVdBgFbZyks4zdaCNHPNjUpcjwyw9kNl7j+0i+qmk
cWpRJexZe7SL4y9j3R7LhOuHIWOj3IQszhYxqRTi0h1bQq48Hu0Wq0LGl/r6t7DDxqLzbs4QRkeL
y3gxqbB2cG0PuWZBLrje7fFS77oIEfMcfTbHoGxBkBTQgZaTf/tLWJjK4tU3wFW5z+jEThkKrVhk
ZPBQQ9pLDl1bZm7VUbn+0HN/ClmIopwpZX6mfthF3+/bo4mSMM85IXtYR6jSiazm2nL47L0A2IIj
0mRU9W8AREujqv5t9HoyDgsmJpfQyhsGZcYshuxX2Kt2NYdjmrH+EFVU9DMjGUpSDMv30aWMrKx2
NQozAdLxOxG1OcN+jg2AI3gRnRvp4kXgpvOfCz1ECjh4Pc8YnabNyViGtx1xD4jrsbzj3OHO9Kqo
DXAFR0HmNv+RDZqgzfWWRGf8cuKhf4/zF4E56sEcSrslx3WJUrYwLFeSgCeOH/Z5EjupFAT5FF6h
3GbX37iiubH6HYBZOAqdAfsykVVFDKrCNvIL2UbAkOP6Ge50y+grUHInNAi69CwEkF20N0jwbisW
+En+Jq477TTfmFQywCGzTdBp6iN4yFssM00hKHH431Eewl8rStCjAEbqeHJYWT8Y6Mk6GSfMH8lm
8DVcCDoxhgfV70DrjOX5nmOuVNupzAyqolzW4416no6kv3oiimmACfxXzFEl/zlr2NHWNqO+Bfh3
1N92t7Ii6dRua/xA+ugZQTICWNJP8iM0oEy6ymdUgVa7PWE1BrG2E6rCEW/CvdM3yyAqch2ISOSY
addaO6N7I38eCmopwAfSLcsDB8YW3SHDS7E6MaJvskNnQop5wFm1dUOyzgs4bp3K0hXiIBGMn87V
MLnnmAIaDj9uXNrRf7db+VdfC2UqSxjUQp+KdK3IBwoKPslv2AwdMtlAghAagqbOtzvVsyMaFvsK
4jYirK5/WeXxnw4LayRawrcwCtwWO/lyWrSTqFdYgNa/Y9b0VLZP+ZfUQh6OsEw5mHztR+nyujUG
bOU0Dp3D0szolQbw+KGQhWEmjuJr/hW62cmtk/oMdb3TPrqCsMcHKp0wGUL3rUXcJOEtH/cbkbzy
Gu42r4tG6F4b8U9/0g62rcWKJykPv9ABq1RiNbjv3nTbHhp8uYmPyH7r6TeRtMRSDcLvbNHm+UyJ
CbYhtRn9plSdtu34JUrsnVbLWAePzFTzQstGU95Uif8h16v7Bs1YZPM6cWToeqt42bzD3EJuRg52
UPsTTFXe7UY1EcfltSdHZMc2hqZ7Gn85ScddFELpUgZEhNspFylrbe0ZfwsAaOt08gCpm/u3aDyw
xuX7Vs4CX5Ej6NgczM2sjkUfNAjbsFC95O7Y1DyajJGMy2uOvohvzjz6NjoDXvCMibcVVllpLoyO
GhaCNTTbM6FDEo1mKFEcW3x02TG+0Avq9z2V4jJZ8ijjKjw1QpQb5MpmFaZI6MNysjkul12Vqa73
D6ZoO+9HuIuL7tqp7lF0dkcbSjwaCzdSOAcJCrCy0q5NI9IFgIzpswaHKJShyNrTgIYRkY8vlvKO
PpaMzeGWZ2kp7csDz5NZVYROds45FqwSIf1nNhgTeCW1XekR5VjKxLQGBCFO8W1RlvkmPCXq3OH8
UAcy3OdwrTc1x8P9oBFQ0seG9jKmwdClMpgND9sTaTyCQxZ+SGzJeDuxEmordM0Zb9TxLf7QVu2S
Uw+HGlweXq3iQpFUd8PkwR0BBFZRtpa1OTuYw5qQgH6eADCZJmoTMkM9a2f4NYveHMgAfvrmT3cN
8QXyLnNTZkl05dIOSylA0vo58cbPiqptn2z5MmsBSZcsXXO2Pw6j+qa+kcD8yMvqOxBJV0hmKu9e
Rxyx244ZmJDKXRk0Nk+4Vkb1CL30Ia9iqQZ41+uS+pysAgJDfjX/tBJNJi4aj5Aaj3KEalTxhx31
Ah2NbNJKvvPi3BFquMkaBDnxY8/EiWomSlATP2NKlwAu0t1ANhCJw4URm/bUXMbvuxFrKLp1fVng
hCGpylo6wV3g9Zr6Oacrn/O9NCjUYPSU7CSKmWQ4+fYdM33fLbVC0aYABbg17ISvtOP/7l1NPGKK
esgE02GQW2jLHoPOOXf3ggPds4d3AmZdk9GofDHmPfwL+Mda3c0s4HboHvR6Z1nzPkDaLhFJJmy5
W/uNyFkiQjv3jzhTlvh4Sq1qKY06RXE1r9v4fxxJPHohPpn2RQQfHhTTkeNkippgCTcDupJIioXI
nx2SIDPXq+zNx7nRJ5We5XAHVebBXTaHIy4GyeCztqmk21qHQV0llD4rxulhwx1AKydtJElZOaRj
Ao0O3bB9o6RAzKbrv+ijlyzSgFCS4ujwba0K80eMnvEZPPw3U0vKQ1WUD7HfekEpffSkku4WzIJ+
KbUJYtkrYokqRtFYcHInR40YxiJEBLEO5j+Uk1oNv8nmn8WmvKDbqDreEu/ud9Ti9GGQXs9dEKZI
fwIepla4sUhqsf89D+gCEuL13xMjxPBZAz3HNGigVx81E0Bj/v/Roc3eYAL3LbrnkCi+5lzbv8UJ
J6RW9LeKSNRBl6JHlTfC+ifuaTdIt5p6HYSmXifvNpqot0D5g+SQs/iLGPFWecMUaowFKALujDu3
yemX1u4atNI9zNR8BlTrxcmwiz6DmLH45Ad50UQsDM0VxK07kCXZVybrjSko9L6TqBYhAymlV2Ry
tIng2FT9Gdd2mEYGcBa2LLUPR05gbdgE9DH7M75qBQnLYeD6zbXpPiMF1uZlrpAWDJWkBdkjrD7e
rjNFjqw7rnIpEjJ+Q7wNlTrabdkTZpO4zPlnBBQUTssy00KxtjMh36t8p/OW4KyvsBtfUnsJLotV
V74QUsdIG2la7tBXBnoDlAJFxY8TZIufVpRwwmd5K+pKvIQMMKCZQ3idnHI00Se1ruz8HlxstRUK
a2PMkwIUlvPqBW6RNKpUToinwg8qbe5fFu/AjDrrk9IWepkaus2CtlWB0W8L0G7FPTwjKuZT3pzK
lyd2Ir87nwhNEh4MaIZNZBGM6QNRh3MUeZvQo05v9URVAIi914LrkJoACprdn9kF5ZVHvG6IIvby
oH7RZhvsMuVGC5M/6s+A1GaoUOocapkTU6JbPxGK71nf1dZMwRvZXkAWPsJRMHom6701nZhdh56t
KnRdy76Dmf5rvzQn3piL7YTTVJIm4FlRSVgPAo5kyvDAe4qlwJh0AomykogKiWRcyDwUmJIoIW/I
mu1LoOQCp31jUPgqFaNouiGLWkrIq3DhCnmuXoRhvgoiSqtUIa14mUsKCwqYTr517EV3HpCzFcw1
v288zz6X3+u+UpAPQgg0TVGuxOxWrr6nemG7+ftchYVVqKQsDwSRS7Unsv7n7gsSu9uF1KLMAmMe
rVFXE/GboA4uFIO+MCeDnM1eVIcX6+3RFaNXVcfa7UFUpjGXSn3LpvC6SEmo68vI6klBVz3ba77S
arA9bk8eKTmnpknK4bPI/ia3JHKFSEWMCXX+5/L2LpCIvmLkawzwLveYP1iBNieAPISnT5ZQhxHe
rg0sg8SwS4JelckRQ8Epo6GFh0mD6N3EMnIi/IIO9i7oYsuGd8zo4XCMllBTMyFWnWSGKRMar4qj
yQxPz5gJp0gaTkjEsv0vJp+vCyhwyJHwd0h2x8u8lBIEYc3PAbOqkDXA8L+MbTwbkgPI38od4Dw3
zutkolROSMSppHmACnKvYM6sSlTCO82nwCXwlh4dH8Nud3dMVjNmQwcUhV8hEcCDm/XGyvd5DOum
e9pQ0+I/ct5y/XXxhJCQd4mOJ2oSk2s1DxhuYvBeOcj9nTnPgLGFJVlxPvePqM3bV3Y39hO1stQS
icEv47cO6F8X1WsUsS4YknKVP8GRNeoh1fS0KQT3a/GETjFFSnEuBTk7B0WcU1Cpz68MMDhH9ENT
vMgJI+kEIv3XRGda08PdlovuwRLBysINdiEiEmtG7o+nWzIr4ycBd77EAluAjRjyBTF9LKPCY429
mwNG3w0HCHlVWAqy/bGRByCUdzWnaquaQ5/Gkgoq4Ssnj8FjHVXOD5aP3yNRetquiGxXNttZp6Tt
11o1pWXJa9S1dMcfOJO2Pdp1QHFJ0w7PYymCr6mR0dpXVi8n1ZsihE7+wb/ZZNBRA9gbxDtQ/m5V
ojd99ZilYiVN9IQV0oFwgPvdhF4mD0FN86j2lSbazvp+Q5slVYIMlcl1TgAABPvJcpK0v9nCJ+71
tZzPfEb3cWQBaPLVWlWw5eQNstKyY2gb18MoALNbZ6g4DbUDb/fi79PuE4sGzlMGFYH7TIE2aRlf
MqhNN+j28S4WtkO4TBOhkHZA4C9xB1gTU12jSsIugbGPM173mWm8/SLvOBA0xxww6ns43qz23DJX
ZufFfNPez8bvK+QHi3WUguFTEpcP0Ssv7dwJUht0dlB/Zeo5DVsYRiDofkn+KBjX7CMMuGRZ88fi
D5hCqnxHYDebe0vnFslM9GqJ/61qfvy+vHXqfKzhacgmcrL5oDhg2AhTK+Kp5uffmJxLWpqjP/S3
usqRCc0f/Zne9df2jkOlWlXsYbKNoNF3rJLRnlXGVL8EramnFN4l3jNHgITu4x8aPOma/qboqIoi
zXzdXOXEmkuIe+Ms7auxzmXg7hfOotLnY9nue3TEOGVra2hSBRe9k4vuGTjk+cnmlaTz58BkvXcZ
Zrg0noIFAvCSiJSuriDX7Rn967kAeLpUbEXqf9ZsGrLsrX6y/qA85pRMDJBcm2CtbdbIB56/dwTW
ONwwc08idIZnrOUxt87qxUl8uGr69sasz/08qOUO1gF3FDae8U/BIH7WEt5i1GFI/8XudMxdNd87
s+D3QwQrJbm424R7cS//ythK/lej4Ki7iJlLtwVQCYCNTs+My4hanJGSsP4DGJfKTmHngRG3J+nG
KxwWV1efOaPmITL7YHc5hlDXhVIW7c2t8CF1BQ0UMZUWysdukrX2KS4Ws3LD8TkQt4oPkq2jNHlg
Bd67uTmg6h3BLf6Ebl2kOSyjve0M9XhqgqRbXMgWBJB0x8IryW+V1PPbebC2e0p6wfIWtKn+2xW5
cKxx78YplirVskpjOAekeuc65stzfYdAFvxT+f1d3bTs5sVbL/+kLYX5l7vseMrXcnpua04V4Adw
GJneliYWpVOx/P4UO2Z23WkaC7azHLaPFHEur8DxUvoQNgddhjBMtEHZZ7yDecWs5VyXhe+Oq17j
UnMcq60mgqb+eVC6JRJr+q/kDdTo832rO0SKcfhDWoZRkvA/GYrmW9FsI19mbu3M9tzfYwBJ/xTV
Ra0J/dcquWTj7A9mA2EblPR86saI0L0VHAeBygXE+sMGzb3yhTuepOd4u1ufJ5S0IO+uUShCHPmY
U3sa/rMJTDTNgaD+k4I8nxXefo50/4+qQUEAYFgkXUla68hKrT3Gi+b9FpV4RgenR2ONuu1jXuVX
HP3VLJ4Up53bV2Hk0/FfLpT8ZQrzWWVspxeL+fxoa2IEEAJBKWkY8JCJWzC4w47iK86VQmchOFNw
IDIwjRnaGMoru2tpBwPxY9OlTtDwBBT/kht98cdO65OB9Tj5PndcTlnc9KWMOEhGYgbVte9HI3RV
B9HZ146BfuLSI3ZO+LrS0XOac9+2+ykMeM4CZ2033BGzycCr/i//hoMlLpWNHpMARI3x2EY1ITZv
EayhBmQpF6hKjDpUIXDu1vITRoFuH58o5lvs+BMIhmUOz0rrlFmgaRP8lffFXS42cLDXn4iYVeAY
67Gfm2FaGCp8xVspPyHlXTl90IqsUxmcU3CzSF/vC/dXuHLv8ZtAJa9WC3qwB5HRrf3eI3Bvk8v8
lrq2x1PxF3sV4o8WwIFWDEccbmFu32k+IBooNgHy94UpbYO/ppfNrj4hOALqo9Y3+uriouQKqdNx
fJSL7ir6SaOby9Q2tkTICHRlq3RAIEXyRUNXSy5vVY+1ODO1ZywgzYeHZqrtbvgIAX+mOV4xL/XE
2ZjYfYIBZA9DYXgbSGGZwaHI9qV+fX4aoxdziKZpyFooc8QYUr+/IsfwhKmOup2cnjO0AgexIKf3
SqBlCxaEQG4whPTE1h25Zo1PoRCS5NTTYqE0o0u9KYxj/+/NHw7ywyjxdSEJUQkxVvJ/HkpNefgT
Ld4Mlc5gk8a3+fRoYHbJrLEkBDOu6YzTF4wRsc5Qm2SFI9e6LjU3bLIExwNzu+oV+9318sy8Apzd
3fzceOUaL+4rGdL4seCBPLJQVRbL/PeGSoMk5iegDqCF9UbXUw0u5ofCElEJoDSqBntWk7vUrdIe
VbF1dnqTmRA9EctfsOeRxqyTm4gVB3EQrmbCZj5w4ZdZ5hUYIqlCD4dCPMAA3WOZgzWZcF18+tgs
h+MlCJmBnx3spfmZ7UsAqUQkAGur5t3E4Hdk3Rm2HkCDOotXI+LCaeEZtjQ5lzhLTdtr2c9yFuSR
VPRBNgCmdpW+UoMZ85fTTAccaLhsXlT1MtoAmO3WTQ7dtDdnDU9cgwOXv6waug5bWXiR7gvpK+CJ
ykDtuScxesmAuGz+QWZIrlJrdIUCRGYDxCKGPyusfsLzxGIcLn15A6A6E+fAlqTcJNGij4maltTS
3v9SZGrQgO1ri/Jrsl1grMBZsi7LRbscPjOVL6i/Cw1fFoRmoPEQGcCkAdYpx7AGwcu0BnGGkF4r
pRF/2vBtExfGpFJwFrlOCIeQTSV+A9ifQVaa0cYmBL4Pcsyf+SVkSFlSbTPLIrYSvAp+NN5pdzdY
LGK9PFcPOJ/NOfqw5ZWW8LAlU2VXMyKIlJe1O7xrUEe77OZCf8iS0YRzx8Eok808IupYknRStF6d
y+qZ+GKLfg1g7JeNUXIwQUrj5LHHFB/c4qmxcllOCPqghFRBS7ypbE422p49pePVc+Xu95ydD1/i
9RMIA5SJ5fm6EyOAmXmrd1wpxQZORF9E+7mHXcTMNrED37gN3ULuAvMwzNkp7gHr7VHJ4mK9jTfh
Xg3mC4YAmjRLtCT3WGnBXl6HwTL8nRfGTQApARkaINfIBtY4JzID5IX/YlWvyHzn9pnecwjZ4wgy
WXycJnVqY9Z6kizfPFl2WMYvp/tm/Ua7koLwCPomCjEowa1c68lVfYv2BnD2ZPjahXfLdeqAy0Hm
vKSyROokTaV3OLDFLXgugZq9qlg5+B/cuTdn85Z+DRQ1uKs6bAnY1jic2h7lxEn88n+jVmcmkgxy
yVJDoCMYfUhw1yvwpK4cltKcPo+N9jS97YVN5nqH/LSfCXZWBmN2Og7ZmI3yq2IPebhRIdNBt/N8
t7erGjXlcxgbvX66XAc88Ac/lcez8WTLyy1UWb1owqzAMwCgfGDpIiQjRKbfOIiDOozIo9TcpPSm
zzzXpYu7u565/zmG10B7htILbl/f7spwLihrfDaX8Jf79K9cFB8ym5r3p94YPmQNjNHe6mC/5kA7
5JYKnqG3+lW5VubEWdWm3cci5q1lUmoivyytzttDf1hlfopnuQqFyviFE7VazROebUiiaz3u1TRs
XAkslj6Oq7hOyi21VJZYNW09U4I3NdJGaCaZ4LssVwUts7dA+aLocQYqaiEdbfdDY9Ft69WhbDFi
lbWzu98HdNfNZ1PP1BilUAJQQftuhozelaPhVi+Krl8QA2xNRw7xhfnVKfYp73fvK7wfi5fmRHzy
7OGqYzoNDF1bKoywE8X8L7Z3MlwLKQjox9KVtmP/i2BeQpxqeXYkPfUme06k2N/Dg6NtWVpcem5t
3StsmUEGk59/rKoaUGwO92rLahbuYRvGw0IPGZ6GkOkURbf+RqQ7qIs1AVj8dudJqw1Ig8/0pmLh
yFniPruLVYaxh6skGJ2DMMgytcAq9px6uZ257mgZ4CLasI3KnPyvsxyEb5VJbFdUapUrJpZHivKS
/pCOyhbukUAFCDPSkOPzJ4GQS5n7DN8G+8PoVpz8aFJwPo1BNZ10+3Jwr1Df9H1i1FFWG9xOBe5g
L0bPhWfvw5v95wkf2ntV2fuRdikfgHKbe/urEjd+NB//HFPTEjIDMTgLWLK5vpuf7NIuur6/c9vt
7UYphGrgNXTHkUrsDg1l+tbyGY3EMxldDzZUlRyuPEDgT+Zh+u8GSAdIwH1PABLuVLZuVP6f7wfJ
+WIhB/30biwxy5ii22gVsrqvr59to0dVmF7OiE2bcC2V0W9PTHnmtrHOBnYWxvVcdVwLjLPZH1jm
QIgKXcxWrWhtpgBT8h7WviWRKw1fDXq3coVrfs4neD4Q4AznUv4goFfminiWzq3U/jmzMsBmVeyR
1TiPkFl6njZC1JcH995aozam/zRVN5acj2TmraMgrpeV3Xg5Be3z0onWzvdqvPDM4l0KFU1nEyif
AGtMNcAT0Vay2F6FJlZXRM5lpPSWud4CBiBUToApj/udcP14KwPPF8dlZq5D/zLLCCsFJvD6FZer
zCfkwScCbx3Jg2/7IBYhT1EIFobaDG/xSr9Uk3R/+jFYOEaPzlGu+JhxlqedGK+OfoGLPH0W+2O3
cdJ06sDelBTegfdRYN54K3jfbiEqhFVotfDdS9H2ZHIN9h1TMb9B7M02bD4rqZileKlRmPU0lmdV
TjIsJqRDI6gEufPu5whI4ajJfHxTz+9jFHXEH0XHyq3frC8zf1EVxtjP+Qq2K0aZaOLgupFKq+KB
KpRvTYQu7HdGZqTkMPquSNlZHcvHeKjHs9BZFN0+wCBHzLg5G2xKxrzVZYU/OicawyzKUzY4Smei
1eu4mHuxgcBvK1kpviKSc4/0j/SU5UmwA2sFzQeaI+Ups3QIXIryg7qdvVSGbypCIJaCcT+bMCkJ
JhpLfpAGpWSW83AHuG3q6LXdRZxIP4MnYsD5V8BkQc5UneW5F3RthSFjKVFYZnA4yZggp5NffDnc
L0jH2q53+DUDhzZd2UU/HPcJ5NENoxVlyBvymamBhcfs74WRt3SYDe1J6XfEMmRy7ENn9mnIWgoB
AmUv0TYsg0S6bm7gBledTCBxAfHpXfBcaQYM6qwONO2bp84D90YEmIWuqKSMTRiWp8noDjKjLOzI
ueHu5mAednbbA90nZcs2YI4aTFFjPjHziTdOIVh7CUXJAwjzUTqpIWt9j8hr1asgvM/dgoWBezeh
QQblq+ACRcQfdWLX3ZwyruMm8K6rwMVYPwrIhRGp4Rl7w+JJbCURBXbfXouyoibxXIWZJK9qWIyD
RpOMomO7IzoedMpkxhGcQHJdFgsLSqdzLsKUsOTEPv1p24qv7klwTidj9TrK0v71uyFiC6WwkvlJ
RgG/aDN9hKeqSLaZfbRHj+1/wlL5xpN1OrzmIXKGAYm/k33SzXXYh44TMZaka+7OhSVSux2qsStx
PGXoSb47Xou+MUuSFMlBcgaclZd4kEmwOpxeWEv2+vG5PcVzIaZbDqisBbc3U8Nq1DNAGGm+1SAY
B6AIeE8ld6VlvMMOH0lc5+ocIEets0kcLKl7lZnF/Y6/7NUx/qOruTi0oHB5dx/yhFGmP5ZSNamE
GTzX7Watnuu97UCQPTot4yasRqlqXHA/LDTURPoj0Z6dskV+48hfknRA33BBiMpoBHxBCMwkOof2
ekGXTK0hKZLXV1adfeYsl/M2PcKRzKUs1bS9JM6qwNb0KI6CeHoaWAUaeVkEJrgvk2UBWjUCbCZ7
9aAEoasMO0L59Zj9EDhrAjfQdHlbsEJia2edFPPjzWfDhRtD/SeqgBbldBPkvSyGZSichYYFtnwD
TSevvbvcwt/Rovt3j3J06KsZtPp/gfX/INBgyKXDDBu2gNilSZSoWdQxOWxfUYOWG0V0Y74m9Po3
wAKr00NHNQRD77M5qmJTObnLiFqJRirJw9KPisTcQWhifstm0iR3LYpMd8Apvy8J0/PXWnXrGfrk
AQPiza4GgZkcM5Jv1qW/5bKMjOkRwyiwHRh28lCvHyQHNhp1stOIc67yaNmmMqO1IGDpT0I94CLB
fu0pO+zquO/lzi5ZhWJr59LIxUQQMnwr6cETFl5PIMHykRpXv9+vl7u9S0CwPDtK0VaFQyWgIiLb
OqSX6Qm3pF1PBqogPOFLiJa7OKHvzJztPPwRNSNF10bML+u0/ufD6GV1eI2QyZFkfocNfhE2KwEY
xONX+IJYKY4rsdzaR7e8+PhRtR1tpMw4Rgkay4JhAPPKTTQT5ckwRlBgS0YAdQ1k8y1mp7N6Hl/q
Mx7BUgeKnDK40ZdVX7+tjNcGUGTbG6hFW0rIna1K2egKkrz3l5yyTFwomakHjK0f+AYpLnNIvt29
GqQsNOfIrXJzfOXp/vSPut3VtQMXag1L1lAFOiw1EnpAKw2sQbL3EPRjOtRxWJirrsfd29JNpF9Z
yK6ddb+apmByg7TFFjN3GttdGThslhwK6hlAE5uFStDbP6+IGn6xcz+EkLYt5J6AM591AVULU18N
e54RQcv89xim3b7E+rzuyuPr3upVXppuSkfJnrYrJR87pu05nRE6epMYauHc5oRFoskoQXhjhS7o
WkL9SyC//liOH6MvXXsCCSBXipy75G+Orbd1CK9B/zmDZm6kFM94Nc02pZfYzJyjEBpJCbAqJ/53
xnxraJqK9yTt06Iat+tGwyBSOdSfrjy4E8lx2xmpFPJY4FLvcgIxe7IF96uSMOxxuRIoWOmPi+I4
dBz91iUPfP8cVW3eiQKp9si09BQBdbhMyByLelyTV2FtLirgrvFxkEW2zu9dVUWVgZIGGxWqX7dN
BneYyA6m2cbHoXRqL20Ga6YWJLxVgC0RUkw4IzxFh9f/KGDRVgqeMsP6cOlGx7gGW1eVVG89iH0p
BZ2v/KTxPKnen1TXuVyqfn1ajwCwUZpiAk5vv8cVkbkBb+j5Kknv89Y7RuV8lkOib254CuhR8ZTT
MBWLSDyw42k67Gj/DI/9VKcVS9glVeMeq/CmorHBeJuqds6V+P6zZGSfbQk2+lJ3flfqN/aGP5vj
1XLADnB/lSUT5nYfD/BOMMinnzI6ZABlCWNe9XgEt0XyzLIlOTHbztVX+TaCwiQgod21ndH66Lvi
pT1kzTrZUE1FM0GTD2xj/wxRuJYckCMHzuq5hJhz2ZS9z16vihSVhTxhiDEzeF3R/vXJHAsS74UO
5+hKz29yl5Ls1YvBydilsvbqh/6D1bil9qd+bMIWY39SjCEExEhl9tf9p+GNMNQIkzkpI7fxT10L
cNCY2Ogzp1nOllBkgbLUT6XsQpJA1O5efj5DAzEpYBIyaCelth5rTwopTk9/XBLod5wg0+XCselu
gZHBNAab0nrWRmgJNc7WYfFf2l+G3PmqDs7DzvUo+hOu7n52J25pTiWGL71fdd1qiNS6A7bH9K5M
ZSgY4Aab6j9AyvW7/er88wVRaGn47nCLPnP3qxFFiNFIm5txqkhsovuJlVxDZZvwk4biIhaQBwTk
/+P3VJS+7kT6itqEqNKdokmI+CdStgEKrNwGDL6fKTP2eO1WZQEp8OwiDBr+2mD9/8Kcw1pXBzM9
5DPu1gZnNZqcONniFPx8pOBX0/7TibeRVX5klOXrbsiFqGPiq6AVGREejfbpHB0t3ikmASQw9H8n
kZYfzf2pewDn6vZlmhgaiKvz+ZFPYkBC/aF9ru3dn1mKNdDtpkYl8VbO2oc0BzYrwEiIbKHxnUhz
bzufGL0q8Nqnd6ggNX7geGg2+wYZa54eEgtOenlX//O2kMsE8wDdpqldkHZmHg+rA/CbHAS3JzCt
e8PBF+MciDa9Gi+GPkui+i/FKJExPjX6Hnb6lXHYU4Mbfc+XS32XUIgCcA7uoRrDSGm/KgICJAZh
bbzDmYPHa7L8/DNy6QS5R6LInKeQB6KuCM9oaQFWrMOpnF1SkZ4FhWTFjsnZ+VhGqe1+//bD9pCI
Kx9mgplO0JtjXsa7JMO41RsPfI2dt0lBhlf2P/a65Drq76tadhoVTyS9FLXeFo42Ez1EqdxnEITg
7sdn1op9eNkZVz1ygXBeBjV50ql/h9Zr4+NYeExCi+SFYLJwiyfcHDlfpl6qIjDgl9BIvETcSHzy
YLZt+DFIqFS8cu7/V9boXCS9HAvCTWamwC0irb67frkXeRy5IC0jtC7nQhmQt/z1WexdrJlx6HeC
0YbBI8uTgtA5dedYugpm/ZI+fobk/I2n+qMTEu181Z5q1cy5GoxqKpDpray5NdxhSNtP5G2QLafb
gJEqmroUojDZ46mJ21NXDLPnTMGvf5uXvmN7WKcIBLxlm/chhTtP7KmGSzu+6PFJ/v7RsMGmHBR/
MawfsSEhRtXf2jnOC7PAZh3BNBVCd3Tl4UyLUrZrykHeWdnnHyLx6HtClbUmz4TS/jy3AKmp7cCN
IsU+xjJ0/ZcaSv8lIz3khE80LFANEU3O4MSYN8Gh3LXoyMRl4xsUF9fk/6DBRAAEuJAHaP+DZgTs
PTMhXv4AtdLXeMYLNNlFlyDZsxjs4C5+tAw8SW30FF9ZEIWnL0XxQz/da6fSiE/DPCw68BHE+j6U
+3jbnHZQAAXPbmssnpYcjZQaAANEGaHvGFX3o08IzXcOw6jXBk3fTA+D43DmmgOk+/kOO86nkLK/
qVEIaYGPuQ9WljdP7A58bTLBVpc/HAWcUhdhYM1pRjqW1d1OSSehtPH4MWZcsnCUVqa8C6LdOghK
d52/jJFmzS3eUh7lX0KaMcVeJc114NmYp+pESY5CYrzkYyX0rGZaux5BcTGKJSYTBWi16MrkWIeA
F46WrXIzhbjTSZVzDaJLY8OPdd5pQIw8KAB1/CD6nLBQiFrt4GDmAdhJsAMYfyociMD0fxacN8aj
oQ5PJwnq6S6knrZQO7Ku/6QEo/s71w7tW0soqWyl6Rk3SY5Zsso2jbOfF9UVM23qXViQcPwXoV38
ZZXxevpFv2rIi0oUEml6LChiZbmcris8qPsXgea7l1j8OU1Hqxmunv84HfXurcZgEIIqdGwxhQN5
eOs085oOp1iIy8NHw76nAm7HyQMuRQQDKsxWH9ctniHIVApseozDhGMC8ujHv26gvdacluBX7ZEu
yckaeJVP05VCuzIsDO8nX6kmobV9I9uLDhzvlnf4wCBXALIownKpi3XxKRUHYqbukGmbbAOnJREI
zEUzLoLWO88DnX+m9rWoWWze3dPV6sVrzKe2EGCtOf4OYdq1csnzJWQL+9+Zi3j1tNUiAX959/pp
Dj0qAHl3nos+96M5EYd2zfkJ/pi2ziksVlLHpZS4Wb+LoK6wGWzq6sl7WN2QEM8Pept36s/jx8Sj
gz/gm/lSr40jQAfx+zfJuQLvdvI6tn9caE8iIxHyv1PyKaeTNKAjePRvobcQ6LNcx4x/pHzB0WUc
iGnzczXf5Z9qs3V1gZ5BM7pEyUmV+A1aJQpGMVC79lmJKtvM9RQNubxuC4VLYVDHXscxxXqkbGgs
JXxV18VrP6b3WDnh9ZyXeRzWQPJtmRwQe5qjWKCsNTPjocqs7xOZR3MZxUECeZf4EIhV1ITbg79F
EAd6/bRtr11jR5FhqdMGUNYeIuOlS2O1gz5vS1cBxN46OKXIgvEhR7O8myP7dRDR7Azg+2AEW1yN
ibWUNBT6gJexM2Y/zCYNblRy+xUV4GZ+S9DdYHr3puByZWr6uA6MLf4eNagJBv2jZ3OFD+eTo74X
EiY/aF3VAUk17je2vTN50wNgGDurVtfnjUubiX8Iq5caxXzeT7HHRSpqeL4cJbTfjxULGSIshoO4
v7IrfB83icNjx5qNjdZOsLUsUbeccvsN4w3sWpcD16bTlUCUAREK3ZUnyacZM3d9+TR78wtTzFQF
jmHMoW2zRn9d8eyjPOXf0sDq6rQZuz87XvwHW4B74qd0iEwIpHxj/LHIAIOiUdAjUjLifm1GG2nR
nl2cHEgk3HlP2067nOyXtE37fRmkJU+uG6hJfajamYl2U/inJCGsyTp8pd9Ef80MSdleJpJbQi7p
IUB/1KrJiSXhGapF4pR732tI72IoHxqQ4grlmEWq2C03Hkt3e19UWujAZavdg5jLdZCGbj6IC9IJ
FsdahswBQeCIDqs2jZJSInFhI5zc0jxjogRzvAS2IQPvT5pw8Sa7ajzv0VoJ/rkYb1oW94LjhKsJ
4pEB2MW11GYrpLYsUV87WjmeGoapP1a9Gxy/yIuc7SapNUz21MUHmkvAF7sVcBIGNv2BP/1/8wYc
eZk5ETtv6pcfci/sAJOlWmXDwc7cBl1zDgwkraUDg7bFwISoL8xbiJCqZ0clPIOdk68iZRfKaRRx
UOt/3H7R48xQBvwo5F+d10WCY1fmtUczb7j5/lm7w8z+8btwUWAoxiJjm/uVyEEKcuejRiShk1Cl
0k18zQ/mVBZK0osY2OL10Y/nS6sA99mUfzMcxx8WJTHMQe2GsZcvwOPPd6mfjVIA0UAUhv5n0E7a
OErg3SQ6BvHgWey5xZHVSgux3NGQ/DEk1JiQ7Fb3VUZJ8pt6dQXA4W0+u09uDNVPSltyCeGkyBRM
r1g2x/VL5vxIupEA/u3eNqNcDcyabDguc4olJBK0Yt19oe60Tvu/pcbmSNCOcSoCjVNaDZrLOZsQ
/gbITFH6biaGFgAh4SyMQ6QsOcIzmciNhkP2K5bDd3vUereweQn/TaBypIPqkX9+ipR9LxjvMq2S
HSMwrZ2uY5VwVCOcfpCy3RKpWZL6HWf6qUS8Hy2lvh8WLTWDmteicHjMmwq16Jqe/L5c3AaAx0Fo
FcwY5ZQhqFu3WYIf7qw7qmUBW8hMoavJ1t2O5pZ2BWMZdOCTsp2Y0L+vRztwA9oNg1G4dNHc0TDA
yjVfWkpQ2JW1cx2QQifZkdu1dO6fSt7EdR7FSzAeVnsnyEwOmS3EDCxr87xow8TVv5EoocYeVN8c
jTp8imQPOsjdcDNniMv66po3rCUKezKuBOQHWihuqf21ohFYZBM94HVi9JDcYLJxn8d+hO2o+oP7
ZFGTwkA74vqZBuguqmelt6ivh9vjq+5kYfHzSYyCldEwZg/EiRIo5eEPYXQFAkPiWRXKgj+Nv48f
Dk/e8DDRdA5R+toGfGk5N6QzyJ71PBFMm/pxx+IP1r4/BuZ04lzq9VDjRL66LzVm395q+vw61FKk
tk0ML0YB3eHMcePMipv2skuDZVyeig2771sfhoJGnqNZxeV3ItUv395RT2/qGlBbq5dY8li/GYDy
23hl+lXjbLmQRhruyMpyXYsfgZFyb+HNrDt2U+Mc4Bl2i4FxGXvtmNUB1AfGtEyt8bfhfxrqTtsE
q3wULrIuqOzS2B7Ubj6D2bnW/DZq5nCiIZJ9bAGn9oKoOiDD+qwMRkqgFxQ3Yf1VudB/CraRp6xx
paKyBsItSfQmWv1bASS5WrF1ZkJ9DupmsQMqinPsL/Wqy3qwWs/yjySpKw19xhb2mVrMkUnX2IsB
r8sg0lIWa6PzIabAyCvE4ZM7VTAIKLahyBUtBCjKeA76CU1awrzysO8Qh63erl4d3Bj3FuVRQS5+
WtyoSf6+FxeVa5+MtxrnP1TpTPNR71kGfvhWBhC8yrxWmoENb3wj3t1hz3t0ueyA7FO8Axw5v57u
8q8cx3TIkb5YSj9TgLWp+Y+dqm/hD6LyuhPZgi2a4klvepn6CeFZ7v6DzPcbRKVfBueKZY4zhlhg
N3a2DBeTCZop9ZRqDEjN0CZeZGZWFh2aZf3sqod22bzUL6nCmh6R8eO+kKx2C+CzV26YEcxZ5Ruc
yJ1IvHyMVAtu1rHYwZJsP8ghawTakPrvG2LhrjPL2ve607Y3LDS3kRjAKxoJqw1D8B6gkZyAWmde
HeUNciuvFBlW1nIR6k+d6nGGrXw4w3rUww5Us0iZEuynAZbzyQ48BdW6c3DfhTkcvYi1US34K8/2
u8X2U0/d3fboFE2dVloNZ9m38M7imEdhCLsyXlG+QioyBxmLeJGAEs8sR9Oz1lE8M6M76ijIZdad
Oyin6MSdVgqvag+Bc4Ln1t1cPexjqH9UdBiZhZoA2NEIFKAR8Ja3PjaZkxbZSPq5v8FnuaTiuT74
4+VLrlz+xYqlalDXcJPAwcBUFn8OXra26cTtEZNJQgTE+TRsyOYu2CAtOVLRPflp12l4JwMDnfy3
EbLZCDn1rF/AJsD8xOQM37yFuilU84ECD8e9ibQCr76pRpiI+UqtFxvFU1mC0O46Vm7QoaRUpJwk
9mYmUeJEap3Gm4rrHagChinvCAhlSPS6EFI3/fv78ohBn2WVfzCeN6u5UYrj7zSapcD17l4kMVND
wvaHIArWo0UEoc7RK8JazuEJrj3+h/0jnmj6zFPif/OfoUCm2yJsvIJpbT1uENDckZSsPaXUZnyY
FGr+p9OHFrC5SxjfS83Jq6kfCPoZ9o/clq3lQC0dsYb5hW0BPHYqePh8M/aPcihH8ngI+fwO4u0H
0/FcZX9dg/xvqfIMjPT/7mZKeh50X26Xwxeh8XAAI6KXzvAURyiqJD9iNYZG0tjyVpEpQr+BrlXw
a+mluMPXOhR3NG6xWYubXoHIPBh95dH9QwsNsBfjk6/4maxzx3/IS8jb5jfFczQ1cJKJ/WIjuTSF
pNCitH2sY3TAPkQkLxBbOQGFJhVdiD5Ys8RwKel5aBFp1b2qwdHfxewmTN8AjOyCUdByoYYE98Mq
9rE5Ak557kVExORy2qwOqLbper6AAe+jkOCVkpD+EHHOkdVnuZ/g/QWk9M1yef9T832ES5c9Ax+H
kV5NXh9kTMhuS6hB85ZBnA7y103/Be1Gw0Vvql6PmhSJkBFcIWGRIrkdNPWRiAgu/CV9lMuSkySf
ml78qtR8z8ILbPFVo/uN2JTvQxFg9siQ1knXnhuwZ9i2dobwlL0dRaoZRJlFvEXV9lRJPqnTZRrb
V8Zgve07rC4HiLWYcxVqFTBeyx/pG5gUY2shsX/ULRazTuQ/tEwGks4xz5Notqls/H+Ze9WuRR14
rey4LvBZlh0p0XWc8MiVMCAmgP65ibYC/ahJd6EAOd46B2tnl5Z/+gQIUrZKf5otG4J/i8W1SMnB
maKRLHh9jZbz6jJLYEbjXA12RlUCg/Fh7wKNmwaxzTFSqRC48BufxCLut4AaIKxdmEPyQgv9vbHs
rj5i1sVGwQjKThOjuTnxvYpxfbZ2/8MpMexkTDsfTSaifiBYWEwhQRoOZVN3gXtQAk338GZCiSaV
kDBkToWVIpcAAmp5/LkCS2ZA9bERlcy4O7biMp50yUoaF/WJvDbu8Ns1p9qCCAh1OymI+15vsiFQ
4w5dn9sXUln5nfqTjNaCp4G6mEUdrnqNEPB7K2PpD2x6Or3/3oB36lLclN0H4z4pqQv36fXke5Jx
KmHPUMMskgOp+pfEX6mEd8vsv4/o/OVFaNfoQ8oHstOz3hqq0a3adOozssLYfe09y10JXOgb60JL
pLLd0Ny/rpOfhmSFQCRR1vi8rCCki6cqaybYKmbuuUqch4VrmgmiBWjqd23FYVaudXA5VhdDPnbg
1U4r+U2N3eAHBMLZoetHt6lBIPV7OQl1jQYIO6d1s2rs0s7j5ek8SJspLRN2EsxELWv+Z4OQb1df
c86aSMzRBS7iDdODZmYMlFyTV7gVy6nAkF3HUak5lYLO5La9+TJyAT0D49nhgvFJlTUtrz1C/FDW
E4pAUXFkNkXrJOHx3cUAM4MRHcTh7uMtH8AESLhrfvzmxbdo2mXYBCRwxST8Wp6TioM38ZHKCHVv
2Z/XR2820khNUJCEPe7PUhC5Uc4xkInteMaZwrfoae+fQekeomuJfI5Cbbz5Rrf7dc6f50gJ5SES
XVp/F5EIwXx3tGBSo+LQZUFdlAnt78/anl0wqp5xfudJwM4PincY+nOKbrnjuQmkp+tD7v6bF9f6
CzE8fGkA8DrsfwJ6nQQoGkf7tEGaDDJ3/MBQGTPx3Da+6LPcrQiRae5Sd1xZmmeArJVupnU2HMFG
xa4gKL+KM2ni8Ywoc8pVruu8tCbsxi2DAMxRQcWERj17mFKr1XxpvD5mBYqvek3TK98I5FslvgPd
LlnhjzF52nEF/bybi0OR77hk9O5cLrycWhS970WvU296PFRJYpRCR7vLXRXRLUKS62yP/dMTu5ir
pvN0KBDj/TW+fn2pjN1/R5TZDUcng5wO81Nrc24h8aXDegXCJh3xAnq+6ga+VJUM0tpGRk/FPzGj
D+HQmifHQeEuMpsh0zEPB3gBjCG7xfaqkvgIZYc8yYEcO95qGFHW0nv+VlE20w1hkDL1nQcQ/7yP
+n+He+gGvNymV4OYFxgOqn/+InEyKP5chjeLiCdiYanBtLeTn7OfvlXsvA0BfHhJ8bBsujfsc+sQ
3mnysqgXmz6OGNaR1KqVFN49XXCEXNXttO0eLhrQyNDV1C+BD1SPvBolfVc4npc7bbAPbmDfQPz6
Hc3UR9axLxR0p8NPms1eRCmv4sb8V5PJXJ5pMCSekOPyLOWRLk3zQ7W/owHnUgRywPxQnRM5kmQR
2Iovy/7N+H4ksW540EMRDKENwvIYnN/18hqIHCcEIfQta1K5aKJQvgSd0/QOsd0IvlOzRpDNqfuk
Q2Cvc4G697LP7bWJ7K9O3SRTqlRzutY/fQqM/DCNCF96y+wnPny2/9r/HeFBe6mXI/9fSTJMngjq
kATrs9DImmvPxen9HrNp5rrM0NXVazIBmyBHT7RIshO+yxQJdAi7DVnDSAUG6GD8krNc5Mg3ftSP
CRKusGC/r0X5AqIFSsAa4Ip7plYnpo9BmkiHAzEoNDfCA79Zz5UknO/+nqaXiWiLMX3D1MZZfWTu
hHsV/yzgnIx9cUQARxgDVMg/merliV/dvQa0XRy/qIRQzYyVMMwBRMtD9HxozAABMpRSthweRpCK
rDFgCoUPSCBdMDmU1cbn6C3JjNkPUd6QbnTLZhcQunQNVIMF5nMq5OH7RPuNYnaCSnfkTdCjhqhq
8Z82Rlk0iyRWiuzq7qY9Biy9J88XtsQe/zcuuqaWCSdBDEuS88zOvISzba8FjtFLO+6DUoryVLBk
qO6+zwHaS/8XH/5XbOf8SnpPGX13lEzkomdvrXuJ5luOuq+5C1g25wYPK9bIhD+SSKs9EnyDWDK8
MNimuL23tKYgrac48nCaIVEFx/pNIcxu4y0lE6vmG8JdRF6xZ8wI+FkWGWRGDqQL/S7Rkf0bmjKO
XLeRTcgpYKpSLLIkYH+TndybP6EubQWNFtcEZtpFwALW/HdkfStjfLoOuf7wriRDUE0DtVl/7F7A
JaAVb5tam6liJGXpUd1aUfnzgkXaMUjTuY+UIJ63lHFTF8edysdZtN4D3EdztikHCm4fgxjvMi0n
C1vcVsvVLFx+pY10axRVFU/WfMV826lLdVM3LIW62rKduntjmdXUNGrsezLofdzAjeluBk3H+uvs
yjj+DbmFp+muCnC/mlkbDgesS+4AwuVfk7G164JQyVgC070nWA8JRQC6B8oN73V6pNrBjqPD0uyI
Af/5nuPGgp3QHQFE7NIQHZMkgpaxNINOPlo1YNuh1RWdh88J2czo87Kf27MlFwXRdYyDB4VArFoq
R0jnyyFEwE4T0Yu8VwyXpUdSk3iSCYEdSg0n8ouAjwI/zhx78t467Q8YCXIUyXXudJL62YAWVb74
Nvq2HxwI3dN0XHPshHbLRdwP9wtcME6hhRGI/KvOlu60ndX1vm0q8Z1kD6au62i1u318dkozU6Bh
/lUalhMDDIQ3Ak5m6qCrP3MBM/XT1r9cLEoLvreUsdqdnqN9qigISApke1FeDc/sDg7/nyAv1HUI
u4S/zM3eBlzcmWNcDBgto42Tvl57lN1RK5p/rwiZwMgcZ1NeHXYko3OUkEAH/cVuYLBiZO0er5bb
x2fnjKjQFXz4HXxF170KApQFs494YWnbj+7ZAWP4mWn0Smx9duMMytMv2Dqs/edTym9JAhI6UYK8
LGcHWKZZ1liU3SdBE4j+3KORUODcXk9/lFyd9WNrm/agfEA87XnTCF+lrjZFrrq2aq0JAf+mHSw+
KkzjYyhLderVt1tFQ8Ia8kgqgFnHsj3/8leAGPfnKCJfx2TEcooPnqV4V0i0H51X//YDdJCy180F
/O2W5qYZmyHr6rIMFjCCSOil+r2I8cxjNGKf/w6ybHmlIx2dQuEfkL5Kn7gGdoLT3hrp1AOzy3hV
g/TUnn+ITIsU4oTx4/URIFR8V8Ri1Lx8MaiYZ8hmCYbBCdto0Zb2d7D+iCerCJ+70dpzqUrOEJ0X
+QuclkAgysWLgZlrMPPM9TZfjQrgz6opoOwe+tiFMlOKKH/wQYaBAyKZ9Uk6wlCtXkahCMG0pyNn
Ul9MP94sZJXCVXYDLZIpY7sIpe8l0l3CAko6oyq2qmFrkXWMZV6A2UEVTrsd6DY8ABLMThNMMvMj
z20gith3PNfo79pdEAt+R9nfb3Cp3n+zNdudTHXGq6Jc+DT/ssQxMLpx2RrOzQ2DwQDYtAVUnL06
V96Uf7tXw3/7+Du1ktF0UjgAROKoHCcM6b1sZHU00TO4CkHzLUQa4GdpZWkpqbAu4XBOugiTCHyG
1AMKY3Lp9A67fgE2vHWh4XltSNX9Uvj1pmRomipvML+Xsn/Jgq+YnQnXebrY26nSrxRZ1kEgiNQg
IVF8PYRx7sQwH0P4UMltZSiocqGgb1rU+KnU/AzRv0P9geZsg9YtI9jsrht4ZTbR1Yy+yYvOSpBj
ZpucHd4ZAkUjTY5ZGftqu7nlym6d49AidKPDQeQU90kJldQtt0K3+tSZFDKDELRHMUzc49fCj52b
wPBZb3oo9vJ2Lp+tQIPzg1w+yVwq5Z3rPcR/MpaMIPdorj6q49bMGThj12FE8JQAympg5NiPJvcT
MifsE3pJW14+hlaBKi/OyXAtIIk0Bnxsa0MKQ9Jv1jkvNiphU1AdkNO5U8VSbsIEt+UfskLm84BT
1sr9wPzfqsg9JDu4A1YQxb7JWkxkmLPqZV67+1pheMwH0H3OK+NUXIpQ67/4ZLTnhOqzYfM3xZqK
XYleduztGumY2wr8BsLvOpOSI4iM+R5Q/dH5oy5nv97DRZSZQe1GY5pYgms2cb5bPzKSxS8ORaNP
gLu9nxZXupB4NFgsJkn7gO17GoVMdpD78RVRxiBsE6FVCqBk/qSFBWBCdi/QJB3l2hRV1lXGjduY
fUFKZsBUWFJnJcI8XcRLLpl05z/9URfwM9wZgHxsff+4Mae8z2VvCotq+9ZL33Wx3XrhwJUHI/tw
2nR5f7rpDJuIOOO/gq2/hMe58Ex6VhRvNu1XEgdQ/N6paKqrqGT5RE058jr+CurjM2/1C6bmm1dg
l+blMFLfCOXSEne5bAVd+IW5fLQjE/o1l0jxtKTYJFzG3PwxnSPTKveSuNCaVjt1SBNvEPA2S0Xo
QZPHmZMT58x/gx1IFg4F33rZpEAlOGucfGB24z5EMSJZkXu4WK3/pPHRRhWlHyRz/DtY1EyLZ7mZ
bWBXHbhVCPvXja4I7hjg6TnUgj+82hkk7Kegvb01Lof0yUiIetKRItZM34+HTYO7SlQgmXMQRnbV
WrR75c5Lp+zFnpomUJUz1WgbOUh41cRKdOq3dMo4WktRoYRzfXfvSScnfQ5HstKewaVYHMJ4NLZ9
RG4xGo6zwZ/kTZu611DCHaR5HFVSUs1U81jk9fromPJUR20Lp86SJlCX0yuuyURpt3tmwV/lIGwJ
LI929QbwrlNuAisoQolhKSxvVs4u2T1I5VB6tjnLrMAIy33U2oy5BSUZZfLNcSc/l3oO63kGZi7+
n8c+EHAuFbdSoN01zxxpgx30gRpHISZbZlhoNghf+RKaxT4lgnBEmZVKQVMUzfPqW2dM2c8K419F
WcyS2y9QNoXRbIrJ7HhBXSQ1lhzoENccIIPHaWovB8ClDqgsDS/jS9HWaB8gn8E9WHpzUm2v6vSr
harAoXsZQNxcg9h3U+4F+WXD0DPiBNN5Oc64JfE68/pOXM5pUzGg3v5OwYvxEY83eMRfdzHcn9yi
kSKeG53wMJ2Wf7+QAmGJ5vtbIzz0BhNlWfeTwI5qLHAmC5p1kIbSLGjEAYWhvh+zc4zAPnnpuUZT
jvhk0wBgB5UocbHG04JXgP05pu6rM2Pp/F5915vIB9IuJGF+LyMjoqMDeoFKJEu2o74O4EBbj6fg
IEEvHII16sjcnk7kg7esg/rgAFhHx/jtxin8xwnkflKIXqOia2FohwJpbYYf0CVuCOPs+2JmXmHI
BCzRkqe0jLWw0dUN+mCCfQ6dFAPNBbYopdJ/dsEioXRlhstPk45K/d0z4OzQnfTuX97EW3PVifrB
e/o9gP4chVpNkCa9umUHGm2a6i8lIHdSBXeq1lY2kwD05NIcc/i0U3e92naB8mNuFWEThmsA/Hpj
W2xd8BOKhliJ/bgveovvSaFf3NzbLh83BVNSQndeJjvIIA937lviArqgno5OCOuJEmLTOW+qTYxO
7Us0Oq02xyWhAIfod1vcclrPp8ziKWfTbhBxGsHgo9ekG+TcEwsT1XHsSNF7x2Tlrb4HTH5SJ7CE
h8B4Z80LyGATZD4CxRiGyPTXaRH8kdkvUWWT9FPEHR5br7tYt6npe9mZGOuBpWtS+VdQrahuU1nw
0ONR5SUGAYmvffkoVlcaBdk1qR90tzzMSGHOShOM1HGwNl+UENxn5sx2ygQPnrW7cHPhVGJjCqVi
uoEeTpUFLJlTsRMeF7WDmIOeiKx2HSgIEunv6g3OoqLFBemsmuhH/HrLP3kDcrNySDrv/MsEfeFr
/rx5w7tGsqDcrtislBlluCN2/YgCewv+i+7L7X0RBXbqdB55Nqm25a4TThCz6WJzv1MTGiN7BUTf
tK1JVYiXa3Nvl3xkBurLxtrfBjqDd1TdX2/KXKv1TK5c0GdOInRgY7N7fw457lwTd/RWd0fpgD5v
6QiCMtiNfzgTnvLcBGjqmQNrPw4q4JyeHH3QZuiskihcTDB2JcY+Pe8ZFC7DIZq7eDhY1rK9pzXq
9/emJ6BDoIsrWpTJxJZ5gQdqmEYLz6s0P3jPcDr5MKbvzpj5y1pHTVpjK2AFOVpk7U48kmmW+ssz
Ksxbh6lISY8E587rxkGzu8E/WTBbIp4gpEeaarYgUeevqIAw3Vr46lSb12r97oiw+L90sfz0TsF+
01CDYQsYCS95o/UG+70KXEjmHPtesgQWKgIGR22HyxqoH77DDiZx8TiprgDen1Cx7MS9KOJW7q2G
DMq+Riaxk1UOJ+PJnXWoGkbiAzOz+lFktP3EuYyDpkiU4cm0PuOBO1lkeLIBoJ/E0Dd4r8pHIx5J
EnceI8qoEmPuLqMmi6eKhmqzE8nlxKWVQxEPcyKN7o0O8HSSb295Fadee9QrKf6tpbRH4SMauD4Z
Abt+8uFeifNMI6ifhPuUTNn1WZkYVi9gOAw8IuEmFbl9S+Myqnk0uEehQ5Q+VJaHX10SZTO4G3ZY
uZcFzvZITygb3KpQ+MDMTJsw+671o19HnhA/MNBXnqcNRiRVp0utMV4I/nPFKYhaCsw/KqCPFXll
5yJJCivRcmJYERQHegObOdVdPJRuVm/EoysbrmtIpXsXK7L7Uq0L49aktb2N8jcsG6RjE9WI1r1b
yKdXef4vqVrNMWplxUPxFpcfABmOc2eUGpiqhysDe2rpLL/7YWh2X4qW0C9oqcizZ8dACJISpeH6
I0hxqlRC18y3Q1LOdvtKYAr3FaAnE8QLJN+/chBOAzl0UjM2Q7hJEP/pNj9dMBiPbA72k8MV/hdI
z9yRcN6uJv7JRgvOf++gp5PNwaADPhKWzqW1owxD2XttJa93v5IeF239KlWiGH72uWK1ljwRmlbX
KZ3xMFm9jU/qLWqLJ5JlFKAVJEQmue/GpamigHcxRtAGR5oh84aVFejYlW0ofsdtrerOkVHmDVI1
imZmbUifO7JDbWPhgMAd3Zzne6o9VV2F7ZmU0cJKBakKjZMqV8KTzzFckcztCKpRHm9hVabU9uYV
DUJCeevNCK5A7gKsZkOqdRiUln9pA8dFsLdObOewMuWzTqkFd0kuoS9r/x8cF6LttGmsW0UYLHHd
uaQDMVWQ++09kruhR1TPDbWk//w9FgCtJn3C/GBBpzaowSJ4xkTpzSS3PfsxvGWhtcuFLBNar6Xn
VY6xGeIcup2VNv1mtpKCFJyIW4rSmHpPNgVhXdYf0d+uGMFwheVdmb0eWvBrM+aaED7bpfwlkdQY
Qo2Bs6LoUbAAe8DjFwIG7TtBa7H+qwK+02zqzLNcYPWhOsl7kW8MzjWTQuuLwqcZFdMcDA+gxIHz
YiNkzcL8tfm7IlpWGEaAfnmSYhz2n2/Xz9cvC2LBzCXZrthOqpUjPnQOLGDsxgn1UHpgkXUqSERj
QZmS5EcPx+M8IUZm2R3AR7Vo0Ol4kH3szIDAyvEUVxL7T9WmYTnQcZFkCauOBqywZhp1p9lTca6C
cxVcZhgHTLkDxxtcxiidMOVn+YYElZxarowHYnWwKpbPgOdj9pLqmuBSDtzc1ev9A3kBLmt9vM8L
K61t9kPavXvOgw1q2je/EsXZMUGtuLzNJyDZH+1dYyrX/xrnl7M7y1s6niFTZzyhLbjovfRwQ6+/
Led/xRR0ww5Fa64G8mP8Q2ASGBHXXta/BbQWGL0tfgSa4HJOF+HVQbVH1l9loK4Kc0nRuzchYDHI
30SawAF80KC0dp4toAjeE09UOSwahjH1GXzFz1wVwXP0yGP/I04bdVzPF5cJCRAUJeGh7/PZz/TN
l8hwyG5Wi/LusSz/1K7pweRJU8uKIUdnP1nub0ScHO70g11JILcKJxAoJnRlbwQMs4d0VSqnr6uZ
SyexDryIYL5Q1W58E2s6WNhGmImet58HhUK80h1NSeUHXvJ8hmxT9n652xoQNPtddujPN1uqLvdD
Mvz+r5IxJCDWSWi2KYsaG82r5VqTWQAxA9K6qFVvJOr1gkmQlDLhQ2PLl8XC7aG4JmtPD7BZsRxI
i6xJGU+GAW0kJSnb8nPSyvKpePagV9CGZ1NfTsYblxSLFSjwQn0RxUrnzP6RCafyJmXIwzmDeoYD
A719LhG5OB4XdjoUxVbaHY0JKDV2ioLt5eRSdjTo/ewmgPZ7pEBWVxSv+ZCS9a8f3uXRYM8Wr6p9
W0uDweLCLPLM4lA/ph+Zur8kDBVlYaqD4ENJKIRwse0VBRuC8F+6LeTIA3KqfJ3tRktDJ3670u1c
Zq+vjsnkrcT2tBOBe3P8/0CE5VVl7WUMYQw+MA/zEW5ZUA5jKPnWWQDcLpfb37bqTKznfaG+XhdV
+9vQrUYtyjXqmZVwDbXwPOBPqu9057iFEOPZsZsDTom52+aWsKQRgvYBjGo2BoJpJFR4K7pxMLlm
IPHv7Rf2VYYKhteBHH3Nta4bzEvYRCjN1GtdNqZ4z6umaRkcQbmzsz9b4EMXUn4WAThogkGDRuFO
awOHGIMEww73p1XdrJZvnziEFSQjdASnUXb43RxX9dLLv7YqSGGKGxM/w1fMoOBV+G9Iw4vpm4LP
qt9LiaJxb0VfRBbHVZil1EymR1/U2NEdeBfEj9Xwm4PciMdC+bRLUtQkWhhAf9qLSlqMXiHmhp1L
lKJvwZIJxsm6YiVTt7btE6Wv1DWddfirXqbZkRI9/KaIHk480Qd1NWHeVc+jYSJXLn+VDZCSAWBi
fxx8Y7Oju74unBZSrp9aK8vwMOGGF1xVtk7OOqNHOKUtEet/lKwP6NCbehelnSS22+XJN6S6LoWs
ErvVlXQImoaqnEMzqEJxCm1A8xeFe9WCJGEtkXUoQh/Nd+uDk7ZlfMPg/qsWpTChMh2EMAx8ewTZ
dAlX/HMFqCnkZ5CGgmDOKGCQCaJgF0enOaKgMqIxtmtH5ek987iHon6B0DiHW/mBqCWbAtx50B60
wHmmmUAfncbVqeyt1pv0ZdvslV1gZsfr+6P79tPv3FcL4V1/LhQukp6/9t0JLCRqK9La/phJiEY3
JLCANWSoA3yFsySholkUs7K8Ti+SCZj+//yHzUDNb8aB8RLtObBER85pDfARTAmTxn3GAUTTpcF5
P5qJO8flcbIzupS2FAkUTjd+X/pq2R/xPcsl69r/JUf3AePu5MyVrYkP+3/FbW8LLANqXJfmWMz8
AEEAB/jxdl0rJBcKi5gYZJvLiiji/I0l2XMMiFkMPVRUWoEQUpkPaFgsachwf24eF+lChTUqF9gA
i4aujWQ3yg7IvcF/ejYpPyY4AfLo7Blub+nT4mdPG4LNdzPj9XlGWQGCsA++KhS5aN7CbgkWhnAV
DdlhuzmG/lkKBYqQMt+l5S1PoCNCkCQio/GzuFmUAaOoS1C3m1w/gBdX+rkUHsrp+zVSDprXtpeQ
DxkeN4K+xu52Y744CUUk3Bw8vWtJLhSnk2iJNzr62fcgD88gMP3Vx1/y3KrWjodfuFft4YA2ppG4
KT0xV9heJWPqCHvAxRcq9l8mc3jAVThwFz/ve9clJqcCoAjAQm8ksUBYOjwb1PXkzwehfmQ2I7v6
SodZAfV2jh4xWA+ph06yNrXhm6C+uZ+ySFcQgf+v7jB/vR6EUSv0VHXhczbuW+ugl9PA3mDQSGeM
wjSA7i08yA2xcS/w5WuW8ePCW6dHjUOhdZolmb/eBgfg4c8LpYKABlMXW+KnChF3VGfCn7NIyxW7
OuEVtpz/N4S4RMVGhPCCBe3ubP4qvtp5j5XzGdWSstxIt4kpwikNXdC2xfUNBLDUmaTO24QhwRZS
O/+xk50DCzIwCuOuYIwydOES7JZOcI0rMqKX5KcM8lMiL79bn7FszjI5iiws7tbXB0shqPA7lDIj
iM859N8G/V+AJsXMOqXuFowgM2dpxmd7gitrKw+ROMQmWhPrUZcVGttVFzsFrbFhN2zj/XlhNRVi
6wLLPPU66EO0Cde7RGrmuYIr3/aOUOGOoP4iHw6r/HYE0TtmPx/OHdDuvm1D1CbIBO8nFY14tArF
1xkBpl3R4pNq4UcVgZzomnSWoGj4UXVIWY2FYYqYZISrnu9mEq0dEPuwAv039NC9VXTeeAkUqF0y
Ghk951rQKLFQfNGcLA/VF5d8dj/w403856i5EQhlPRx1o/kh01DsM5pTi0Zi0rOiwB2RuFQKrYPv
dfF9ed0KdBik1zJfCdZ3Rz+WPAt2z+5SizQMsrrcRMYDyCbRL67QBBJVacak3fbmBltSpaDSiGHP
JAbMXR+4w5kuvzdFh0l3b8BIWoMtAkoNrJcDIFa8ZJAsVW5AizRXJBU+CVVeiAf+90EHaJLOO+N5
1DkNpEcaYwe0oVoDbKkDsOR08aALFSxb3ckuBnCDzfkH+XI5nMseBkRVnP7mm2ffWEKJtOtMx4P4
8qKKFLz9kdVHaInt/3Dw99Hb6gKBC99QbEcFWUSJul3btzvLvd1smk/evhQoKhfNYfMH7JTkP7ze
DdofWA9UMlV2BvdbY3SV4NC/bolpk5JXZ8Z9zLmepCD5PtL89mOdAYtFh4w0BzIjWMTeoF73r16G
iqTswwLRRwhdMOhV7Vpf8abBrY/0cbWlm/11QjgJSygtb7BgSo07xQR84Ngz/yVrGdzK/RqJj1ws
W/OdGFrRnOqRm4DXOMTDdHghBQW5Goy9nv1g/HQeW1keI0epn5dz0C3MhUcU5FdttKOZ131tA231
V4j1zW4EapEDO8cu+AyTSN/Wm2H45RLJyTUUVB1TM+5Kz7A6LEP7B5EQOxObFDf0gZpfbJohIALm
AvWdIz6PWrdJep89pEjio3fPjnP8Bmk7/r34bXKGHJGklmeC4t5DOVLp6w4hyoBAgwMzjG2tooVt
jy9CfurY44okIKPvPrgihaAXSAL0z4hb40vIaSK3DOTxlLnkzKC585WzxFdqRRF7VcMCVursyR40
E+Ibdy04jdUCpG9kqI6EYNE+JRd5hPuPLPcZ2K1PM2+eSHiKgSrtFpYWRiX5WasbjbYgFvXYGfuy
MiDUHjwTYvoO8V5E/CQZ0fS9wi/VQnX1txTXirJ2lqffF6gisxvodSpRApn9gmvvFqfo/EG4oXu2
dIMA9qRllBI+byGKl2VlXj5UjSGI8uW2oBwDfx97M6F+CpXe6Xso50DPIdUDYR4vVzjwY2e39Tsu
Jasxnq4ZHreYER6biYnc4KjoM6EpUFQgluBOkMjJM3S4MHkc/JD8t1JcGzuTY2Z0wHsBrUN7Hd2D
iRlpithcwM04RtCPpXKhWDIYM9vtW0zuG8NSDtDibsMLyBfjSZ96GrLOz7W4GTK9W19pyp/6duFv
eRxbYW1QIQ63PMmLSmVhlRrhvUsZ6dInBGjgTGGbvuH02yNP9mFymzDpSPlhqLbkT31fEuXMCUb0
k6mGhN9Gf27CyS51+CBOQy+xXCgOgo51tAvg/gXcXDKM7npOlhvcjhlTGB1LFrfXNQvttwGcvx36
tY0kbqH63C7Ud6wBPhP7pijOiccPtOaHWWM61C1UZ7LJTXWVYfnNEEflmsthIZujjjXYH0IZI0U9
l9wYnnQChbchW9GZx3tMjSmPzMrqDHAmybmc8CqJG+ID+9fq1/LfzApQlKK1F9Z/xc8y5n8JT+Ji
K7YcyZRFDVRlE+4KEPwJ4DId2D7dk+XvIgUTpwINQK7gvrgYyvNDOx89uda2wNEW+0OB2dGkFOK4
QmpBUiePs+R1x4FsqkB0aQWS97YCRXApIF2jH4s1Vb6P7N/zVq2R/K76BrX1waZ3psubLeLe8yWl
JToyzPOanupMy6WhpfLX1WZVXpAGWaetSo/pn/W11xdKiYiFU4pQuXJAGAX9h7mpHq37f3WAJtGn
8jPyIKt5iktchRzMWgVcXf33DoeETruWcXrnCskrkyUG9CnfFB0Defss0CFnejsBh0pKZc6XeXP+
L+vkfiofiVRdkBG1Wr5cDILIECkl+FmHbylOs9io0XWvDK1SiFGfR7uyXdzKO0NU+2G9lyokQdu2
CsoSfPW2DIERS2hHGTTvQLApa3C4ssjql4NLO90wan3LubildnOnrPdc9QpCLnvFNcPbCJXUBueX
ixyzbIVgk7XuAcnvvh8bL7CRzIJxjSs45r4k2xZ8+3Yl0HtluSuu025vJvVP5g9tlCmhdNUaJk/1
fEp7xQTW5wrAqsA+nNRUgE/s/6Vk1UFm/kf2x6tJCriJ9nwwpd7Tz3v/ZZkrlYSkA7rZ9k3CJy2j
IYaQg3Lk9tBbrOmODBtjUsDk7eISUsVFZmhaPY08HT4JByR1PgXg1kR3DeRbeVVI0yff/fCz54z+
popLhthfJTkgRQwDiL97XAj9HZFdvvfOt6mKIPp9X35xJqJU/Uv7dHFo3F42YhFqR0+ooZ1R4EUl
1HhIMR3f8FmEsiq6Hdiu1cSJTEcM2gQ3pziWIQHTklC6IkSm6gBBmDiDl/PYTUigGH/Z3SLYsKun
gTGUTrAew/A4u5dk9mUSHa7JYG/RvIbeOBxAnVEUy69elVRFz0bb+oSHRr4CpSfJnAQsIzMYePDY
b5IljJb16mtIXqW9AIPhxIZwA2EaGQgXrUc7q6re0g5HfgA5nCC+YGD6ngLhz3n7BadXhYiC1QIT
RliOUdcugE0TrxzNZVcyhbXxyqh86zttv5wJXYd3nn52I1zW1evS0b0jSk2GfP9MoHdypj2ucanB
42u9gNjEzYrTfbCNEh+uULx7ZSOcRaPGQcIUfrn7Jd0oEdTEAVWPLFNOegbEHWwo2cXk7vO5IRPl
EL1khap1vIZROpLQzOLBL076EuSv+jRrihYbBzSW9wqfaLpaDesddyPamvs5OuVw+1jdyNWwBqBB
acoNt+L01oxKmIbwGukwF+sV2kKRhLpj9mvJNsiw4wHcU9Q8HHiugffOAcpLH+w+bgHQPew962g0
g3M+k4D8NLUTwpZReFe/tDnHb2F8tM9Skj7GPCcG6oBxjSnCaioy49CtMHa5aVPSOQIBL7EKCRee
4s8Vn64V0Lv8L6Uy+Vs6jyJn0L1xY4N/JCGb519oa0kWJtHfiAsn/KDM0c/E8pzmg5TFqL+em9bQ
ssZAg6debiXfnbbCbIhA+GspCtQAOu8u833AZKE3YwdRfCefGhJPJ6kbnj9/I8//ngDaPGo1rGQf
FPAbAQJbeHmO5L8KMfVtqB/+I52tuvxkyA3OwERIQg+iSqg2FkAGgJuQKL3NQU2HuhgdYbBU1LOG
WzZrvGNk7dK3TB9ZqIgdfHmWvpYIHFMGL2+QYKaTmDbTc/9lXo+yJW+mqYQmT3JkSWEdvPftXBuw
DScjap3k3jFg0usIiHjAFMJLNoI0cbPhKoZOvYmwvzFLv3OhfiVMhshV9zgjZpNeT+RFvEvO6QjW
6PQbU948NVACz+WQjYpE0QbdULa25StrzXvcaFirFhZKwgGQknSrCwzMGxK3WL+n9xS6IHkFs+Fm
KIVs3VqGSowfyp1hhmi7DfV+9QxX6fP77ZFCeeazgCs3BxaysOOGe1+NyaC3EIAbehXay+l6sogN
vjAegNk9T3rpdHTzi3kAWKc7eQNyH86ZOCWsz9XB1TVJIN0ErRcZ0kHHKP4Ssdw4G/B1+5NPJFC1
7HEdA/xsImDpy75fsnumUDVuPp4RTlkp0ovakygRHZhlY1dWJ/55+aWlBzMGBC658bSeYKFemsBY
hyWoujeBlcnrDFZla7SvBI2t3JVi+Z3MwYE53L/AzRARSZD+zVrHHH8ur7ObA4F9K+l0WXP6bVUK
uiaBHS+qKdXctlQgUhgaUxpQ1SPFCIAz8t4Upo7s+ofPe0BDLZYzStGhO75zoHXnrt22Uhbg1LW0
hpnZUBl7RwBr2KISHapzliqCL8NE0CHvITQfdFKggoNjSsOayRHrdz6Ywvwuhg+r4yfrKkincU0z
7DRYGR29/5hZR1pwRr/UPfRgdGVMO49aCyKkcPb4oTemWNq2XJRpb1RpCHWJsn6hLbKAkEqYC0K9
FqpM4ARtWkK/Fy3/r3GzinnwXbsmRgggzGjanF1/4pvAKFVA4NJLsxF9wcEG8OaYURUssh7HxeV+
Ly68pfYrhnZdjqOgAlyfPF7Rv881Povee56RniaEsvdTqQnUCzC2ETJxLOiIP1ZxyQ5ZD6LukCON
kTjJ1jPE/+dGySQNw9BDC/fZ7Y7buEd+UFs1aZXR1WIuwv9pM8fg5c5Jtcw44UK7EV1KGeOwFcCo
in0yGl8AQTsifmE47DQpaH72awgUXJkS8g3yEMs8kixl01JekYIs3OTrNxwsEKNNzJpAgFtGd4Wr
wKg9uE039wBdtX9czFD3C3DQ2yLRfhQl8JvQbEsztEm5DQvLbd5Z5kNZGog5ANSP9P2JSubYE1YD
pVnJ9U19jwvD6b1NfviLPgu/v1u2Q/SFmr571PqfFsF/FtiZyd/Pndldhj03kGRDdE/hVXTIER+f
Q8ldv9BIoCr9iPI9/Ey5mbbTCbbVO+TR8rBPhqgNDBVboudlrNYiYRpz8qgc9U7AOQH6GGIHm9kz
niGIHV+2z+4a+2qH66ld+iBnlQa56Gw9XjedKn9EH9PCgnr+3J/KFkvlGvfH7nYP55vTLHsHWv8s
1DYF/vkWUTL44n+TFqyIbkkow6r4UbQkKyc5a+qyH63YBMKvPHsHvJeFssvbFvhuocwHmQ3YcUq0
lGwQATkRgciJFjEeOfejecIwcdk2j+btbV6UnsN2U3li3hlotJv1L7YE6iD0hWK4DM/C9Q9AgEqv
D97VtoJgdHGk64wyeKo38QmoR/+IYgpNKHiFTx/Chy7KG/2qXGeAfSOatEXiSVFCsQGf+F4Yeqy9
F3Yf4qR7/mAr7L14/pItlkXT9PGLbXNt7Is8QO8TcbrlbSWs1rVr4cXeoJVMtmY777PpkmNgfJOQ
tddDCReuUlJq9nAPEI1AHi0SItiWLwrsWw+hV/SKBnf7o+0+5n8xVbu4JCdMWYdU/9494Y5mQ01n
taYhmYTBQMspblngjN8CkMmDFH0u5utLfEnVi7rExP9EC7vG+FAu0rkEFa+SU10P7Su+KwBytAgp
ur2xIfLNCnuBPJ27/Bt4KJDHR2yoFqtQzI2+9JuCvI7p1KrqHNXyVc2jU1roJ6Zg0VhWGiJ5mJWU
e66OqxcRjVI6sQacoGBiKv8a0GPYbYHgoJ4n7/3QLxEjYdDMpES1X9/Wz4MjRgQpeGfzKdb6fuQg
WdmpJf5MlPzYbFWPBoII8Jbro8+ONIHbJTQxGllERBod9lNuGKYpT/x0SrYPR6jDmlPwY2JPfVDU
YTa/XxETZFCaAW1AkscL4cCdUnj93DuJcl+KZLjMtMdYRcx16zMIoXFPnZC/qRjtpW+QgZaqCPhe
+4ZD1esM3DQAy+TpPeVuIPO3edUhh9Wjp7wbyvW93RgscmZhACmBHq8QaFsajkBeWL5O32Zqzg4R
E2Lhb5T8w21zM3eD/MYJHI5sem2d7g9BaIngzXoRM8mG01uVDrCuKszQsiHqJZ9Vvqqx5REH3ob9
UzTE6IUTcND00ofMZUYg26RwM7yyFCTydR8WLmU8FpHStXiWPDROvWi4v7NpLdWJXaZlIqbw508Y
M+3jDdKllpclzB7l2ge4C9cbxsFgnYtyfGjPEHQtkTpMLgLJo+FKWKtgZ4o8TdLOjUjrASTUuoEP
Vmm0y6CrHqMIIM+0AbynHcivtlhMuJn36LUFJnpCh1adb+kdo5kbpTvE2tv8GOPt4km/OAku4tO+
ySWvcVfVu49SOdfZgIAGLhWKMfQTZbFx5GkGsKSUpGkgduwbz/ILnRYuE+5ioJ5sVeAWXFcxl0tf
RfOzUW6502DbsipYiKh3yRMVuGhb7Uccl4ij8B72mMJICyZOKUuNj6Godbg3+AbiymzatNaac63B
jghiL8627PUw9/BSCv+67h17YiY4Vd7uG23uHPjN3DtuA/ybqsk33GtxbhMUqHhpvFsE2K5Bkg76
FA9mDIVVEL5mbqYJuDw4yycyTiljUNNNb3/fFhH+Syyt+PJfP60N2LNArPFWRmoefiQ6hZebKuHF
crCxT2q82NDOEqTiO3A/btHeruQBr28hfWFeVaCm2IrOaZJtsnSvBHbiobZdIK9V+W0eU8WT4Gpa
W/Kr1Ugwo+n3Q8EkDWLoHkWDf3iDElrhNxb8WkiYx0tBaKXpYu/xyxgdXS0PRc16/D2+GUy4BEVz
QFSnWL8g1lCbRgomwnvq4e18TcT/aFOK3z5MILR6o1tVf/YvywXbe6Y8Q6m7zWuYBi3SPn0pTjUp
lJTT9nGOIsdwB+yXiDoCJeqQ5oVRteKuJopRRaLynroZPjuUY9n+kKUFONDnJKs7RXXTsZA/O2pB
QJCRUFW7J2xoAFhg4CLlrZEEnKRs1FaqfqE2kG2E0w/cMiO/8pDSndFcEJLg+WhzXNP+YxJQgSQi
vmd65d6fI4VbDzBn9EWK1h7mti13GdrEzDvpcry6kFyT/lIyLz5haOrhXO698pQSG+9lIpHDx/jF
xJbE5UHTgs5QwEsRdxVuo3hXA3Bpq6Mu/Xm5nwCN+rx88PTa0TYJlQ15w6tr44aiDkKT1sXPMYoj
6XzzKRd1Np1PN84v5wO68mac/Fc/tiOQbPVK0axt99nXnUiDa8BnDI+cAHBUGMOSfwXrRaw91F5R
4IPdLIKZw1fk8o0tc62ZNmm6Lm/sDCZiSqkf7TamTvlg2lIg0x6kTD4cp/to0iVhC/EYrm6lkg/B
S4wRpSMo9uuDFlkuH+QXQ5GHxVNxhoLg89y87f01ER79YEL3sveBCihX4mBLj9xGa+8DEexejwgR
D6+RdYdgSyBes62uMK0OCI/IRJ1oH8DrpbppMoU+X8kTRWVgCx4NugnZqHaOKFXox/7f2dy4ToYT
Dilv4Gw0QYBrMLYOx8HQBpyGhEkgg10MDY7Rv0gCQj6jzi4gQlrakhGsC6wE0lU+su2MBrYBsWaz
EJJPg+Qd7MAkPOVIjfeRaeWtR2eYGiYFg3US2+OVbZqXmmcleXtLaFfIzIFffrud4AuoeCEmXGtk
eeZ8MokqJDMne109FgzW1djgf0dv6g+PqOoMLZhEpKgo8xSWjgKtr8GahSq5MYhakwDUQZ0gn4tT
Nu04tyOttR+DFU4vWCOj1AO+Zf0roZKMriqNtnByxkEwujmMDx2Udm3SSMTeuHg77pOfUNoselyi
ZVqP9Vz5MFL/us13S9fpIUtsFvMtwBsFzYZSbjflT/iXME9qanEdLZmJOXznlhry8qz6//AugHt8
Ea+VoPoRiJ1xiOb+ADE4XKFADMl3nEUIvfjWx+t/9jn2ViT9lLbHMrPkatWOKauCpXPWR/x4DB89
5jNOeoMhJoivZ5hekJjVoaHXMEu0Q99wTmq6TM9S+ph1rPZBREMc/uTc5o5BUlvPychE6Rp+u1kj
QCs9OasFPz4bAKLWg77/49cvOeoAT7QXW4hzHcBHFaEXhRsnZq6tjXGkwMKAJRmqEn6qX1FhuyL5
lAawgAlmEEhmlDva9zDuocWXQXN77QFrQd234WZEj4l1jBCUeK+dgA+edUSF5MV8ZXemQf00mzu7
AKfTbGPfg6v+121ysIq6kilG/Nf26OvJd8+3tJdsw+R86+yqow0iRi29+GiL9F5WZV+jhI9DE50X
gxQffK1sGY49YODtPPIyP1YWrEsPWQ77NjjI0ARWizwTruvDRTH1zxCUSfAHHpA9TMTe6KSZYCFU
KiQp7gT4/P6zxbhfIOuXCCpLFl32EbVbmVm4lqxvb4w7Oaks8okTqPqtUkO8GCRTJmwoX9emZUI/
AWS9VzDvHOaEoUQsGS25Lbsn7VCFM5mOBDBnCjqy+2+lANWXeeVHd5eotYDLArOnwAK2cqENwMIN
AbJjyJ1cE3UGOPcwENi2unqZrY1V65/CAh1rEKb2nRSZ2q9M9Wnn/hff9ZJz2iVn7oTbCmfHVW3P
0qXYQN2Grkt8z12aL8H6qFlOTOyRUnJB48LGXEHCSN7kLYihdE7y4uuI1zqp1pAS49Wwzkb/nJQO
EKDy281VEUMKH0sdAfgXZExqHnJphWnRI6OhcVDpLpcQ6OzcFNP1lDkyjJ7N6ho1ATJy2b3XvlfY
lGgPdxZioDlSG+OhyXKdXYCaAkRkgQmL9aAt2genbPEp13S5ghu9jcg38cFRTgiXSXVyJ7hmcdbk
QQOxOoVdBf2QfoONMCOA8eQnan9+i2G0UDR0PSm51NTE4TzWBKs4MAgFsh5wuSAQHwkWuhHUiv6d
5ad3+2C2Hbg+uGYKNWxynT6feCbflk9lv8JpvX9mkMjX3K4S9Fp02TwnwXdBFEAz2zy5Xp7M0nnD
4Eb/Uqv7W5aczqyBltwk7quNiViUN/eu1ATu+0jnxfphHvLCLBlpjJ5qV7XqH12F9I/4ZeoYlCrI
AI/jDxQrzci3faifbdcjh+gJzRe76zslKkQyQD0/kfZME7VdcrSikwKsAuumumfZVqwQVY45LDWV
JK3S2/IsFMLrPcRoQkcPbQMLd2jqXXm/FKmyXUPxOJuQPWTn9GrGLCVjT+fQj0MLOwRtVXVHi/3j
dBiB21SnPq1k6QjJhpkff6gVoJ1tydtcXTd7b+j0jiJU2Nay7VpjnG8QVSdaluw3UF1xIWPwlo2l
NNCllDsNFvW3aR7Bc8v++rhPjTsQvBcnGY0JSHzuKM3+teN3Xy9oxKeQXFvNC0IWEyxNKqePFb3N
vi9qPDhEaYpzNo7qu7piIuMkwQBdw8sXDJXYFPolIZaCrvJRIwCnieU1ONayjBvdRc6UPZmYjDr7
z14B0jDdDewUrlYQP0B1o0a992cUXwUqgBgDIk7xgA3ysvBR4oQvmiAig1EUX2/F4N47RMmGZ+6J
A0+W0N2/atFC+JWAOtmlNULaRdzgLLiFyQMiHoKfJimHQOPBsIrEllic5RctMGfMBnF4CGnTTYqB
ZGz2eVg7AvOS5YFkYJK3uVxIjknJkg6lLP/uAi/VSbCLKYGNoA3SS/JJTh0MW8kierQgPU+52Rh3
m8bA7pWwFgM7lcIP0Bxoua2gZCOe1UaCNvAEIXhoWak7eRXAe8ui2kYdcT9tw1BFDVJHbgNGlf5Q
t8+1kIOgVrKM/Q3pPIjnfZc3hD9Ngiua5mXIndtFmIrRX3LDwdIbhljgAR2oLypumLFNkim3oUKn
sxop9WUeJa/Ta9LGyij7QjIVNUGnj+LY740I3ErFU5O9zB5G+vYH9FoBZlPwWVydcLjUh2PCUOt7
aRimrPEchkp1OU2Heh7dh/cKK3ZsXOZU+dSjQuzDUOgpd5e4YJiYa1uCNz1L/I5y4dvgGth3+goi
V1mgM1A8P5ivrXYG6dl0FViY8doKyIcAmqyJJROoxKPjsQjf15rPy3zyVTRzX2AbqwBoYc5qGPuv
W8e+7Y3YakYRbrOLdXXECDW8TKZslUS+sjFts+mHOIxDoaZf1WSDsOdaEPnptw1uslrwObuatuBK
BcbFigGu+M7xLUhq3OqZTL5ZDa8wZUKptL1A5ldLAH1TChd8B+nTrPzA0pYTM9/R/gBz7EzkL/oh
FWswS/WtYwYetSGrejFDrKm9Xecupu25GnRUpR8a+vVndofj2RQxO0douq0OssIz/L2Pw6hyZc9d
gifd3TqDgMy8I8S0gDgRt1oCSNYnYQzPKA2zLhYxi6GVx/GCX7icj3CMSMgUtgJ0b/TiOPUAnFmj
fW+47obbHsj2uc+oP0e4UzlWCpfQi4iuW45cqtMusvA3lTpnDxEiDYM5dtj0hG4JVLpukMfWmT4D
ijo8PfwAfDLdi6XrPI8JIIE2e4nQriPWOk0iXrIgAWq40OVT+M1CCNC3fVmbGHSUEm8GIfE/eXui
abetwGKgKU+dWUs3Q4OXILTLf2PkKfNsLXKZvmtskpU9hnKN0UXdbUoqmigsKA5iRPZC1Gl3jmWI
kb+QqViHXLSuJPF1R2ORCTbG4w7ngsG4VJ00/TpWnDIQcpcKM0a6nP2RjNJqIinIdlrDAT4IFHtO
MMzd67nrRrXIIDF3eaKY5gcfG3XKMjyeLD7MO0WF9BHvJMrm9Th/U+7EGu/mWlCrrMu+8L8mGrh8
SlDGY5wMpxWQQ5p45o90rmtLv5YDBxFxenNhnRqJrf0lMJcERGMSjruT7VIcLVcOPs/vlrc5BVMb
6b1e6nlTfdy1/2kW1XspRkojy9DaZrWj9+6Ckx6Dchh2bd97n9g+mxrYYIDoWRY1xM1NwkWKFB4B
Ieo+WTGRnk9ug3a1tUcvCiCNcgzqf2Jw0410cdA4q/f7da9QpFQXkgrBCLOccR2r8dYbwbmHiSmU
YLFwqVWnWdVTff6pbqtiV/53OREp4LkzCZ9Ms9bW+tIw5rnyujY39HIzYhCtkfaiutn7GaNPjGYs
jfTbdFNfoUXQp1OUVJ83lRKLsnhZFsuJJALsrdwnbada368Gwb4xjtTilb9YJM+lJFd7Ixe79yCC
DrZmg/9dRpjUYX/Hj0INn1wbqmaQ6190EgYdvIsG60QkWAgf7CWk83lvgoB5h8A67M9Mxc7EpiJU
UCcL0V5MIEB1PqM4HnnJA+7nVuP3DSOOH8uPxAC3YFLRbTWT163oHQnA3Mvuy9skMzSlLMiJXEEO
v4UBMMkWNwXAk2soKU+JlShe5Z4Z644BS8Dv+B9NiPLo+LqGQsl9LT1yyXVPiQzpsMxehmrkyVAg
UvG+EwOkUwLv3BlQp2GZRQQjonByH5iV/FfSmPv/hzHds8aPgMGPZkv/9/bqUh2ClKEYMmPnOofY
qmHtlWxH4mU4A9TmJcUS2goK49y3dDZsQ4LXj9ltBMD9YEKsFUwM4Qd3hl7a5TDFuJHHG2s15noz
96egVq2Ql63qE7610pccLxOrrVvXPx83mFLto/QYvmoUCEZxvYvN+/CulVbQDX29x5kIyB831sTD
nkPw+p+kUF/BLdV8zohTVhMYrYAzcBU3BGF4U/1DzsmUN++d+J4qieXYJ3X2ku8KaBx7HaX5R1/P
hS2YZo2QbP35ftutaKxxRXjPc3cxhLnd2BC7jzb5PrO5lFA3VV5HVSwhGFhgB2VSz5F7S0ED06Og
08RhFZOD+7psLcvMpZ2gUIIclkI/1aMWDKRbcf1xORcJxzqHZxZKDWkYl34ieyfDhinPtu+h2lpM
dXu58DhbNBlomJBIGZyDpPcv35yryyECgnnZ2JhbsJwRS5NqiB1PCZ07s0Htvbn5vMnWr5CfK02t
DfbVB27DAMGqizri8QDeqgwX/SeXnSg6ukJzSrH/wLTplM1Y2kUq0PBIgrAvLfrk5va0Fb1gHIPV
hMQiW1n3+/Lw5x1ZV9MWGK10BRxeqEYsCXppqIexwVoMeUTL+VUpldH7nyAjqMDVRVDkVd1hyDCC
wic/PN7tb4BJYxJYy1Q+dLTo+OKKgzEcnxvZ8cYU/uEQZeAqi32HRGhwkG5vA6OVRMJiiiWm2KXS
Pr2tUeO7V0X/S8ZIvI5982R2rCMKp4rhB9Fh/RIiX4fqxn10K4ZUFJ+3aVd/kKlPEPIa+pGd15vD
dkBfcVxopcRHvg00FZJGEj4Fgm/OBMM8mgWv7xSvB04Rf74bwtkocbJudax4Oox0uRAKrH7AwsOP
/eTcyj7tmVpcqZIMKFoUo7GrB/ZSH0A3zwkWON1drH22oNufy7W1LRwSCEEWQok6T8dpPl5PySBd
vabzXorTWKiA8oDxn9T7pprTe2IvPmc7ORLYxSQWckrPlww8RtNS5aCwdf/gn1X5cSQ1/NLJi8e/
6+Amu//s31Ma6N43iev56WFQY9n6mQ5psR/bhsK7zdfGX1ixetW25SdcJWGtQjgRv+UN6GRuPxyW
WmM2CRDE0Jyiza8TEkvWlOq5l2o8w+KIVakdcVA6Ft7lBMcIOnxXpwtlFXqSLRD08AAl+LyQRO+y
lmBaEl7xCEhLTLq1fRNimRFMd/MgOReUTz/d3gk/biufPgqkbAQh8CDM223gLN0jq1WWeugSLN0s
zeN5uZFYCkWfANnpdPEXB+GV7tg/U0lBzY239CTXwrB/p6A4lPxRANOjWHc5GQTGcRaGPv0pPcaj
5UoWT3GwtojJ8izhJptkfjC6m0z577HwrX6VOspgpGZBfDsWbRveOI8u104EKdul/Rs6knTd0+vQ
FaL3G4r1+sIh7eVUFz05zfJGMlWou3C9cE6VTjJ7w8FA86HMhu6gVnAY6rQS+XJggM2W1+GDEHGH
KO3j2IkFcenSuID8d9oBx6MGNQz1istSdKziTCzctKS0JPYFXTNexX6rGUGsLJ3T/i83eP5+uxB2
qdT13MqtrormZDJReb8S+8Xy1/029s+MRJr2rCXxT8fE+xxZ4kIVPBdz2VQEJBGb0iQPIKZKW/fg
4cog2aiPXc+bnKwQbzGA+nd4tKy8WfRKJleRXqgvBv4iTVgPD6h2ncJ+DKu5VGYbKoT6td3wcORr
Ko5xMOkQrwaI1Mxk1hqOq5nqojCBXgPKF/PAI8yoghQDE22g9QSJCG477BME50YxZXF0vpHDUpzR
exwgrl0LFoxAXeQBhVlb/kDGOJ5Fk3cRRmngmgvilowfqzr0L/VkNECSqw5mU/zoXE7ffV/RgYN+
494wUHJ+NK/Vhx2cjyxnsL5NhfXqB9Gd7jIRcrdkOnlb6rwbk0ajwNAovPtd+5zBLLVIrwxz9vOJ
iHwWnkFliZKVNTnlxCgX6BIyvXtKB1+ikVKkkmhRlG9HaD3wCIpyTA6nEVc1wrvzY1b85xeDL+p+
ZwxrxK6rK40eM6hz2A9/nDnawU4XaY1cXXzHsjaRJdEUH/KCQwOLoFpcllx7FE2xeFE44/275NZx
/rGMWA25RGnmiN4i3r5omYFsYEpi75LWg3TrbKHg0fGxzFllHXysprxyNc7KuBGxR1GbJ0H7O/iH
nVz8Jw1JAt2j6myCiALwAPvja1qeApyvgMaI+riHxqmb55ZGfxQaAGEtPFKGoAq+gwlGUiKa3gTF
Uq25GKTjrysHxP/Eccq1btYysxuhLU8qcEP71WzyUf54Lr4o/qy6CLPh1E3Jp83cv1Uk3+oy2jTO
MoMQPDAwu14gKOg28SCplc3x3D2C9sfLIZWQ3ncJK/x7ftEs0u3EGtH272w0kbWF5bf1B7Ubc8pk
O5K3N/DblwyPwz3SL1uPjnuJgaDkz6CWkMtt14iOSlLyi14EB0yRm03fgTb8buq03IsyjeRiiB+t
ZFv8z4CY2MQ9BuI6vF0CxrlK1ulS4kFCcX272IcwJsjj/QyUXCo+7eSHO538vES0CV0tXkTTzv8E
T+vL/Ui/aDZr6L/FKXwyJKA6oZnjNRTPIomYH2HwqpWnch3Ath88JQlX0ITPa3/zUYlZFv2Nawpz
z73Gt1PaP+K2uWxpk4NVirSb6KgmtIFEIWdYhG6CkOd3dUPFrzpYFCuL6ALvj3yPFxe7s1YcNWJP
SuOXDlese9zzuH96m+V3BESOAigbBxsjeDY1qwRnzemc0W0w87/hUrCaLBNADFb5uHD2QnMSCnSE
EXlqljBqmTLsdltEGBmg3OhEzWwYTk+jN1e0uXOSQKehXFJlzG3o+EXi3xyHDxj9Jd8RQXDpZQ65
/GMZiKG1Kk0eo5yUchWG3FNGlB93bh8mcO2iEkqpg4XbrLysIFmO+5NXBkcR8P9+7hUnDmuU1Ywt
r30CfNQOygUbGvtBksdGYwknZooEIZjsCqeNftfcBkdTU2QprLZV5DI/OA9PslYvuVz4yPIc744C
vjSb8VmfXaERnyZXgUGRCkCwkLIqFg7HvZ6uYoilRAm1mfAJp9fUEWoN2g1m9mrU7qIx+7GsRvpj
nxlxcHQ/dDbgNxqqXSWoqJBSRN0QYRgK7YSDV0eES5ngq1cr2Lvj1XdWCTv7eFR3+JCZUyfKy4Dl
UfCPVFnRTyqPnHcAYDYZoNTtJgtwL8lQsfr2aznFGGA5Rs6qXG5MpoA2Uj5IaYk/d2GvLsbN6hde
ohVhhG7kqBMFeQI5tjK7kzopAYU0kD+bKPRcV4Wr/KMnQcMwrtxqcR9k3+V/hWYz0z1BU66AiezP
Mb9jSGSwrtSXLjP256GolQf+3lsBLQS7F5+qqGz56osM0VT8zP0FqC4dF33ZA3uvMeSGqilb1+sa
iUZ0qyEuyWZZ6PEl4Xk54thVEuQUFYDZGA8/F7E03/V9o1DN44NiHZOlCATe/Rn1UqNUSd12Ne4+
vGkEOFqtCwDSBlXOXSMc3ti8CDr5nKLpjoRCs2aLpnV1CkVvXiyDNGxThsIYmjF/q2vHGTYX0svD
/g8nRNfmmclmdWhNty84lp+BugNXInsrfMHj5mnoFI+Aj1MsyIWQmbxa6CzVBN86UlxcFTDz0a31
c6DwC9GD21x2HLJPjM5QXKWmAiA3tJ/hl/faZxyDWgLoxHakuk0wWGVIPLDDrs8CuhzHiNQEZHXQ
UWKYrpgbPHrxlW6nCaTZflOyRqGWowCJekqSGL0//v76tExzyqFjYDE2Iax6eYfXo7LheTOTVbsx
5YsdPqMVqY1YYbbhzeHRFH2Lr/ELBlrxE1/L88XyyXGjo+Kse6Xr948rbxose26nuLsWxgFmYVvN
c24rDUaJhWU1jBpuVrPlgJ2Vt6IFcts2kXPbKjxRJQhcgTAdBJ60qajULtaW0CYjeUixgZM0ZdrM
guedsS2VZx6RlAkeNj6+8yQV+wro+EDAfrfBncfkFc9RrgWc2t8LQzssXdBwk4hxCYUFZDUA2Wk+
rZ3MoZzmhgP+vvVm3p6HdWv/+9YBQ1SgfulDZyMhrhU6Nq7HxzUJSi+Zqr4vyKrrii4J7V7j2koU
Wbfs0o8LRIKTbchJE60QXu1swnsV2iTAiLO2Ua8DNwxF1m5SWk+RjnHfqptbmoTZwXe/bzugze2O
DKQczbH3zMXUK1a/FqfCEq2nDfMBaxdzsbTAn3rATPEpf1nrdE9I53P5p89O3KgNWfza/yzVavj2
7//3u+0pYsQMIfkn3cHPZMZGLH/upKnmClbMckAOwMSZAQxo464IFY7ca6HVqMSiNKZzd75pLae/
wCAr4o2p9v3WCHUOdOWLOvRdlMxdh4OqkrBQFJNQqVSc5TxrPO/fsGetUEF51Hsy08iQVDJsrPAn
58drPaVvH4z25RSC122YDa8IIKjyLubQMbWNLqtC5IppK4osdQ7BJBw1cpHphoIKD06iXLdFPAwN
dBbCIBIDTbydk17y7j+CraBlRKqdqbeI3dx8rrVb3tIhnYbpDVNaMs6OXLwTaTxHby4EVD2Tp2AL
evLPJQvzC8tPbBjfaPdE/8q7xyuM7wguo8TRhuqZSIDEpneMVKhlFHRRHgyjyh+hY9Q68g5j1fw7
BWS/vugWpEVU6WX6I0poc5yzc/zW0F0qCqilIkrqW/JOjFTMebiHYiG6haMj452dbjhbpYmkbVL6
62BXrqZCNkFQ4DCai/cla20b+Hx9h/OwjNzcXi4TzEzSIrY+fhBHfmDOnRVhKnuYpDAprI5/eOec
M5qmYQ0HxZsuy1UsUbHfb06HiSaN+qutKK/GOvwMo/qShnyHvLoI/K2AIUQ3xi4+QCGFjvudVvkG
OO8/lPaCtDugTWfjgJFHrmXCJMdfuRUXAEaZdH3B9ZwxdFodvQ2NbNBh69b3yXoqa659OfTmJnEW
n68nzJPdH8vRJN8hGBA98aDz+ln16+XyXF/Ios7nq7I0sAHwudQTMQjBwqV+YluY7oqGOMrivuui
D8qycV5X7s+mztVkPIN6rI7d2PnzAtWJxyokrunQoSSA/hyyiAuVl6lTGxg4l6pSrtYU0DcWOqV8
UmIhu/6o9IhczeDG4gMp97h6skqs06G6dgfCOkIR/uLz99erMuRaneAA5fI9tqO+YtDFe5H4hmOB
6cXsqkDAiSlChh7it/LfUgGPfxO17esvmPy6iCu4ELf9IZsNHYd+eZ/xvDlp+PIcSLHykdzSvnbR
Kn2iL8Jrt6r7zflkMpFmKoFVV/635UOUiPOpGLuh2rS9EetJbJmF3jHOXLCG6IpIVO727SqeEMZy
Zyeb2hhWoNt58X01V5Ix2i6PGqFd2hNcVIwdH4G7UZPV0sBEyIVfzV20pKSMFvnIxC2ARokdwr6h
hXDLtnGellf3wfqnfs4NZdeltAS8MhGaW22H5Hiw+pxsnLq35c7Zqr97UyfcZSL0Nvzx+xZaw2K3
95Nm04da7xgdJ+ePm8Jk1wlKkqN/oajS5CARDFWC8el3x/MwmXGGMEsfQl2TTcXqqrvF00fllfx/
dvWCchSTej2Ll02HMSEg+KEOPMkEaDlwnv+OOcFY0dSwwuXpVYUmJhQ/f7cndPQkgavzPjDvULu1
/5SfJgLRVKkVa6vflV4CKOCLnIhcnptE7dtgql8qEd58iIG3RAPPYMscdCAQNWZgnOes46OJmNZi
t/Iu9D5iD9P+NrY69LthlsJQuWtCApYo1YaGbTW2Nb09shFZQT/uIzA3BON0wfn8e41hl5+PM9Pg
vcAn35MQdXwHhrG65e1tfKMFzPFVADLJHn+4tth45FOV1avAr0SpduKhV/9pEIS32uIIcb1t9aa2
7RgXGocHs/ZvcrWZH6u46LRaWqOw6ER7pvIu3DWEtt+VK6E8tr4baVCVREGdIrEawN6Anqjj/upO
j8JnMsrm6hxPazq+6//tWM4ofQXVvuNoyushdanUliigrLg0UeRp7hrT6/0uAdPPUaVExmXBmlIm
pje8k7KiOMk5PK/+/V9v4xq3BGx5XnY/So9TKKLGnO2R5uiRwh39wA5gJoVomnFbW4K539sT5Ilz
f18a9tb2qFItXX6a3bUXeb4Um0VGgZDhRQjLiARoAgrXvaoFdC8Jk0TyajX2zSFDx7Kw+pQ+J19O
tN4mUBkCaQKfw5RZmPIi23eF11uw6szQdTbkbsHYAM0T9uQjsVsMEFTH1xDM+nf0yERUZ5/Nson2
JwTH3CDCzoxTPfLkzVVrf0Du/Nhc+zdWBOncdpphL4FGqts/MKTp57EmykOyh9RIAMoHZlv9qs10
QemY+JqlazArfUjlE96kuNC4eYf6+0xB6FOob5HYKuLRSEVQtDc1/7cSnPGqmqWPzsjIA3VCvDWK
60qF8gb7ZbH/P1oM+Mfb9ctibQIN93Lue2d6YcpWUGuoXJdY36m5Cw07w3VweLmZxpvEk/Bfc6zB
+bRYOcWYGWQcoJhDAenicR/ZnywCibvexu7bb5nShjIdMOoCLM71ZHGThaTgKjuBU0RhNKVH0ssl
OaKtdYLIqqEVwzjSI9nAicKGgECRDkSjowJhS7YLaIHq+Cza+1e2wxIXsA49U8KL6MsGc4mn9Ku4
ZBMI/LZnKIowcZ8Wb9DtRrO69teeqn9tmCf0WbZu7exPD2kDGkGgByXQFgW5d1A7JHJUs6MphIlX
HHF3+CeEMxBchcV1ObQriSzBH2OLHd2tXJFyvXRauIWqlBVvcz4CLA2Y7e/UZIH4GSS2ge8mb+Ko
lS2nMUFLZV8xkmj0MhubWcTitulEWjC0Pc0Vt1/60xQNJ8e8+Plktsx82aOnIaXLfbMRaeuV2T6J
iQ47RI1pwrRRCY/TJxhsS06y2y2394P5fG5f8peBvH9P5Z66wVXq5EaBemgVBeWmuFSx9poQqm3T
W7+j32M8MPxcL4p+NUOvXY95mDsi441jDTqikPMUETvl9Sh/+SYRwsXufMb0T8hHHZtt0my+ozOc
YI8n26y8LCq6IL3Y+OAXlJ6vMKvRl6MneGvpXs6JFZPOVVWLLBBUIqDXsiQNgniihupxBne+PrLV
IVRDfFX7Mh1vrbKznxAYvk9ZZzo2htX4fpu+MWiM6KGPa8ZB9C2HVeSdEHXf4Fh8IbNFyfTTrQdu
d8fD1P7AYQw6mZzkY8GF3hta78pfimDCpuO8TI2+KuG1b01qjDX0THgsuYuOS19tbBAuk9e/+o8p
bnXgfcpBcTPoQOfgSPTMMqapvbX149e4YfyxwqrufJIzUm0gW1lfid6QN5g0wdEADBdm3M8Tym6C
mRbUQUv95Ub8baKTkJByCxfqieD8p4PheK3OWK6quSKXliEbVmsUWdQPYw1BMhttHShcCUwJ1Ga6
4H56Nfxv+G/VARHhu5oUj1NwwOFFvzd7Xgc2gGKBX1FgLB6Kjrqta+kHOdROIa142ZfGxcXBlAjJ
gcx34zNb6/+x6UvBxPIVdSga0GSDqIVauA5PtYMVSEDjj1w5G4D6tUYKU2GPmnbR399CGLBNrRsw
tZvzFBoZuDHCQclmsLiJRk0yd532r6ghRcp0uWG0gpK1E/sWFHfXEdnB0kkghqsgWd64xk6QEQDx
rKlXfxX83tmwka8J4MPyUCm7DhEYonHiTdUVAGpZPNNpEqUUWuFizbdjWuVu+S9xfuve9j800qOr
u503pC0HYg/zdMTBX+/dNgJnl3DNqwwz5VPmpGwfav4I8DZHB3he9wihqnhP1OjoToTcVXuHihCC
QsgKUx8xWLiYnoZDId7wkRVt6g+Sl9caOS1SXoe+LdyUP0hZGuxkQg5blCgqrIfY5/qKnXtt3Z5H
Bv5ZZcVTFQU/nWb6Q+IiACSnhRsHNXI4xMHqIXz85J4t5jdeuwwg8ZJmDVJLoMVeOZf0jKXNCSqA
hVso4PNZFMiNGamuLp6ycaL5i1o2wdmPzWdWgCxJEHwbWIUqWh99LibTf0JGAFruTBPBgsbYZqi1
d9aBrFUG8d18bKt2cgBKXOO8hh3uiYDFpJu/QlTwejjqz5dTYXQ9H3wfFLHRRgy/stouFEXh9GKt
75+IdXn0VtfwUb23P60s4ObgbXO4i8aHpPuSZs4r4rXvT+Xz2G3CzeGCvvZNxnrAfe72BFzD0Ylg
AnultMmHKEtIDL8E2BiP8AaOiQJ8kTeWnGyFqmFQjKvxATze5wcQVLDrH1w0l6fgxa8gxUTSvdYJ
GHT46BUbLtHK29uM+EJx5vImBSx/vYuDuLYHNsVjareU3IVdtlqhwbujNDoXjsmhwNKtbsRJl00T
JSDF6x7+0TVUvPU0cTax385YiymRRyZOjNJ1NlpMNbVQq1e8PAgvY4LfHGwk3kETOLSJR5nmqPSH
eX/ZAeArcA5Fe71+Uxywd+raYZmLcx1wDJurtzkoe8//hlckVIWzKIcy1mrTzaBolDTl53QBPYTU
xinfwKCnpJd7gfzxOzW+Sn72uaZ9sM8n4rmro0K4KnvkcNorG2z8xPjaS5+W5MDEEARPYDtLIDI4
6gF2R0r64ImDm6aevuNe2S2x5EBy02RmfvAgCXE4RTKHMzm00y7WXxBBVuUnEUl1xwN8iM/ug1Ir
nc/CvUQ7C1Zf2qABjh34BfMdTFYTYEMENenJdJvOvMQFMxFg15D/FLi7Rt5I+qyl3BQw6OezdAUh
KSZD7l59ezmqdN9XVhvk9veOOQ3Iy30jkhaQgURpdjXvQwI2W759JDwFv3xs4EB/oIVdYOXcAGXJ
tbok7Y9j7X50e7Hj4tuxQN4lHgGt9RaSfVIP3rkbzkT3sHad5mHycjnJ3rGaSmADWjUIPFuk6t1e
U7jbGatg8WU8e3Kp1SRp/uIOrd3AccW7Cf1lGiBSksI4q0X98DKA0MUdxqzoPJD5L7ebJkFYs5e1
lUIuPewxBzto0IG7V5+9tPs0CRfhDKaDOsCC91a0DmFpTCS2oDKEz+LPF6IZVRWOlbkE97Yw++qT
K6EMrzfs6MT1C52Wo0FPSmv4S8pPW2UglZsv40p/VgX4Rwx4UKrOqisQ/P0aJyXLLbtbKnBbJqUA
uGDrcPw1W442hBHCN1m4v8V03KAgzyMWi6TXTug9krf8iEsPjZhGI7V4Qd4uKDoqcCGwkDcAmB1H
NzMfOHctax/+5f+R92clUScu9eKxWezonynLn4XD8vE4YpE2XkAyBBP453RGJuASSoEdUgxih8zL
QUhTUNgAKDlTFxFz8domYYv2hXyvB81k1Jq77WGHtFM3L29msjafKj6t5z73GHiAFLCiGqPpWB70
4Ggo9a8WNhCLZt62X0AAHw3ezJ4fncq4gxE9aAsOHOqSrWzxUNGFQ/SynjX9/7mNS2/gFW32SszW
Cussuz61Ek+XAjUXMM65hsSOcKe9bLMfXhoRMHGDGmMb+dl/DeDxVeE1Zn+88V2krKU6QECqfD5S
WGBSagAlJSDpYsA0SLh91bxVRqkWVFAJxO95eeGBQAjBPhKir51lXAIDANL0ADOH3h6b72IeS+8S
7/JqGQsk+n2QICB6lFP43gFo1hYOjPEcEzXVQYligZApAv1nFeqxvhMwSrAhxxpQMHHfzUxFdSdF
lwMLVwMT28jKdx+ebe0rIvXxg7LvQbt0lQkOSR31Ufal3ZIA/ARGXoCVq0amqVj836ENlc3zb02D
fhw5fIZdylNOtR5J6wFS8qs/UzcbHVca1nDw2S2qMZvOEIm4GeVGG4Oo60fnFY8AIzlKPJqZJrjY
M2gymUpL81cNQHV7v6yeDOn+rVii1aIz2LPIpOn2ZE6Dlm10UAfRT7MJ2pQ+tv8HVC8Li+hCZx7l
922pCmJoFW7lOyM9R3lHane3+9icLWzb1+L8VqIXChICwyq6Z+ztUfvwGVR+vch63g23K2CrcwB+
D20E+i+3RgOl6gYKbKI0Ihs6IRvRVUSIdBtogdNCNGF5um1Ep8B9/cBomThl4Q6fSHHy8jY/lzi7
tpd+ujc6poiFbHo70YWHAPKdOPE/EGMw0Eg2AbjL9yMJ2MWfhx9P9i2XJaTPuvh1YkxD7QiV2RWB
kIERl37ALuL4LXXcMxH3AbE3s9p+oHBOCITBOeBi0QAcVO7sluCeG91dPEX7tmGEqxx8W4dCYP9u
T/UiCbMWZPRGy9uDmzMsew63xFwZMZ+e2xQkq3L10dloljYTj7ReeXxoTcDPHGiCUW3WqgL2I2wT
8ll2JPxRR0K9n0EK/S46bYHPxO633B22VTohrdiIdt9Oam03WCaLBNSdECvoGHRNQ+OTi3YwkbQl
bVIGxmVO9Sp8p8wT1OnPwEJ4V3OenPkhHWCi1w/BlILEpG50dGHef18Py6o62xEMXU+L2GPJngiZ
7KH+N2hVafsw7T55dumGn8YpcjYrcE3ye5LIAEHLubfuZZFwdrOIrR4cRoYW0/ZXKdimChaQyS8E
MnKuiMotOF8cvi+bCMtg3t5OXtMj1ZGv7LMUyJJD1xC2el2yOyfsZ7YiT8SLGEFvrpwyFjMR08te
q+JAyfMi+6L0NFjAqK9WvcdDyrOSvMDRtm/UhqifZ+DjbJBAf/uYFMa3TaIQP6jaLC06CeMv/1Zm
n9msB+s3WdXlhP6diBjwD1x0ik4C26kx+nPSILi523M2J3NkmANmsF4TPf1IF6itM/FcnOAQov4w
dl4dUbnDYYSyqQBimd+G9UmWm3NHr4GhlgxyY1meS+LV13FiIMOEQAZDrxO5jNnFMo4pF5i2v+hu
6IwenW283483We3qnjRdqqJ8BIjlhMv4eJKQkoGL+Kej9R3cSRdUvgUTLXfb3ExXycpv5hgZf4Pq
IqwQX27z9W2lFjcQjMVpGyJLgOu/Wt0r9pxDeW82sDEAK4BIEIL9YpzWnfvG7Opzr9oi+1pxRjkP
mZtPpnQFj/pUGvHDORb3t6dhXQSonb8SFSu6Oy25PDPWRn/pBlGKLhntRaQZSPrVA1QHMQmd+Imi
moYPfSRSEyUf870G0shysCIl6rj/MNsmceebHL5Eg5nJn2Y92V2QlZnUXm2taE1kiXznwb+P/LDe
8IcQ513GJtJNUA/vNSIsj+YRhdknkF6jNALvbV/IE5UGfZlffgoiG4WB1+k/umlcRdTBJWZOATCk
H/9N2iT1AAWQbcg8F1j4ynYvdYBpW7++xgSsFffZqf/wxB26QGra/YZinaR7fIq0iqJPjwdpmsVb
7sL5UBhw0ywWfvMPOJDbCaKvtb+qFZrhhrxGCLriSfpL5lQFr6FVU7/U992b22HKb8xHe6TKoTYu
Q9wpZDvRY8Ty4OPKbnbB5FaYYfqNCwCCHAMX1jcFXoN5TKYr34xo3gJeH2dDXevF3hvJZKmdWW9r
OFOiXlM5KHh/4k/D3DPT02cW7X8b1Kj4bbNh96dz3tC0WH3tYlBgdr92Mug8GfHVv6LUe65gIaYQ
o0zHOs6Ut/5ke+5mrJPowE/JYGPACMlAe4jtHQPORX/l+fRBhyMa7P5/ej+26gOiq5R1YxXR7jXM
K5KGL+ztRYNz3+FUA1mR9hfDwjge9U9/VvSjXCZvQPWRReYwb0aSipsGLmnwJWbMdv2GrVcpRbnR
gBOVUU6WCOgvROThBegaRwAhnS+Etg+hCoa/EKKjA+LEbGXj9q9z3crxT8vN/+0GrMw47CEgB8/y
MjC6uqTQ+8VsoajjamvlQi0EKC1Is/T5VlRSjdI+de+yz4oPto5gLalXigxWE4fwEdKWAp8zZ65R
FxpzvsYjiAj6cIL998TMyGXQCyMT1dmGQKt88LuZ+6M6buyMH5l84Ab6aB0Kkm9sVCEL9J/ecrwE
Viiuh8L5nLAEFj/+ysGE68JMDVHzwUk9BNlGej+atULyj59Z8wvSu6BKgH7zRPuXsYj+S7beFvKr
15apHlgVpZXV1dZATAxzoHNnl/zvvFj6dj6Iew8U2/ujY2lnhGwCQvwLt6F217kZvOHcEnY8jnqx
kf2OIrEBuNgFwCgFEzjvJd+jBL7QYa47z8BDvQZvdpuDtCCoIT0eHezlETcrbttgsBFd71nWXGrd
wqHOE9lnsDYEEcuWSTHmQEXTmYN16NP0FDdTI7h8L/lujmYqLyaQoKkNPTfZse9O7wFFnH19XT4r
tX9p7dInCU7VA7fzDoyEgbbxIixTAywg6+qHaImOpy2kGeYZKOoj6g8JathKUtNOVvuq8xNrMaLL
RLo3YrsGvv70DJAkl9658M0iVJEPpozV3+/yF+UFOKtZeOtOk1cY9c7+MxIqHYeXzvWVharM0nmL
/ePlJKbSG87oWxGTc6MYwwqvPjqY+NkpsRKF17j6rlAXOsvBwHPBlIBsBpwLSsXISfbPHLgxZ51J
F6qHcLGacEPQyvCiVWh76ZFrSEmY89q5bVnV8KnpQ8qP3+Od3sFOMR1qNNF0amsF9ToBkkmyPqYw
VHxgYP/WGje0VkBcyp0bsFdYOcpCXHyhNR058LYv2pUCLUuAb0G7p2/yppbjOrTiHqBQCT3a2VbM
zx3QELKBkFcLXxGjrm9HclskRv4Xe+xI/EPodmX7zdssKQWKi2TuwfJX0CQ63tjCFkghGwxoiCRk
a9Jmb8Zh1E3HAuDvANHPqD9Z3tSayA1bsqtJnj4A2MkYJH8HsFIhB0z3IakfJSTbADDNJqTuVJO2
jBgrVmXn9dffzRC3AzD+n2Hl+k0XaXhl2RwHkyMCrH/jM7NA1eDVBxasPyP5cQodWBVn3ak+Cgi9
z1XfcjYy6O3FJMqJWbPxPTgjwS8CUwUXMtVO97gA3EzvQRO5f/HTJvtLERiE8Feqh7oh4RGMgcQK
7BG3/tKMv2IX5qrynszDAgJMj9ISSN8xAnVrcsK+5xOuL20lhc40FjCEP8dN3F4sH1Qt5yYByryb
+tMdvHSpJjfhqaZ0IJU1Z2Fuc//UXFtWFUWEzU4PHa/FtjsAL3PVcb8XFz+VE6pVX3A7N85vNmyy
/Chc07KUadMN8lTfaktoL/ND/Cf8Hm4RXdj1xnQ3zgywxiFWWy+JO1BpKNDGesoiTHs68pJ+SuNP
Faj+WvusvUX4VobpCX/x1NnSYXZaI/NHmEGWFTk/mfG/pbz9fMx3TmR8p14mb9fX+FIy2UjN/Hod
FGQeeQERJvBQF0Zn92/j52R6pPib3+w9o5iZzpvNAsceWvSWiU/CV00qN/HxWRC3GWbmvVG1mjbB
T0SSov05mn3ORkEtUZFyezpBKi5FxnS3w8OWnLAsKSRzVqFI6tOWGy1qgN3UlAYjWVo5/YZA3kTs
X3o4mmYXpwV4JRfV4al1dbEd0LJOPENLF4mF8W2GIkxQxx9YSN35WfyE9jlP0VGlab20BiiVwn4l
iGEY7iHAA0rlP9hqJ8t50msKgjefDPLzzpErP8q4s3Xi8uc8q4AGL01y2T1/7N8JeEJEvYpLPNLy
+4wMCFnYxVYl6bXfRV2Kxu7EYn8YRgJECIlTYqUSeOPNvJcQHLrT/bYiKQjkk3iMWxOQ3fnuhMf6
xKmedEt+bcKAwhk99FrLamOIdY9TIBAGDNVEnjEFFUzAaJ/b10oIe0GmUW6IQU1Bw0+uIYQOLCxV
v7a58sTd2/iFToWJW3S0XwiXbpcn2LiggYwDUybZrf4l+UcNYRA1E/xqyB6aciVbF7phMIk/NXSm
wFCrJtdNqFyIUepeQ/5ZsJfVe0XzCkR0mOzgiTvBJDFbF9n+Do6t3oEluqoW1jD9BxxvZtHhAN5N
ct5r3HNGQCnKOUNmCwVZIj9JP09DnqaBNxsOmCZHYFYaYt3Wa+8rsh9CN7O1buEio8BOyE2H8Ast
MhJ7IjKVjsrhtSPxrgm0plWFoGx6G5Y6IUOYGdmIRJ74MlbUqtKWSljg1irCR1IQHD80PwYDsPiD
jmUHXgNoxuL9rUBwFdwjxRxyfF0WL+RzYfL6fnQXkeJIn1T9EqDAO5m7H91qHyicGTR6G1rYfUn7
sg+eNUAs9IXd47zi5vsOTBeeN3rT5VDit6Ysss47edFFO93MVd/xOeL3xCGFYk4h5Et1BnNj8GeJ
JcOAIkcUvVjapwbW7t1+SQ/gvUh9jZBLl2whRoyz5ni1gEh9R5zh0dbteo1UGfW1TGyYtGttE9Bp
npK/kt3fXpxzmAF0LJUIqelMDWZaq8+Eh9CyYBHHul5VtA8EHVprxNfj6e4MYKZxloJLlwjd/thn
CA/chhgBQPXXRXsb/sRR85WBmjgUXO6jihNb6V+T6Ae1vgDS6zaDSWV0Kkf2gDn15vrIntQXZkFj
+qhm9S2OxAYYxHyAaVICoxaoi8v6VEuYY9MnDFQBBqQwDLM+ohEdMwO83KuIRLSo0EnxABgk+ax4
myxa0FaiMzLMjc+hdj3uqxkyjkdVQhB+zZ8IJSXzFp6m09O2Qxuf0EobocsnPIKWooj1mTq/vWfe
h7CvvjI4DhGpqCXjwo89p2c33XaebwnjbmI9fw6ONfRm6CV8bHKyQTCP707X21xx1Ueu1c7+F6ns
IVAzLP92j8/1i6qu+x4jQ3JmkpC3P4ZQRFzkeJ3mDoXTFIvezYmF+CkD0PQD3rlVYO3USmyYp5o0
VLxHF59s0dohhkKz9ZxhQgOZvtb7CW7+WLdKBMIDptsd5oixUDTdyZ17BoUFwVuiZPbpNIzuHy3O
dtZZkLcdo/5mLwXUfXd7EhV8G+rcl1eHI11Y0AyW2SZbecaaKhJbu1xdqdhw1ZQdYoWLAT7deu09
xjoZAgszg4tZTZqK0zB7Ffyh+TCJoKC01+exBS8mtRKFM68wZtYS0j2R/+BRLCagnOuhlJB1Pmfu
VFgwJutJ6WueHiWXBzxA/lz1JjrKg/0qpmgYyLpJyx2t1tRJz05G8w66l8tY0jmu/saPuj5Xgs/A
1jtuXk47rVVgeg0sYykPiBZMwNyv9IPILBuze3QsaV3w7/mnmlCXS6uwMZdpGDeaf0a0zl0Qih4e
biPYJk2Y1XPNmdLQ3tgEM9M0V6dJ2+qtzEucCLcUSpw5PYjcyRb7mmgZ/9i/elgZGlssaV/SOcuy
I89zG53QOWfxvKTr51DAk4z6VKbTIMln2W8IrGZ4r+7uerccBEYdYP0Dp1hZYmK9i4ArbQ4wcW34
MrtwvUXrZGJ8DZCNYMQo9APzAdNffVpMlylx/7d+Yhoh3CxxUH8xXNgz8fzQn08EkSEXvu3pHOQm
ubxcjhoioZQtWiv24v67oWjpjrMVxsxO2B11h6Nkjh/vA55hNvYfz36Mwd3VD5Q7ThXhu5xXgK+s
vNKHIFT9PRvrJZDIz5Ka7IOhv753MCWVbD05HyRbPccZxWcHR07UvoU0NTZ2Q0X7gajcQOWxEhcI
6vhqPTOb7z2EWiHtlsyA/Feo1xlPQWTnUL1corC5XamixORM20pQDSu1aUXNcJbsShEzQSdVpArM
Kf6QOE+xIOTg1kI4L5EVoA4gAONAcrYEibpJEfwvq8iW6ETQ78ozmW+KeCbCgYAfhd/PWYvXBgLh
KY3KkpWWU86/efui3Cs84QdEVoy9gi7AZW5FPbQWsqyAMTnDjSQofTzgyPIfQ5/UfeWlEAHz2026
D1rMkHrx63eu0GXHhy2QJ9kQUDNLcA+1kqFtrXzTfizhL+f6ccMN/e0capwYE8phD1Dw99C45Udx
n/xtkS70fenGFOPf6N2kXo3sGfnVKJYkFEmFrpEohlJMycuNltDK/YY5HqG/uzR270bXGO/O2sbC
enkuGQcizKph0M20R5l5BnLwiFNVPgyKlFC/RkOGjPdEwLptxFJTWPuM4u0p+dLFa3kMOjU1571Y
9FtnJHaqaCtmb1X1dQYj1nzm4/TQ2JVpkCUqSzaeYAQepi3wDJyo5dfvTcUaFP2vn/a/0VEhWGm4
hdm87jx7vVca5OuYH1D9a4l/RPeAgayBdUdcN+DlIuuKUHv4EJ92hIWBGuQ8D8izgxNB9zmm9hr5
SktVAEpuj+nDc8cCBwtg3PvPNSGN2h2nL4BhRtIb2k+Bv/VCh3OTgezKNuNnL2q6NXBNcJZQSW08
TgICgc5iNc3x0u4ai8MHAujDv7NEMGdoaeLCIKyLtpRfndfj+FNJcKIMHpZLK6VdXEf6rhx1RE+J
TQzFC9mzf0b1LULtgpXmlTqUvLEy3Zj9CkHgD0A6Yt/NNmEQWStuy/XMnZacBFYtjDG3wumHrZau
0ydqYsCHQXmQ0wjQbTEh+FPFSZwnAtjhXbHhWXUlnNS1qp1WWqKThqD6SHUBIYqIXWJ7bMPLHBSH
AhihiVl9LUITwhhmQ0b0mkCKot9cPFAklB/1PpuhO7Hcl4qOMNLo7FhOkU0JPPlX4dYg+U1vBym2
U37YKI10I/ySFp/XL/4x1PLZ7PlR1HzFJNt+ao9Mc+rjkkkP2g/bR/Wnn4JlsLnUp5r7I+RClzhz
tYjS9zoOz4i53Ef+ZOFAVcZ8Yl/hBgKnpEfoqY9/Kzd0ooYhDCjk5z6pDCVu27kMRZ3uzK2lT2DA
GjMDV2b/wA6hzQkLTxyljUae6gXP86oIwxUCbOOW4EWkGgGaQwTKyJuQ7n2teJ5i/1pC9mRnLhKL
fmQQVNS/PNeATQQRWbZ6Qat/k9qxzquDS154ZXxhZFYfofDQBCtenHDvF8sBscYP3LH/y8L/13iF
z7z6KlfFaUmJ5KZ+Qxn9LBW0x8R/3mEvOdiVIapKn3KH3MjPTGBnBU9NgBoc86quFMAhpvBfKFqu
dvZS0QEWGL7v7j4MmYuTcA1gJMCLbQLtkjuSBZO6ML3pHoPNghdc8APLRAUHmx/vw3B2L5eIwTLZ
Svt8Yl2LKh9kEie4uvbPVaZgbhM5ghU2rJJlUU15rM1CSnZ/lqbqLZ2aWkd3KkbWX9x9MwYwnVBC
ewlPFVUCl3BWoE9i0ejgT89QlJCHS4iVXF5Iv4iyap2TUo+dlbsIGK4GC8+TxEQ3Tyow92rku5ey
KHTEpvLYTjW9gPJWGJ8xSYqCSyq4AdQ0kJpngWeaJoD2zFl/nU5m5N7p8/0Zwk4F+bEQgYT9f154
LtXz64vdtA35kJB3FrmSa38aIP8sHHV3BCLM5Uq+GjCvol++t1xw/4rUz4J7hARtBssfVi780GpQ
iemEj1Wnxdr/mickY0sdcKEgzT0nby8IUP5vZsWvacvM5wfWpakTEx2MKm0Ms1FVl8+f/shOGNG/
A8F8zZdQ/mjlxMpOflkg7KORRgtw3I5CXXgxz7ZZLlGcnKgGB0XkY/0BKWANvRwXxRrc+7Y0t/f7
fv3ca/fDwdybb5VBog+Mg4l7ZDquzI3LJu0rl1pYVC4OHafFvizAcYYr8D+/huwLW/heqGt9DEjP
aGx5v1wyId6mOBQcAdGnaJvCl5PHZkOxPsAJmA3ix9oYwrmMdOE9tn51clazFT5mwaW21KKUPJoz
0tKMhAW36I6XjpquIHRxmPgH1OgGSjBX4J0TJA2sFXCtngCB9Xw0VkErBlETF1loynjcsThBawbi
JPqkbuCN7LT/WFTX9RU6O/SwhQ7zeihXjmLFlWbdgq/EBKF3PTRDXfxYBb/0xPbNItIwuHjCnQE8
AccX10p6R70SU4w+g+jA110E0amuKnRKUMKKiZhbHuupplDS8bczTgVK8nf3ubP3/4sYhQCbv5x3
72ly5QVbF9+WersaGxdZluN0qScGYBls4rqirRM74VOV4sqi1LCmnvc6dCaVue7rvoeXG0UDvE2P
tqGpvehbHfpUt2x6BEXpiOMKUulyEKt2S2jC7Z+qRDlr740ux7yxOTg+H8L+SmAnIv3D+rX+OEs/
UtoOKzhSrxKmc1jy/aTQFP+xU2NtADglUvYWF4lPSYrkj855u7cbDF2BjGwHox8bpaZV+GBI0BeH
qB5jE/SGxBv05mGnHeuZ/ngvs3R2yQjPqHdXKBrCMgzUV9kz5hpM2y1e8w8w4/ytyoJmgEc6vXbN
m6gHxuKKtfdah/nyTSf+FxX1SoFtKm4iU88fD1q+StEJGYg4ahaGq372QUxoPzGV3lgh6YKqWplK
//Sz9dkIGSvQiO6Tg5q+nj4hK3Whv3U7zjw8uW/4VU/zmdjnx1/8wnJUU2Ls/JRbmfaox9gAwksx
SIyjaS5PAkdR1ptiYfSHGyGMuPD9M5xAF3N8mloXfEiauu0srdM5R33SjijDmn1tz9Vxtn+lbzek
ma4lTlSKaFRWNSHyRcV8TSVMH3RSySUvGLgEgH4HaMkUbyva6YToDgajN89V9QCIo0e+7KIW5Qrm
gw/Y52zV6tlWSGERv3fS9Uyzp6wASFOS5zkdD2hMD1s5Ou0N2Q+1HkvF8O93F2iEr1MkFWnCQZMM
0bB3tcLyNnNTVzmFNft8+290prAGSprLayqGMuL0gdvtSwGpwgTbGpxmzzCx29Bg5vd5sHMPNOnD
jmLT0D64xkEOkvZPn6luQ9h8snsrC+oqaRoYEK3Te1NkHOA6ocoBoIaYIOtZ/vJIku50ohfQmxWp
3DeRD4sqUjr0G74bYPwG3Cf2Wdla4CoEFR/JOlUgmDADoLznU3hyPU5cdAaoy9FkgNwIZgj28qNU
sCnQoPRcTDg6Gbpn+HpgeL2jWSFLnbESEogYzAF0EgG0B6nhVQQC0+ngNZjOFRHZb8GNDfGSfv4R
bfl8bzh6Z5UZgokmCCWBhrOMtE5aJsFQBh/18w7ignFqmd1lhevIJZpyBa/YHMM0dpO5bILKxqIf
rTdvcqhXiErCSWaGpHT8C25Y5VeK97qkk93nWVlUvbgq7zQc8mwMJgfFasNuVsid/Qbtijwv059v
lzmPQG6hSPKDNEi0C8+uLJ/p2/upbIO7KfOQ+IBKZOhhYkU/zLyoLYLfVj37uQYBAOEpAUuYrOAw
TPv6iVcKSbiX/vZtxJJCCddSdPKOBjLUC6su8PEVRXxZs2GVOHs8zagfcKOfHTFZklax3Zpzqr4k
0rx5hh9/w92eYwufvvLXzTwAiRP1ekEGiK8D4OBJfK0s1laUGThvMYv6qFJaHJn0UEaayUpZJxvO
wDzUEncuIk1BbvCx8sIFsIaMa72veLA60WWkL3mYjGqcXtaQEeCDVerbbkV1HaYD/k2VYCgq3T95
753gFcpfDED8mKBWamUZnpG6FKIp44bGmEkoNKeJJPt+LMkaiSG+z9z8fMh8LJifjCkDoZYPK4eL
tYJHf0SBhHkW1IQVaz0mtH86O/LWVlXSN4m8cOxhn/V+fou4C2ldTX36wQ9BE8HiI2+atEHoQpeH
BTTD20OoWKBtZEihDlxB49ngR8/1BVPN3JtdKimlOlMJwzH8IWXnM2e2r2yfMd0PDCE1iqeQd9B1
RgjOkq3AqztgwfvVVjl4/X4Wx+QQgnKipqVbQ/EoTG2ShOrYiRpAo6ibiGachySAS0WvYkF7mC49
N/lP5uGqBRCv+LiwCoerAI39TkMuYmTCWBGImqX8xkAG6SruyrenBC8UFLC/h9VrcVb5tOKXQm7i
2DkAGeu+fSNX28puMQHTsSnzmSjq5pVQMaxAnStzrFygqcYQWNyT4ARst03Nhz9Ea2g5dNvXq0/u
AS/JKHJ5dFXzvhZLdN4OVlIJYc0fUffywZuWMD0saKMR/lnvcZT6o00tliURZptKcB33QFkcRGi1
uV/n4NEX6AN2eogjgpbp3xxP5VnpkCT4sQfRtXlFSsQ5qy5jeivAZyR0g1kPwkxbew3h0pnSGLq1
ONmSoYVCLWkW9my4NMbu7ciUTXUnNJaPEErZg5jYWGkvs+UFf7QiiTaNxi/01yXSD8EA1/ZBGq3H
YJyWgcJur1XWx1ddET2fOt2+sziAHCsiNEo9TAac0bHRstMI2USYEC+/x5Wlw+r/J4wBy7YvqLwc
bA1Gso8hZTfmDliPmjvfGdzo+1Rdcnp73wlgZY+NCHHmXFrFgtXYlHTdzTappDJ03cZHk5gONes5
c4flgGs+0PGu6CX7cudJMjf6XL/7iNg2mnECrPTaWmQfsfEe+AyRyL0dWQUi0ABEwaRmSuZsxTL/
mlCTABh/54IXOkKp1MhjJHxkZytBDy6LNcagi1MG4muXjuNpYLHS/KzkqEQT8yqGrj0DjSIeZMqa
sBeV+ndj5ltnAoMazsBRkwkkwP//ZjoFqPJUR8fGE/6MV/waAgyXXMe9bINmsTkD0Q3NkkKFNEVf
MSDbUW/iG9kizt2PSs4y7oRHp2IipfVrLc2AAb8Fy3Jp9UbFwhEnmH7srKAo4oh607WIiZzRittf
6Y7RYJ66SKVr0llUSryTkVwWvfPW4vdd8Br0LUifLQmjMnCNal5u6hIyUSrQHeRMTDKaL824HgYL
pZ+MT2FvhtPYIjAl41oBRSsVDBRf1bLsD1cRIYMFJlcQu69XtB/4CQMoyfuT6QooGtqoSD8bFtHS
tVlRg2YjpUqkO4Eny8o0x1TWMs6rA6htwMyBa6frx/5q1hCAgTwwsnJX7gcrSQSy33eB4jX6EYhb
SSCPLTfJ/yotjlcnjZUAbntF6biIffIkyVj5G0YLb3ovzqP+SxS+hCei6QpeLLav6gALp0xAYdiO
2JtVjf+XDKck9iArqIYw43HDKvpSiRm+xcae31xXxbkKetS9bDg5iR6uKvsoRr7j4f3IDRS6WVvN
juB9BIpXu7cBrJsziuPANh5h3ZFIY+LvSdiMmYU7Kkcj6P2cl2awuZSKf7Xc5nGMNDYOjxqoQ42I
HbXNdmz2HqH2cYvT7/lT2XvNkIJq5c4uGrVerpus1VcEoG+xAhzXyO3n5L7Q5JAZvN+4f4p9BrVw
YOW9Qo43fbezNXEPtYR8h0jJhknunKQAhisFJZaVvd4WhdowB3xbTwmsU7Za5ygKMHXRY+mq4abb
spz/IBRywFG/RkktBjm0fL/Fu+Yu5+1+larw92LM2ylofiW2EuHEpXrXiPXqrldPR8ThBvTHN8PN
GgAphfkvjGPEjWCf/ebCjORQuK2mgbKbLNYWOiEavSKuGLezDYq8oLswpjULv8jH7B33XTZBVzws
FFrROzYCavmm5+LE5MFUgMOaZyLB3/+31XVoab9aydbikSaCkQPktASe/33EFmNKnB4C7aOBGfo7
KaBzklVrv6K1KvA524XFdE93ifoVByY6EL9yCTvGJPikm8iZYeh69muuHYBIjdtVyrunW3V9IXIs
Vjd9f3zSsJ8+3pRvO91rXozPpnnO0KvG7PgzXNmiyykzpFPv0m+ZNLTTE2Tb9cIqqv1Oj3PJ8UVQ
1Sf4FfSea3nto7GVDFNUYXF5eNCOLtRsGnBVzi/wJiDb5DvS8kP6TstXrkbZucwbsWSVcrKtv32+
w6NiB3MldgE3OxOVSWLyZXvCbcpZRpnpu8AWJWzZVpZvxYNaB+yWlor3ZFLoUGu7DmOji2Q+cjsx
QH9WPJGO1qKbp7n7im3/2pgfAY1zlpZ8pMxPNZg79bs/ybs4WoBBJAK8W2WVZLK+5Ifwj1dFTQRc
hLMNVlmxbTo1CqIOKZ1Eg9ZYZ2u2vAff5sYMwcMS41xsZ3uDVekITYZu3KZxcTIVj/MY1YCVi8hp
qYVyqsCIzWINQkGzwGpGxgQGLXA5OTluXPMmXMVU0mt1qnGm7Un+U7nn3jf1v7llUpYEj0+7W22i
f6zFCedYueSlCVXxGr5aENNNHe2vLCd+3zR44ObYsR5EDGDOOZNvZWLnF1OpV3v5VEy3Uj2VPTwN
nkTdqWZbTqjgz5fI5+egWwr0ortlVSJeJTMmR/XdqG2fSeza6PjRBvsgMW2ZwENRVMxZxIhm7ARI
0O8A1L47Mdpoub4EbcxXilHW3/+/ieTXdVFE9hFZCjq9Q6rkjEMcUqC/txeRqeCSF8fowu1c87xM
ms0a425bRO974Y0Af/VhaVqSYAikmmhQ7quMtmMo6gwdDUX1LxcPJklSE73XGGSqwNaX0RTtpvuq
LDii0OiDEl04ekRevevMQgAzLpeJ1nZbfLxwCHG1tIa5kjyUmzSKxeNHhPg6jezI+Y0DJOIgzrZs
udRqm+TwldSZ5r0isjbQUun77D7sGYEe+TJgPIfxd53OoihPqwkHjCqlD3QwIs0r8kr9xn+AYXEs
t/RFImt1H0MmLs3AC5B/m0GVMXHVt4QzObkKGRFj1HKLXYYUAKTdvExuGyZL30QavDumdx0sKJJG
bhNuEadY+KRv3wCO+2dexxJkj09/pIMuIpOoTBm8EfiWzaUdLLH4A0vZunoxjivP0Rd9LVEzLpjR
TO9pdKQkXZs+E0ZZ6W9gLXOfZ/QhB5rh5ARtiYReuhUWxI8MCxR90YOJkFU+3je843UXx/XCVaJt
ULiTc4YsMjOpJuat1FumCrnBE2KPdhOWxOlr2PpmMqxsKq43bb88kKiaUXVp8enlb7r1nmzamoyU
27ZxAXho3EgHi468jI3T2JNQKB1DHN/YW8AXy+ruwy6DZt5gcBmuQ0mScMuVQ8rPiIrJPAXkvegb
KE+HSvtEvhQjokylhHszPvMBqdhMibe1FQDLTulQfWXeRLXKyJtYLyiO5rPhyB2yN5XIeCbYiRw9
fsAji5WP32q8QLSNo5Xr1m5Z6Ia77dJzMt1D+J+m6mEpp4+Sph+QywoQgfQW6e3AqBrsffl3fD++
dSixOBtlvEXSd/VQMzVgviTxlQp8N1bNf3O/2asmUBfgknVA38U6QCIbVgHb8qJsgzooALIyIqN3
nQoY52Tz+qnQyL7v+XAn61/kYI8lLpCcxezjlm8glVgspH34EI/lut8KAyKYdkFZZzJp+HDGgp9/
VlbPxw8qs42gtwXaz+fQGSgd7O29IAdt+HILcWkaWiI2eVvwx8vIPmkYFiR5bmWum6HXJ4upRCYA
ZtuQ77yljkCVDa3MSPvtp/Jcg8i65g4MC8CYHeO4y50dNTqnqHQrY4DvnVxXFbjCGCIqxul2FMTf
QAN+QLy/nFdgQcvXrt+FTJbnMdFBjzoZ39W7w3DEGR2ohQOsHzcZMVEGOHVFGk8rP3sbNJt0vfxX
ouvkPQS5xxK+Hi7UFkHBaspaQMED5J3cJHQ/DietIUq+jam/vHvyPMYaig4qWJAfIygKcZzhu188
gBBEgpncaZoz4u6XOARNEheDN6ViHhPeFkh3cjH8MR0Q5/1PC0J+TWxpKMHyNsYn0nw4CtIxErIz
/yvmpjvBEmbEzutTINn+/4fda5pFw7bZOlAwsDj3u1z7TKe0j/um8gf1nsYuc6O9wC1VC9UPkWsl
8xCqSsuxDgi7dPlRj7Jeul1ZhXRmwSEIGOyOTnP3qwbIZdQlonbhD9SG4Fad4jfSYk53JoQoWvn6
V12O2TTEJjIH3+dF/fohsj+LeSL6jL6zYe/K8g1HqO8E0DHLcUqp5Qim4VIigpZK5UiN2XlbrK9+
ca4gFx/UR628moOPz9Pa6G6PQjUW56wOCX/Q6mQcWTOPikdw/k+IFR9QOhPDEepC5RiF19vFYJY2
g72ziHMsLkQpikINY6vKzKr6Owv/YSIf9/0bVZ9QkKZFmUOOZB9S675v33rkknZU6+BOmy86oZUG
Jjlxn9W/FQWDM22b7+HuEEjDdGTq8cNdpq4Jujj3Xm6k483lVMDzaPG+SDz4WbSTTJN9chxuLups
cFdgv6w6lyZEjPiengbX1doJynZbr+q+kTDp7HgDwmJ7J7UOKrGqk3XpSSswTS8cXsp+GecREby1
2jBiXY+JpKLLQS7CadEL+rr4s2DgDGZhKT+w5uI7Nrs5HX+3/GepPlx/X3ItKU3hG+8wsFcBMV25
d4pZNnPRy6wdnPaCeWyPyDbHSDou1F24/Y5F76EhA5ChFPdoA49MyNy97fIsAm8CFZmfjenvRfvE
IGoZ/VVUzy3XVm7JlZBmjDn6s/1O6t58zUmBuiQdIIkDJfvehhVneawxA57VsYxY2sfl6omIP9PH
QUX8zPAplTQUXAqaBrcT9MK9wOCOGe6iZWAIC5tiIzdSknXYL3cbFyHjadFoN3SPqvWvuCFYIFnu
Hwjp2iyevgYEh+QELR82VUpIkOznjukwSEyxtWxecxH+rdBcM3HdwKO4cmKXASXHHMTY18yNN5qR
7Ghb6ybVnA+gvF8ZDzFCa/J0uVApw+e7+zwNWeUpHmjz+fVjjXuWx3+4O27Ews5CjbeZW2plHguE
gsA7ojhNvW1ijlYWpqf03vpj2wL1tJgLmvDlv+s+CI3XfBZz6VQJ5gk5MWncbx+RP2uFDUwfCCeN
gN9GzJ/cE3FRs+2ep/Ml8KlyPL+u1Q/Cb6GoHbDf7Ihd4lS88eA4OuqUdrSnofUDVvGROi3BcYfg
EXgNaXx2LWaPtZdR4PLE2eujqSTSnG19PaMX9g+INcqEc5a+aUSdjlhWc65iMNToqB4eym17PJZ8
GvK6fnvaqBItd5eCqcXq7f8AaBYxeO0sajbMr4TlUZBQTrfYmlNUhE/9e/R49H5tOhY1y8fGreIS
sdglm/zlJmKZCO6E0bm1704kbe3fnAYSE2Rs6yn5SeeAPUj9UiHbvZKvkeE5u1wPMR47CDpOrzaq
MIM+2M3FLTHj8R//Et86U+um150FAFgnD7oRWaLw+ioFCUMcLailnWanLm7x6+bGsMGQhp/ou1/W
q5+B8EAZvJVmXA+IPLI3pggAjK+7eeV7/EIL+HL+2Cy8roxjf0DdVHZ3+F3xZqNF8TFakzJaQPOL
YSFgSuhhjb2Lip0rXVFd1DGBjod1vT4bR1i/SxmOgtTFpuyOY6M1JHwQiJq8YUOMHog9VtnWMQ/O
HM6YS4/sJy5S0KGlU5HPauYYekJnMLyLyLYL3RhsY9+v+REPwLfq9mDe+sldWcFFEwk4y4L0YZlU
7QTntE4fC+CcfQZ0Ot2xSROIZak/BTZoNisPK/AzkxjSERY+WKUsLQjOmvD/aRfiZUoD/ozSAOS9
QmWRa4yYdyROPg2JNdn63BKq+DF9OJreNs7QOqVtpygH5chgxY1p2hHi1M8K+03ZO4GL6cHQXuMW
EiilIReKLXiOoakPSz35w7DQmu3S+srunRfJ+oGdv0qwjNid46hdVizas754i+vBIsc1m295ADvo
r6otJKs8VI5nQcdN9MXXZlGfisSjRb/SUahtrISol6hJoCsKBsJgHN78OaC8R578dzAiKLh8HHTa
fEaQBIVjrnBl/BBRW+nG/5MkcGgBOM7/BqWN3ohvkQcGeLcwnVNq/Y00Cv9Pxz1sSVD4oU1Yyqyp
yxqMYixU/OH2QH9vDZBuBUJtr3YLAeZ5MWFzqDVdgADgbBUwCTIhMR28jMyvkJQO/I85l8MEUlbC
GVycUvHjfSr3lUUT6M9aUOGRCjA8k9YKFpdpjLexvkiyThy31c46sNsXBWVaRboeanLAoT2TqvPr
ykEWx1m+4198iXABF19hvustYlMKt2KqTtYGb63BNtIO9iEnRuf/e4AQpG9rAqGn2hcI98FJHnmf
T9FvTK4Ge6q+qo9AuUrTKBSo0SFQEK4yF1pPKdkVadfywi3V4CpM/U86JBqVDTNFN/zU568WTWfE
HhTqFOAa9w0zYTvbb98yMqqCYSVeUC5Iu4EdpxV9MlrnqqiInebj2uKO7IBgny2OVi+OI/0ghoBI
CjMpHiMBBy0PSDLc0CU44rWIB0NRpiHJgjboE+h9helLE8MFdSCI5LhS1JWh3EmzCIoa7O2puadT
Cz1rlEO0xzL2EOBwUB50VKwO1xdGpAC6FJrHH2dpBZh9b2xw+JCvoKhKGpdA/U9GaD5K67d75nzO
s4do6PFIMwacZxEZ0Jklbd0WUxQ6b5jUBSVwhzYjb8AJgIPY0UcaSA6S042H+5YNSIcArtTfdmaz
6s+F5OotAlkuCAMiFhQ0FBtsQjZaEELPpi6bVUuea0f7/iZ6wasRJotYTSY8wvBZhc6AZgmvWv3X
kpur+xVWRwwLNVOU9Fl5Oq5CUdaK8y2W2llXx+anapqt7kXpflu09Af74mnE0U2xChnzXx+jlaCH
yjyDXdHVRpN4DQm1tyC0tkSgdvvnS3GxLwhxE1CZ4vH/1PSLWdx3IV4BILJ1P8x1IFeVYRi+EqV1
gcpy/XsAB4WSn/Alws79Lvh+y+ytVqK0VsmDYkgWQUsF0uc23gP1RIWeSJeI8gHLs65EbyYCx448
M4IrTxE0xcP9Zsg6iPANgM9UapL2PwablJ8UtpmelGxfODLxeFuXU5L0/9T/tAB2bTwDx2+pIGEd
92C+J7pFLaif5N6o4ylNmNkz4NNI+E5CHWviGPPuLbzx/G31ArT9vu6Objs1cBE8ShFytLxXqfxQ
EoXegQrDgSqqrQL//qACfwxCEBRMYrSTtRAll9zCmLlgK/OAXiy5kc5DMARHDnFE5iLkLdGJXhy9
4ZilIOFPc9QIhwnqey7AsMU7HLJtbs4qM6nCiJN5Mf6zkKhMjgWGYWraBxZzVlN+pBvhh+3T/HIN
p0T9eOC3I5jk+F/ruB7bIYYZU1T4MjzUOXPp/a6lEdABe0nd2GtjqOnqdzHllv+zlh1QEngU46fJ
/Ryr77naAwBUXEe4LvnD3/34pQLHKDV0dhE3OEEqJ2EkMhIEQt3ys18z3wxjm/CuyUy2EAvssuOi
7sphuKJKA35an+GltuF1E4AShj7bdzLuTxNaYHWPEJ62KZTrAmxWZLd/YkJK0ehicZBBwbiJrO3y
3wCHFxAe1J/LY4eWC106yiGGLVtRKNHhxkKq23yi3A2VLTImEBtg4ntLCf6VVm72swVJgitV+CME
nfn6anfVRCQFA96kQo7qD8QLob3CMzt7GC571oOhtxXDbYzZVka9dbf5dEolo2mC+3Qli3t0pJn8
CxW3Xncc2X82T73kVLLdXfoK5bAXrSlOGPncBXa5M9in7rcarKhPokweOmd1zCffJLm0kccpE7c0
AGQn1KOe+Jf4g45jXS1LBXV+EmcE4CCv2dong/cxz7syf9h+5zndJAA8B0Pccbcifbxpkk+pLsFW
anCKzyxxpehwECCS3U9Yg8/hbXY2MJDcRMF/oLX4r7x/yu7DyOzjXWbHjQN24G8uFTDIyfPwoEln
3lZKs1+mwPqhZ2lENRNaIXo5ZRr7FYGA6W4bHVrIL3+8qxUmlvHdndZp+e/TVBBB1gqwLC4o8ZvD
+EWsWE8Y+oflcb6p810erdfA5vAYBUU980md5p7iIZuwFCwApMOx3u1D9Tde/T0veU8EFZYCJI3m
SJqMLxKc8ozuAoWVmXUg1PssjMuTqaS2rNOMv4ao1lZkWcu11KHxO71s5DWzlt6CYJF9FpFCgnrS
20fGBBBZtwQvjasQtUslVxzFHFi/okwr4/kmmDMWZvtsPKxgQU5BiUiFbkxT1mBXnlbj2kGS0/z8
i0MmaoDkCxNqNK3xDKPNYoRKy/mpdpMUn4VMqHnW8UOdiKFckwWeQitV83Qs3cYHK0YskDi2Linq
aIsF33BAKGsmx7gsLEGhrVjw3ygUateqsNJTTLDC4eOdYv1X6defXnb3qII48rFv8HE/M1QY4F9V
rwAwzSg/tw238C7fGZshx1D8vcKECR6RCI1ebWwHg5Mgs4UH/1fKfrtP1QzSy0C+a2z6dJs7JrOt
T/4Ih59Wqhd2jJU7MyxT7gzjT0qpOy2JC2FKmydlEKscTy9BaU+QxsIfG7Tmo6o3S76VRy+hIY6a
VNAzKpJwxEVkZYhzSdHDaHULQkGbBgGkc0/jVZzJmqaAtrjuySrdtxIjOkVkp/I9a+96cs75BHB6
CUYsrovgPpR+7Y6+926QhudfQRHSlXeZzb2Hycso2dDODIckkVMBojtVcy3kM5L50hvChQrMvK0r
O1jeZrxinIKsQ/mm2lhLk/Uy6D1xbSoov2Gu0tIGbHGs+A+DLHn3ePp+DwnPme30HsDV6gpbLsni
Yy4S7B2F9drNEi1TzHpvPL188YazfCvPl/Yb4lOM4PvlXmwoioz+mC3Qg4gbwtYDjqyMFg6g/c4a
bDnu5rjBg0qOtcqu/m2EyfbxWlK/8ThlOoZ3ZpKCxH04YU7jQ9mQFdVIbKVqKSMK+MJ8/E+mJ0AD
fc7Xpr0V+k6LSk3/1HByGcfh0bP5HLs4MS4aa2o/L/9Y7IhqrYGcjcuwhIpHdn0yMLRkvGUvTBOD
BGGu4U504RPBfZ5vnamlaMLzfxFYf1r5JBgTb4APZ69QaAvcoN8kYiYDUGaLwRQ770HsxszRS7wR
XZTCupgmaIHItQ8u11e8Aws2vcT7M5Tx2AwTdntlUdZ8L7OJxmj/0gRp9Rh6MzpDW64TMrZyLJRA
SIQT9cbfZTWc4WhwJOl2JjILd8zjX4NMUTibDLmYyRVQbw8+7hUTcwHeMCyV3KDu7yx8A3mcmdCl
S5GQu84l237lgqSot8rVLoJWUgyy9rgW69f+dhiaSovD0yrlcYhp4utFyYeq6bsDrCvKZu2jihiM
3EidooNznvhI5RXKUvr6VEQYPKa42JfBcI8ugVErDSIOUDdPxNkG2A2suFas94O5vs8778OMaQfZ
HG+IkJwar0hhKJ9eHhqBeov6oz37MS31SaWhRdqLE8Fs0uJXnx5tBM14Ooq8XThUdihlE3hUHUHK
JZQHIKGyszol3nNPDSPxPdNAP2VI0pk1oxIRu0RwZJ0v7J6IZjC0EPTVv+8npk9BRhXpnSv0o/pk
JR8h3Ms3jrUNprO2cos1yFtgPSK8UFL7xTV/Rt++hhtVl9EzDgxj3qmZmfLgyK5uz4jWl6JEnQLU
XmwZPmeb8mM5JsyrtDVgnF2ihLBF/7F1ZvKWeZm8qJh7KNK0aX7C/y1LYOoUzxGJdk9tyfXCwEis
bZGokg85YVktAxHjXmuy6lIQPFGDVnfWxq3PNBdRBgAW6HlQMWnPwl8x/277dEwvmm0hiBN/vpAd
gDtA3dbZcDU1uz6pXWtO8mevzYr21wyshPUX1gTlvcHSiLzz47SjijA/nHFI/3EJt0lLbuzpNIgL
rOPVh7ydrNqDjx/jsp6AzLHgU45u/0VY5kk5q53cjs/K9liMfl4241gwtr3NzrXE+vvaR5LEOO1F
CIdNZ1wx3ukEkANPa03esOWUKtTGZChdxxjYeoxYAkrH0iovJ0ar04cCRQ7dNuKKmj5hIuCCwwm8
vgMo7aRk+G4R2knnyPiAFQz4wczR4x3I8eG+rzDuv/1bLA47magmnRx1VEU2qz0X0CsIBB1d0fXW
778U4it+AMUxrtNNUEHjKeQoWQGLD73SS49oiqRvb3cQxO2eypPFSktJUBc5Bp4jlboONfVVqoCu
3p0ibkD7k5vyolhGgJTGrZ2yt+PGlj6MshMpP76fthcz0++9rZA02Rm+a6grqRpMK6NLNfs5YV8B
EoZG8trQ47C6xULzoDRT56yL+qVe5aFs2atguSQwfGAiUqlw9eybiwZG8qi4D9wgIgHah8wKWs+Q
dB4DVOEO+gSlEDAFoXZY7LiqtBuZ8H9JEvNiKu/BIhEaYwJP43KLuOrTCXOwVj8z36rDJ9E9Kvlw
wgamSQ5DkR+AE5LQH3/8CT6kNJad6beVIiuugSXMi3RNES8TZQ3NsfnCW8jlcg237DaUcYPz8ZUR
bxMKGHKsajLBbMFVRvDyfrO0CG2KC9CSkK0XlrhlLfBgzeUWwg8cSEu6yemMmJc+3Sec6AucJQc1
M7TpQRnDLthuNyNZTYl1KImjEMFVsWGtxOwkY9hA0DAXwQzRdXzaGP6lhQaEuXoeOwkbB+qDJFo1
j9nxLQHGZCTS0j28cW25/KoO15qzXbe5eSSYXrCQNBqptbvAENfS//PORNN26wMKcv4OOdQnMSzX
rBGKIezM8PkkaNn1YJ2b65FqDKmedUYbVsO++6jK7CF0A5pY3COSOXbd/ve0EdwmD8lF7AIrxSZn
CZy4pRBeEe/gESSje8D0TGj+6nDvNor1YIJXuoArg0x/IyM2yGnOU9tMfVB/rKlAs71nq7wiEHzD
VFvCa5uweXovDzSd1ublQLpPwT9KJ2F3DjNU/vQRdKUpnC/SYnljAeSDIVqsVm08xaeK4Uu2mATE
rYo6WMIKQkQ2wMmH3KkopW3cGqT2VuitekWLTbonZvtwbLtc3gXCB6QMM2SgSP0khlPbMzxsdzs4
vvHZ8Km4J3Blqyr4y//bOjAnAfhFgirk2QTF4SYn1GAfdiKx410Plocd8gjGLi1uGQpITzCbRbHi
4TyH0HddkXeIXruzDmXd7zs1ixGVBSoVnBKomHoH7YtP/lWt5RKyj2vkPxIs7iN1TySYs/GCg8Af
JeH0kWcOjHMQwhn1vHJIn2gKY6UueahfzPM5DDh9ZL+tr9gIEtOuC2oWB7MTahV96k3jHdO8tIRG
/rdLmlF/5DoN1tYNTSGDUG+xwG+KkTTuo/0TB09AgO8sEweTO7P151u+cLEG3zeUK3ThhhxcjUdk
+DiEdPIECsTJSbf+XeFT+wAHUnRnrS4OX4le+xYbqYv+ObzIIvVguJB/Q7r6M2zSKrMbmV/4E+EU
WRdSqv/TteKYV7CQztg9xFXzb4o/1kPhwdVLM4vRtiTqxuM4xyxS9IcQ0loJSVU0vpMopwteiXLB
HytSmgfvVnsTUYg6bXZ2BA+rnh6moRg2c21Xhk0ffwqaRKoWVFSsQAP5WzAw7vLC+3W0xPqYerww
ssvpASsyLN5FQAV6S3QQap4QvzOz+IzWIMTdgFikZKdWmOwHrFkHm8Sc76FiJJfuS72/VLGenBzV
iE1ZWb2FS5KqYunPoMhtQ3Z+1CarD+ORB2R4zM/+/UpoEUk0iMYjPAonTPDtAiXuHmm9cBTQfh3Q
TFqyP5aKgK7+lhsfXiKuoFinMqsqxLmf+t92mne82vuSM+Uxk9rYT/BHUJrGky7ZULnvgNRuyiJx
YOt1cm/A0C7O3JiYZhHKvXlsxTLZaObJKYXve/IqYYTxehiClIGziN4MtweNUWRnwCpaNxIHT0TN
N5sg33dJlhp1ahrsAxfTzGuJGTRITsydZkeweWVk6S50X7zqEateVqsIAu2za9XOLlqLFPyZgpAp
FSD5v6cAW/nlNp5W/BQ4vBvmo6f7irQf6VgCWag4wToAAVrYNvyJBGcivpKJpcmwObLh9XH3u0ip
9WIsboq5HaQAUGUV1vaixYQu7Z6h8yDRUhBB6p4Er4w2WjMWPMklR0dZ1jS3pxXQdcV8bEomkPMy
ykOag42BYGECKfgWPXDIAasMgHQvG8Ehve4Mvkb2raJrZCtuI935GzzykH95/oG4UNAsGI0Qe0MD
CIf7rbm04luVn0FHOC/n/rjP48evrW8YoNZDRbKwHlsr0oLdd6/HhC6tKaUmhij75AysUVm7jROn
OoFJQqL5fb92FZMSg5fYBovBzYMMRQOFJsIKkxeV6RQ17lBtMlwCMOyvinoxA2zYKMcMoCOYO91X
kI1PCFk5+TYPtMl0sdKJCXMwg/+BNC3GjJIi3QIAv2PBj51zbqFxRd+O/O/JyKU+YcSYXod7wQZ5
XmO2cOUNdyJXMSvu1yc3CtFvdNXW8eHaWhiGgOecmzpYKy/NWYriVswN+WLDLBM/HjUENu5LxJkR
sT7EPvzD4IB+bSxpwpRmC1bWJGFFVNeY7G0zbHgSP/IpXqjUh9W90O45GlAQUfYJmwI2c6wbPza6
LR25MWdsTWjob7LR3pKOIVEyAtHJmvMotv0QQbdui05PWAM+hMSGgtW4b9ZkuwVRMl1+YyCX+Ej3
DRzSBQahMXbJxUUmrFN8p9BTKB1+4pVUzDBQZqefU5VxejdebmXydihFavurrkP3jhmhpSLUofLg
yNrn1YeEgofE0SvrycROOrZPC8oYrf8yz884NehM+mbk/7SfIMDppT+fjgXuNUHpnXtjNzxPSB/a
BDJxvX7Fv8T9fK4ubKW2ugjdHhWFX0PSXsMRVACbFO1ugEyqcjbqq8dXj2yHjw00mhfbc2QcupK4
qLZkPmC6wvkOrwj1putGwDONpztmVO5oIIubt6zrEpAGR2J4RG9brEP39jqvcDgRdOKDAYgR1MQ1
ShXo5XAJNEd/IjPywSSTPFNs61wMDQgJ9GXmVLQOjoiO76ISgDvjEPBfBlIo/xrqionCjakcSkB+
siNlUrIu+vY6VsARU6jN+9R2P5/9Z1jk9+1nLDLAyrGzaZq+eOhf/VolxFwVyxjwib8YomB1gavm
oKAe1UY6g3HnQh35PyA0mT7Hp5eULo0h4myABhAdILWLGRA3j1ssMfcy/TJX4iQ0GCQqTmLlEDka
ixPbYrhZVhEdmQVskBPo+4VuAGAzO8ehYe8x/bcXX09A514zFrlHwoCJY0/PMuP28IQl1kOeD+Ra
GaxU4SzyT1HhjVtt6MnH5ba8BgKS7SjIUWi6cZN5h30+9nxe4eoc7t0h9YHzKq47fX8wxiNsnqkh
Ooo31+mU/GqdxOsei0N7nioxJfeXoPR7a04l/+zWrQyZLc5DG//3Bi6bqTZtNkHEg33XEaql+pcY
AHupQ8eBGfb8JAkUtZVtgOipxYB9B8N3P2AZsq2rVOfxE8N4ox6iPdE9Ld1krkUDCapg7z8tGxzr
dTx+pBJ8pmM7E+J+DDOg5JCqNtLoAn6tma8TLUs4cZbwvxtnvigp/9g4Qo0lOwouYimOVFzNNlk0
Ae8wIo8pMr5mZ0YWkgY1QK04nRJyJMMPHruJR3OpgYrKUHt0n1RTt6iXj8N1zfgSzok0alKzqFMp
XwExZzD6hQZ3luCMP0kBdXKCx5q97z6hngYT9GPQkXEe7z28UuazeHnIrhKiektPUrSn9qJ8DQfa
LlPLa21UPSbNL+FfBtWXKzyvjEvDDcxIfmgCSULu1JffoJ0sI3GaLrxTh3M+x0Z/3VBMO5LTKxF7
pb/icVhQSEEnYsFT6LRamcOfQdL7Q/qlNiai0D6/lTgITsXmDkWalYBQ9N3npgk53mrHPFtovbEP
hig/kRCcQhG3xEMWeB3sszLwbJqafWzU9u1Uq4tJCVbAUV+jMdtW8O+K0RW3d0gODRvv0h/QOO8u
+EQrzwDb0XV5yIB100glbDz5y8Mg+p9BYQh3y9F5YcQ0CdVgI7TUna8HLhCbnJZwVApJP5zyxCNE
iN+k3Q8EpFP5GK50WrswDbnxVQhCOxOq9iRE3wWHCi7YLzLET+Gg0yX8glVdtjHijbVRqTI6YZoe
nQjLc7nsgPf175yNYzeT8gfP8YB1sWKxFiwSE5tla0LBXlYRfKuTWyTk5Y81vAcD3bfygbDjfo2F
8KLfcK8X2DjFT0lbkFENbZ9bdlKxFPjjWjGrDbqSvnv/4rFW33NHx15m89y7eP7UGNFyq8UZVH+I
Hn5SaEC8dve5OZIMqD/2Mk8WBuiqBhGCyVTC3WYCRnHqWqQZQoGun8G8Xd4QmB8om7h1TB56RksG
vtN8RAOXjLYHNGJ20vGl1F+krqW4pfDLV1xp9YtF9RcGrHUW7Np/Cio6V+VAMCQehnfvl0OEBJgN
jA5sCbprEn2iLZRjkL3L9D72lksO6YqMgPg8ro+BXPsjMD8G1E476pfcnaZeHZfKBudr00OFmjSe
hsqZUQEM7yR/t8k/AB4mVKzfJ5xntLbkRhCkxPKPP3qu2TEseI0t9FDPKQruAUH3kkbxYlUR94O3
3zx2LVDkiKUTvxLOO9/Kh7KzqOE4C72e+EuqGYqHuDWf3ardl8PGta4KIejfHSJivFhWnSfw0QVA
ZbKqmr1Shlsc5Tnn0BYyJIMoK6PCel9IeM04RcyQCdMpT8ybpLh6KIaGU0/Vw7AkYVqqpeBHk8Rn
QvqaQ0/1x4Stj/i9LT9BNG9AW2snT11didMZEUnnDg7SnEjDr8BDDdM4XKBpZqUjURoynpLRNr7v
e0a/ciLUqtPM60gFjD1y2nmz/iD3JJQkyTPRiCmCrnWnR2Cd10oGEO2OAAM8gH8DNCn8uUD5AQdF
CUAond1GGwkGK1wCKNIbJMa4RYx08Z5gJqinhU6aG+/6Ow/LNdSrsgbMmkoZ9YGy4WIgZd2Are41
lqrpW1Sge11i3VfjmsIxPIhPwaK/puB0p+m8qNuG6no1g59OFEjaHdo0HhPxX2wjb/jqetSRWGWe
TCunfFYw3rQLOqyGjOnqOFK5tlX5EchsohdvGH9vaO1GDtnwgTjnAgWJkBCLEwnB5XvYibSOCvfP
B/2sMILjbilhKtl7IR2vtwD0in6gyF3iFeA10HPUJ7G3P7lW4Ev7VZB2FUABjPOs8KZhtB4fJUHY
LdOZp4ZiClSn0ef8TWiaDo+R4nyKkTu1AK+modnEujInLkOIipJaCUblxgecBQn5Xjv1klyBAf1H
2MFTJJlc9f5C5JfMISE8p0DckEqOMieHaKatV/cCcAJVM3rZgCVyK+W6C4LYPxb8812ItVl5KTap
Ay1832j8OknL57SNcka4NxjP5jsG54mWIpWNfXy8h5dJsXCF0CuN2jPyjWBAwxeBsVT+Y1OpXw2o
ioZEJn3LljGwpSRPsYWXjPBP3rjKtBkpBJoyTu4LzjUfSCTycSyofUPmRbej+tj/Dkz40f1IS4li
HsPfv1BRAYfla75WUSxJGZjKUiJQZ2W7nuydYW3OIY2noqZxxJk4Ez2ksKtM7PY4f1HbgoL8SJpM
mKVyVZLRuFuTNratIphRz+jVx1o9xXstpoZGh3sIH7lKjb8J7g/VBc9O8ZDRa1duYk4BXp3TAZoD
DA6dbwQ8g4HvEHrRmForLB6XsHxJm00v9L1DOKEE2cBSZd1B09tgeeX/DWWvpaoEMfcRuLTzxBHw
XzzPk+loDjhJuMoVuzqkcOejIJTBHl1qg1iywK3KdWy2ZjOokWXXqK2beFaP7jDn95wPi+Zl+Qys
OxTMg1r/LOxVXhQMHQff3mSpO/FNarT58oI012hlbrmqtIa9rnaGQaOjcCvmYG/LlcBrx5QCtt7a
M5H59mfjBQnPfNkEf4YqN0zVLlwvr+gAKOqKtNHwE39jBWi7SUR14SKqVHcMQ12mOGq0bkIGaFaJ
m3vouo8AK+M0l70630Ptdmew5au+YIB7pBHglHZGouT3gGu87IsxgSEYLkzEOXaIJHrCDPD8IG2y
bzWsyWpvgeCN/chPqywD0aZhFHFMF+EP30NV+Z6uTr/UbOJbMTMuvubRcY7NX02VgHmb/UMe6X4q
PGAHsknJhXVhi75WoYd0+0frsdDsYVW/RsJZB0rachZMEZhfUvbUeTwRcZhTSyXYDmZ6kBrV1vR3
z56S/d5fcGovxySgqlFS+b5wjAfOUBrzTGPDsgDnuvrl/2THhndt3G90565TV4IZ8pPnwH7clDw7
5BXyY3GMGL6vGBTsrI+wSjeg0Y5LI6+jVocSQMQc4cDH5gSMOT4bBAtSZLDWFMFw87T3B2rDbXXC
TBdEu58ylirYUiVW1QFvNtAV/GqXTBgk7Le8l8sUL9AaAN/gIWd3nRYv9id6pWoQcxPS+sIvDqb9
g3NCHbW17QOZg1clpQJIyya2wy+N1m6XoDhI+/DaIgaC7ZKkiRr67wRvbc0aIgBtJSuUTUTOigBY
u0rtvIzk4fXupIyJ+Xscrd+zmqdXuW7E0Yfq8sCHC+ZqBxiykJSGpZdigUfYa/YaELULKbTh5urd
IuJlAdn9HOM/jl0aTKVUF6IN4Rx9S7krFm0EYcaEKKOdc+DbOWoCsppVBrE7UgPZyeo1UvejuoXL
BKafRIlSl3mCerKfzyZ0LOXu1AFiJqU6jApCryao5RTt6vnY9D4MdQC4AFxpfQhGdzmoSRRH5g1w
Eu4ZX6GYotOOD+WJkYjkaQkKNwCIFcVk0TjbVwbqdYQvteTV9zLuPo8eAkCutCjuD3yWPJGtUuKk
VKt/Btcbquu5GftpdlZZuVh0bGxIBRNshlsWslElxI5B8vu/inWlg3e94oJid9PnWri6tGsSi8pF
QbbmLutnDf+Z9aJvXF/B3n7ziqfrMwPAdsJ11b/OmIRmd+W8fUHsBFgTPhBSY1bWhjPUkuvN87qC
KEBZUIrLJ0D8jENj8UCIaIaD3HtrcFDVWH89dKov/QQSC6thuHJEixjA4yf8rSeKmCESmlDkVkh+
kaGiP9TPD+EvX/9pMSRMGLTIuFbiASMnB23qNj5qs/oUM27e5eBQgodG0F+J9zYa53h6/XUykkbC
FsQ7HdWGlQOicYyLW0MZ3PGs7Kgyw/IePNMQZ6KTTCX/ykIj8ownCukjmGJvXSqzZkcNy1/NsRs4
KdT2Uj1JQVJ50i4e5Ho/TWFQhCwsJPB8+GBzEfJSKZwn0BT3R6J4ZdAs/Yo1n0wFom+HOcSq1oHu
jcZQOWTaJBkXqf4dNAE9EmGjmU9CDh73470cT4NiOR1dEnl78xoCkngta4ayNajdJsbKkz/53yJb
LX7fP3gvNrFTYit48nYyauyU5rI+v2rcw8mVwnXiJMv/BtlO5h1PwvqFucv+R4Eo7/rke231GJE7
3CNMaC5ej09tvISEExSqiJKe7Gwkl1G73bu0eVlNKTBgNFaNQFlIh7E/fMnkc+8yIqflUSmOCLdC
Tg09quZ0IyqAhnzlmr1N8KSMS/zYCW4/USsmKOa7lmE845bwEnX0J2cdD3PAMASr7esJeFzpGFXJ
mBLMHFUiGWqZ56teVESKgZLb8AZwZdDgHTpXe7mpw8uPU6KJYAILAhRA8kVmk6pd45et9XfeR4Zw
mMMrhv5j3nILGGII1NlP9XAuBuAcudqYWPLsvmWtj3nVtc+pUhkkpvgbfu86xtH3XUgsqqTKyFck
kiOB/sqkbW+KHxqjJc4Qmd9xD9dcNYR84GBvwc+kQrrBTY/cYRxRGSON4jslSGc5Od1js0nRNxG4
yTxhA/RnD9GBJN6S0eh8MFXZy9ImlTrWEzOv/8TNjN5ptOdI5TuHdzXPGzL4DI/ftry9uVGoXYb6
Nogr7Dou7cGgae1XPeUyninzTEwjdOA07R5fZa2IDiGlRGB4j/1QQ5HP8JwgTZv3L0tHtRmzob3C
h+0imv1K2FqneWOEXJmQaTmPX/8GjJhdqEUisFrTHT9GoVTPfvbjoocEWt4RJl7SulTVcH7p6I4t
lKzyoo8KaeDedIpWl+E8fiiLzyCwnpk7AFuIEDV0G/Foq+u5oNHhoG0eTNIHsjOqK6fzYwety+sy
F9/0Y3hoBXCVle7nqQOosfCNLkuO+BfWhpByQsMWo3F0mrI0OSp/V+GFv09x1NdXDhnJgGcZmWTH
/BS59ddqW4or2VD4Pe3mheY7xrGeJfoXT5mCie1IlV/ot78V8tuJ2CPWHzfZPQGJGQZMsoXW/r8A
/9BiCMlcwAJQVVjp47/iw7y765vM82nH3ZGTII7lXHtjdjcKqL1ifEmyEtUpl9hIxAluw/Crm0t1
QzzhoMgxAOlMOoD32Yco07uoJawCnkeMn5e6NzubjFqjC97UTNtqd3COx2k2K6BE8zIFkpv9ahi4
d/1xtmvr1ySlrrr2V1JlCklA8rzzb6+V+Fbwy0KZBwE0U74kI1xg9K8OT6+YUUGTYIg7hpiwcS3N
O68qM9sR+KEpx3NPGvggymlfCumpmzFpr2uT3QbUtXfxQcWkXWAAEhioUrHj/KFF5RNmvA3bGgSR
lGT53CWYCySx2iupTFF3EgFV0pq7R/Jd40iaz8mbHna11pRKUwr9or/lz4VQYloobfTq4St4vjyo
/jAqfDSwJv+kIkLrHOJK9oCDfT8LF2J41RwjZS2aEH3fog90MnPFYmVrqgcpbpEX3Kssa6MlEQ+7
S9AEgkm+ETeA+0fV1ecisBqu801aI1jxooXE9XkBpn8GHuDU11q0FIrlUdYsieUrlu4LGQr2AYK4
F8srm+H/l4Ey14kW4NSbWsGn0zbz8rAndDO5bgTeoVQ3WXL1mwsHOwCR4LEv/igA/IjXtQitzgGw
kfWRMq1g4aI0gHOGwZFf6ZA1B/1tJxKq4eR8sPXBO4mIzWNizSDD3U5ayOKfML08AAA1LpqciHrb
lUBuC1mOLh+GmlbQLzG7YT2leLjIE+GemoGqgTlsNIIAHuqz3upr2KXGSwQ8mpflaJIMpWxB+zhl
DzNLMOsWc8Dt5aHBi+BkMkDlBBnnzOASbckvx4NWAnmR8TWUnIu8W4ymnHwTTmTGT7rOlPv2G7z4
akwBm/VuUHwmUM24XJzqGaXPoEZFXMzcVBLIagNTKi19wix21FiId2KNqudodyvs+cyGBpdR5QNs
7m5QHwOu128opf/lOiLPn1aiYjMXRivRTrOoKyRbEeO2tVZVieZ/57GKx6m577JQ3+P5BuGiFt2W
h8wrOhol2Zbl8EzApZUPHQtgmLNqR74OrlAs32KEkoMsfCg/EDZJVvpT1boQmXZOVKSyXfEnlNxT
OI3QuuDGSEgpnijiqpJm6PHF8uSce+MnThNFeS3vEVTfH4LylgOA9haEPoz1/n/WoJL/7VWulTan
akbXkxffOeZDG/Y8njryOkgEF6XCVh9zMbzGokH2xcdn4fAEb1agucor95nkdy/T+fB6xpcwk1bZ
CNjHMW2+JNecr8byjdkuBBUl4rvvFjAgnAVVmuntR981tl/0ZU66rWUrFl0MVrAn6gYquwyE2kub
/wkAfIxcQTLaSQZoDc51d3qUqbP/mDQW6PQhjXm4C/7XZEM8978aMMCKQ+70dIncviWtvi1D1+Ye
XcaXuqNAud8tYLsgSoMRJNVQk6t+vTj85UPl3fo2oD6ntx1rx6PF1ELNDABm7wlEH2L1PFKyLa7C
UBDUwau+EZG3+d3h3916jf0Z7uGKnEgiyMrsNhTpt/htMRgoseforamrgNv+djxkTe+VPygVV2Ry
XrgHn5TvRd4vfur3QdYhcglxhWmsFBKFTXBQpCHHABG5XlwQKG/4UL6l2MJQeqRWEaaC5M77i6JW
wu24SZANnEq1fHcE/B5nQCS3O6bbU/KtvlhJt6r60vMtXWwAmNK3P6Q1IurDq4boi6Sq418CtDik
vDTrSociFfk67ZyHCpbn1r+RLHJv+yVPu+9nA+c7FzrMHM6oxf5lhb8qUiHbQJJ3n7C78Oud1nso
pnd8BHX5TzlbWCyRVnyj1lgUBqGiQaTltvxf2HXiBjGTOqcyBrVbOWkYTRLCmDtS6z+0aY5xcew9
keV+7Q3Khqzq0VgswXMVVMtiurBhwLdG96bWvlRZLNC9JONtTKIgLVzuSB/7sY0QEo+TjKlDq9UY
aKU0fF8ddDW7fj94u2rCEZyH9X7egexhTiFtLZsEb+lwcKzQ7b8QraPK7UEMz4BPbQ1k6PEBs9k8
F65S9XDtiqD5Qg2axxg+s1GETQWYRsacVOYN9c/2YNfc1Pwd7Fr7z1yHx+eGf7halZPt62hAGNEp
no1rLuIv73/5oH5y1D4yT/BRcd1h5IODhndcd19R874teVxuwhiouMi4mFlRnmiOYCxTqXtyDQ9e
nl9yCOWxwoIR9Olx5pVwrprGTdw2Fu+nU4TOFzN5QDLt4mItwFA9Ob2DGNIQxPfqwbZaHDvWUd6t
WdWUdjCjBUziQt8dzGAhAL75m6p6v1P/eiw+0mBoPm1dKqEijyMGDI2WefgqcJ9d6ZnCRwa8Y7RO
dkZIiiZmY60JDu3paBbltLoBrDtJ65cgaDiQypaETmL28GwNNh45zNh83LNFcFPXe2J3QQjZ6TGg
1uL26QC5yKNtIyj3GuXXBlvpaHGmFl3dh1RmaPwsRu++8A0eFHLi9zoJthk6ipoAftMhBfkRFKsn
nwss84zwynN6E/iUx0IJgGwToMZR1RbzD9GNyD5+LgiVZdeIYJc5ioSw5a4XgLrHSzr2qbnA30Ki
XfCSMbMDo6J1XmGHJlM4rINZXaxN4e5HcDhS9j238T17RYdB/l979i2V8hTnAknOzAG3L1jPRF0c
FJHvLAuptgNU7aYvAAEZLWnZjIU3ipR/anfGoTS4ZNqJcmTyaqHZZgP9ETMTV+h/WcKPqtYg98RN
xfinPfDEylX2NnPtRPOcGvfw2DJEFZa1vXe67TyDBL/BikAkSK2Oxc+0MovEF0fxwCzfzv5MdK55
hifL+eDLUNypohjrmKJIs6Xx7MUl6FFgrRupsgSWOc4J6+hztB/iBqFGTJGqFWcNco/ouw/g7qeX
CidKPp1ribVjbQf3g5zlcUyJMOIlz3jqtLYx9wLHVxOV7N8RjkFFl47ZtY8hKs5w6UjLL4IynVeP
DTnbEZoFXWHsd6dTyV8Q1FULcpVPeo3g6q0IJixc+WUc/nJW5bkb+H4B3tB7qtUJ4Swp7d1KAwNL
bACDZVt7/MDEMUvvjxPIWPVrOZb+KGLabRiu6EMKM3NpFaybrjrUGaN7xCh16tbw/c+cWQOanfhT
hZSFp2BZWU0PrqfYb/J9UG97GGq1HB8LzpYzz3ffZ+17RrOUR1sKCHcUZ9dsssTAxhPg2wf2EPuk
9m5VMZP2Yt9MEr5TY382i1mqV9GBHsJTlG226uZc1G+Dy1iybud+FE1h+5LU7+t2WCQBfihIbgBH
uEqRWGRojU0d5uFjEGaDc65LEFYZI/E6k3uCqhA/zZbWojwslSGgL4wdP6eov8d31sdrj5CJUxga
88aV2sxi9YpTkXXdxkCL9KBCH4Gm44Z0ElK9pI8JTVfJm5g+YW3wEH/r+CEKGA81wUfaI2bzIO8s
qyupSRMGp5zFwjd1LCefFvEbz7JzRD7wHclh2zJMD4hYgSwVala450+Ni0rP83rj3ClviXbU6tG8
dB6yYvfJJCf/gnu9wVX1lZnJdaNvSNKh8t53pM69zC1Gmn4rzSLTfX8g2eXnMHzqbyRPAwdNOGJD
BG7DcsCnbwmgqRsqUvuHwPnem3PQOzHo66JMIO7IE65cPwtqs/LEaJl8mx/RqZKkNkJsBg4rlN7I
mHkKGfBvYUZOuK3gLK49w39PRj4os/hWxudBlSolSfKwPmJRPiyrsuCPv7qnhuFyKk9YGUhgWYDy
o3mPMjvEixp90KpPy5Q/RjvK03V8Su8fpDNDZYNrK7safrAeRoN1vjijFx5mCYQWGwdJR8EoWAeO
gdc7chxh2ytVyuCz7Gb+pkTo8UgqEnIpN21FHJBy6kppLpjFg0768xz6duRyiTsdbuEK56OuiokP
LuOlj2lBMcRg3WIeClL51oPF0SYEgH0rBhi5Y6abd9l23M24tET3nb1peS1VHavH16SQDmWPY0ha
8yy+VzxfW7XedxinEsI4gZMDI6U3Uekwwd+5kASyJ+nsLshyZOjtRJ1BbUKt1PhyUJfEWires8gl
fDcReggE3zGLqWQBfnt76cOa/LVhlmDtKrpFnUO+JGbz8DVOn5cPB7oI9mr8MhfUeQzvnYZKZYEC
ajlRt1L0XYVNXIjQ5BRVl3doxYHblNhdr/fyLXWnzMazIga1udeKZs8oVPWmeoTTDrQ90GIKSHR6
T6RryesXIGmsYkNxOkuc87d/CKelAdtrW0BpxPFehYc93YXjjLIzqhJBwT0MQ74EOfRZJLrG7ikV
ycAtm6rdiJhGx5q0UL6RHCTEHtRBPJs9U1i+GMlyC0dKCkjkDClgZphG3pv3m+mHZUV/fWQgsyIC
nsb+JBYMeTompPDCZB2lpvm+zCl4bKGFHCIR+mPseT31o+Afg0iaiyeE0PGpWLx95fg5ztC/r0OZ
4C8zBqv6DH4pFgS2cn6aGZJc4yf8nBuEPBrp9N/7ZVBP6/+phng3g9aRVGu2u1GUwYLJsPcdurZp
GE1BZ3dr+4rDj1Vxpndq2OGgmdcZfCe66vxEEmXzfMkx3PWSZIjuGYNvPyx3rIpUk7yhE+S9fs13
HGCrS9BN34mVufm/erk7Q8bMJW5lx9ps7mVX315Mol25oFvj8mBFEC+hi/+T6XtwCBmaXzuTWM0v
E7+UxcnwnGFYlyIKcf9RCqQWtdgr4/dR7ooukd/V+yL66twzyzCFsqILELlti29SNDOrw7CVr9fw
z8qBniXvxX5hDIig2752JC9QRcrWD5DcU2o5zqs5Sc6JmNvoNtGuCLM0vgz97+19G0Tz/YOZtg2l
1PZmfU9sHdGjDbL7VlnzQsfRYHggTogwkXKhyOYdRjx/TPqw/ax9XYkKPK8D/22ACHK02snbDsF7
pUb4ztukyplEKIA7qQbqUrkeWZttiMpkEQrz+yf5nn4J3IN7zgn75G0qfGE5O3USEOmAJFgj6r35
SAtP3HHcwngHGOdTbNSwwCqcjpfASk2r1nIap94ndcSoOA3M2ObP90qqz9cWEwlbw/qNOHJbRQDg
4BM116ILQs7FbshUR1xAxFrGLyjAW8EaD6AHmHFZJn0zcZAXnR1iAAZiGtd7S1NRJ+/aFw4cq51G
hxexxvNkugcylZyWQcOfDskmWeUIS9FpMM9zDJ2W7cZJBNAaz5K06bQ1bOQ3w2cyA/EeqYzU2kTN
QUtUVVvVxWunr8M1EUiD2eBmtpfJuQvjocPPwUYtLSsK1X8/SAjommD2E0p01qCQk9aki1QZhhEj
BblDFNQqvqFM8gzo+O9AQT52kH82jXMuSEy+mklET/qrPaYqjbcs6ceKwPt5jXDmoRjpYdyaEXyf
AZYS92Exfl9UY9B2bIEpsRCZlhou270Yy6MeiSouM6xtTR/dGL2pfqeAHCssnqlaKKVxYl+KaIlV
nP/wRogVOzWx4L2vu1mwzVKHq7XfFsOuj6sE9OaZcUz7Hr0J8VFKSBc/EEI6lEhve1Q6rnGZ8kPj
28zBydtg8XXEzbMRrGwoDu5MhsUVp0hQrScvqxQAvAXlV3N13RggKvwkglXskLVTgF4ZuuggLoFX
BdMxFpk/tE7ZqkJyOGKlVyeQocFeht2BrSSvAmbV1QfDMqUUwuAtvUdqH/5ZMoN+/11riCAxsgXC
DbOvkXoV/eAK62hl1hhk3kyVLVdmZD92NAg2j9iVeyWCH782VbdMMOyIjm720OOY6SQUYHwH98uO
dBzzj6bjs7eGDOGF+00RCvYGzG3PsG1f9FjmBRO1zgFzb+WDpVaq73ynYo4UJL4A7pBYGIOS+eYF
Tdsx5jDMJYebBb/7kI5jqxpb+ZsNNa8keReDAV3w/igIoPD47OMGJjPJLtzWHx5FMm0tQ0hoWi1H
i47kEloqH3IjHTpKqSxc8lDodrvtitCJBVBQS3Vvp5rpP1XpyYfeRI+hT2cCkjcrWHmX8AXv8vSz
hzwr+oqDtGO4lTBCjfik/wnRG5LRJFqXeradmtsJCsiVbHvz6M/UQUtBYi6qljoUnoZXmNZmNyQI
kauptOtiB1Y2Ei3Ev94lF6hnU1rvXkMa2n/aDPFkNGBhyFJQ21j9Sa3i7doXmgg9yk2tI5ghxC/s
sv6dWXqIYcEoAaGxc4cvBq7ODEjkZAdME95jLQfWd7omI03y2SXI9K1VrP2/Yy/U8aaM9ZSFXiUG
/Ix92SeTF/Y2aMDq1zUyPFiJGRMMTvmnioJYp+N9P62t6qWHsmQwXIhj5qqYW2nU+fMZCtqdzyLU
7Dfz+hDFXh0N0XAEMGw9oTQVESK956WXUdUQIprjp5+6Vs2m+nxSwDM/oiNMOZTarzeFPKV+DMNY
9+fJt1o8cMRJr5D2kkUs+ZAvc24sKAo0ggS6cdGJLDizp5N+MTgMIKjFwI5cq1UDI/D7f9MAX3HH
TM1k+Ekvf++++mbXcbUqlGVEoyu3eiJmuMeY32iKHHHL7wz/AXqM7gLZFreNOWYBuERRwScOhTwS
s0WZnr7F9GOIhY91RS3cxgsdEMmN0JDPbF7Xg9pXsg7+CbKTXZDaXVz6s+s7pX+dzQICMsa5xNco
Z3MlvSx5OKW97rusFXEO+oEfqi/2ZwUW26WnbbOeoNIfG9w/3lvkXAupfkyOoSkeKiDUYTIYKvxa
7AqnykOG8UPy2wZ5usOKss1wT57vXRTISUqRPdnyYELpMdSqPLR7jq7346vsiO08fdBknFXywFgw
FCbeI0qgN7+J/4d0gN9Ibcqa4BiGzg27IPsUMGj+HGvFCR+MlYDh3Vt6tgxSPgYS2NaJ+1cj7Dtj
PRcYupjLGbjFIREDz3Gf2xJfafoHPgejTwBcUTSmYejOOhJk9Q9QxvN8HdV2i2vgb8eNDGtipjqB
mWIJCsCwL51KcrHw/MPp9YsUjZEfh+vFO0pZjlhBokaz+z2+GvPejDUVkcS4PaQLaqlIXuE0VITr
/u7NGwO9TOCB/BV8vy2L2VaaNVoryDbi7JKxOS2OPO/CDhr3oNE8whq/4wfpZ6GAquOnzyLVYsBt
7DSX4Lmwsdg7F4MT5uR1Vb4fdT+QwIUHkFGLlKyHLfOrvE6EjBwGHacTBwth66vknjvaup3DdP7V
J24BssHPY8ECG3qbNLXAxMAu0H5LeVEp7BtPAFtqekrQpGQNHL2XwDsgFIKnqI1GHzbtjflJz/W3
7gM9V3xMoxfjDDtUviqpZm+kCGNJIryhAV8vh6cYEpYdGYF8p54H4PpW/DEvPdqTK2WMNOBb3/6o
pedkzDr0okqItCgkVD7K3p66bgMS1F7he1PQV7hKYbnE92E6Bj2DAcj94LXbbgWbfz+EtSDJhLdf
VwtQWn6XudYnwTAcw0/mKhaw+YZkncxV65cmOHuAUo1U4c6uSFN7+hOk/uO0IqoFB9HRsiQ5x/9i
gowsZnjhyC5qWF3gU/g+6Mf7AvK1x3XbzGfhj4oMRMkz0T2psBkS+7tH9Qgbp6LPFbjYxiNXQkmM
kqOzVJWAvZKclkrGSwHHo2v4UBVa5hJZbvZQwraa2e0Gt7iW0qxwYveyH8ExJldEwuQafnvtwoQx
53e/pjFh6V1cOSHneQ9z3IIQTKuQPt/38+ATF9eT6TIVWY//bstmAUHtKqCyF5mG6v85pZ3+4Nd4
OfBQ/dxe8vIpsW4rIUEYSDbryNk0dqOi4Y1fDsYhKALRRW1z19213qZK3XER8f2v+g26cBaA0RJd
RY5yuyojrTaK98/EGsIiE9PQ+0V0Xo/APtEMqUmbPT2GWd1Y9f3J4ncbGsguX+bWuS7902IRShP0
SPmwtVZHu8OxP8bRewfEA14/ZqsMVVEZmP2RIY/x4UIeVwemHM4y7P5Bid++V/7WVS4KUIc0FPAr
FhY6nYiwdi04PY7ExNV53nSey5kXXlFF9fbnCrBILBx9wT8fhrG2yOIcJZz8gR2M2jl0k9MKTvlo
OjGhEiPKVjIHOon/6gps2IG+HI9EBUFfsl53sY4iBvi200Dg9t78iGuZQHX2fv2P3NVYDZ6G8isD
k0Fa1FOyLUsUpB/9L9OTxExx/jb6EkSVw6nAXCsk3UTQCQEVmma4pAm1nZFjTIGc6W0Th0M3mn4Z
f+y59cSGIMIcoJ0Oo/IjfIaicD0h/LS8qfVlsZQyFYcqgbgo4tC1iCa7XnJVafs2mSnfY69Yj5J5
Q8UdFej2CxenhyNnVgHtHu0spNymPSBXrmQpgY9tlmARLCPwKvKxxgSuWvapp/5HsFUl9Dx39cuJ
YtU5QtxulHD0zlIrtPGq+XBInibkaDttr3UyTne/yrcqwK8l9jsSASVdjIqglTjMyqY80OHpXT4F
ZXnC3rBjw7nOPmccB+X2zcNDvh8mbFnNpLdLkcnSgTgM/lO++xjZTdW6PTN6vgeIXG63m/46uQhf
t8p4IsjIR8uidMn+3/0P1KCq2dRAmefFPuTbOXIXCTqvx5U0zqpIG8Ec+pXMXtOmtVsYOqsFR8H4
QJIAJCwbIEWwIgNt8WW2V5cnH1DhtEm7AsXyqsRIvk4l1/y2hSw5JTuN6lJs+ZS7wiCi7drLK8UR
X3G7qpB4QOtizSmL/dRmjO/evHzrzKY/++gqh5f1NXETF6EUE/Zvhunh7+zxZCxgxV6iNpMNJIPp
3STf14MTU+DEQCvNG6sRg0P1LVW76Vht67A8d4LELtDAvc4SRyuzm9ThIm2Yd6m2hJQzdHHV5liH
awHmTKJGFcXy7qn6pMrh478FWwy0kQXZrkfvBG9jKqKk8R+AA9M6NoYGHlDWxerdN4tYwW4vS8qv
FHe1FAdT2BW6aj1R4OxCIuACU8YCHtJ6vJSFTlEFkEnfZRt7PX8FYipZx/VffCzoTxPfepNAD68o
VF+d2qBEECM1M5gD7DJcmdKlxmxK7YdaD2s9XpBc8Jz00EhkY2VK1Y5Z3GgEiMcxPZm1JisLfNmW
KYO5xtjGjY52nSB9iwXUT2EaIxeanlFjzAhzrxraQUfemNxRdQ5sJjVyc/yYQd7A9JlcPpwPfZT9
fL7oxtmtR1dmL2wbhQc3L6wTTpxMAMHY7EeuJlOz5+RIgX/9xICqr6XFn/C5NB1E/ULDHQg7kfUA
b3KgHhfO5sOJjQsLt/ukoZ0ShmYNFiZQRkuWvCXpxnDZO8LDBzyVHhjO86UZETpCKruluECfubjd
hQBCxNzYrWLOfPpSE5aBwU2/X4/yGPP/91ve3hJpfktzhpcZO4uSCSDM+lH6blPqqhXotENkX634
jeEjQFxfWxV9Q0DDcuB9X3SBwxvvGMsBqlXizLRUbKl/TVMO7sUkXksSD+T4a0/MkMKtoqYZvlqC
2kj9LNQVluznJfff/kuhZXFAQoer352j77Fze1/SQwv6XYGq1vEiUxNuzU4EuAYiFJRD93qMPJKO
bJKaTjU5PKczH4h0VSNAgRAGPIQhJI/BbhAwajxIYkoSv8Vp1kFi4czfRk+K0/4hKHUGp+rnKA4t
fKetY2gjaGcUNDZ4uJUV+bcNjQQyD/cK6H/KA8Z1reuVm5xXsDNuWUxm9NC0kuKae36q37H/U36q
fEP1a2ZePSCmq5v40USg3ggbDXFAYmccf+/rAaJzxogp/2X2H1T7S/ZhcKdUcL/PJkQ97zAO/VQg
eVn6w9I47TJSl756zi7AvQjoG1XgFkL8ZlMrk0UPFsjuZfpF6U707xtGpOS9MW9YCm/GTzHoVu1c
OoGjKQgSYLeMLLLX1DParU6KAL6RAGNMkwPO2nFKJtWQc0bh4/Z0O3rDeBYYRCMa/CoQs/+TAB4+
iuocyTcHT4dzseUmGx03Gg0CAQ5gkgmuB43L2jAwCqk1+DIu3fyqhVzKS8841ybBxOxG28vaxCrE
PNONrD+jp3vZFDlXFRC74zBUrHqiMrwKxQ5LJJwXkcqsTB3p5UcFhgRNYj81KAeqlbTTnU3TQUxW
pOYpDCCv0uC/8RGnHqTEnrl0OSE1/iEm0H3dhj4nRor0DpOfHUZncJrUhtxrI9DsLXKoztFR9gPC
J3wcLCrAoyJa1o5pkIhw6rdPsiw7RCmEMoSxTmWFvjqYrpXtWBR8FDO6hrI5za3a9SyG81qyG0Qf
fANzBUOy+Nwgtw8GC4/LnQ39AlhDQUll8v6NVM/3XfIjdsKX4iJCnG1SKG9p7DWf4GvxYqFnDrbO
akXGMdrpn/s4PQ4+YJ5oRAkW8kWD3+yT0R6hGlX7fiI7FpBBZTgMAaTtHWBpufa64GYCrtp3Jxqt
eW5V+YL7OyJMUmvQt/Vk25xHO42xqQhoghjiIT9PYgjfABZIa/NLl8lKWFlP7u0Qd6yjkL1X9ElM
ju2H1JxFpNKud5YfvFjsqyN+qZMfZ9maxs3houjekUEoobk2VTjJgDS7SPbWIqUZUrs42RG0aagX
xUpyausozFwORjAFkCcT4i2wOoA+8mvPrfQsNn4YGKghbVsNlaTstyNZCpN3NA69jo6xLAeMQLt9
WiaQwj/CqQIPPngkffIw9D+zmraEK9K8fXwRPrVHMLpj/O94JbFnx4vH9aCR3pCjCeU+rsp0LJT3
gnXWKCezIkbjaLv7Q7AoO1KDC08AI8IQMdIC5lCH6avv+XmK0Jg8KIML1T6Pm2hyYLXIwowZwD1t
qzFuyGPqKIh/iVeLo/+5iL+PpYJT6A74RZcS71H/mMHkEXaWLikxqkdhjBlDb++Oigk34fUWYn+P
vfq2ta6iMb2eYxI1aKBiN6he6UcIZeDQGl3+zRU9D2RU/H9zMliSMZjAzawDHHw/PIr9C1PP8e5a
YMvnsBOXYixVEFvfxJreVTYX9BxZZwRvKXfwJENf+GMQHjkVFqOC8sVeAMV4c1ymKTzDUAqWJXq9
/YYLI+ZZvpvNeR6rKoXTfHfqtRFilGjoC34roXs4z84hiMkAo06E8N0AyDI97FbxBvHN/x5FhqCw
QrYH+GsKUxnUiDlpOHEX7B6zSvxrPeL8o7pLgxbzvgFLIoWfnAOVVtab6dH+SHFVlBaqJ1ig/0TJ
w495wMxYyqXh1LBOtTlQJZblie/mIA3AcPlslFVTO7tSJp5ctqp56RJgLX4+ifyotwYrAFwFj3S/
xasnhrBHCmneySSI7Glti1gX6nyFg+M3IYT613kO2C2VIUOyOWCfViLWl94yRTAB7jn2YFPu7isx
QB2kLdDjKISIluBLulQPVIo84Bjq+aOYnOMM9pNQV1ITaLZAML0j5BglWYJ5wrBzXuiGXOnmU+wZ
vAD7ZLoMsxlF8bZjFFTHcZcnml4KNHFgC7jK8tKSJDYNEvjqpwd1gi9DL55kSz24C06U/Zw/ce+m
2/7Mea5BHz8d82bYqNnAP0iYNcnfJAXQYasKaPJa2pgYoaPpgFJRvyTCpfHAXOcydHCLZUvMrxsZ
9J/kdlHgZTG6aWj0+GBAeJvAgBnz1sFOYLbsBFkD65IbPkz/WgQPh6YrgSWQZYvD3ydcTqOGHGjF
uW2E9lbHsuFMJXeBAqPMKInm3q1ieQIJb5zl5zD2Ss1TdK/zd8HY2rv+uU4FfZqIMaow5Sbmy7Jj
+pzYLN+tor1L6vtDPSIsbJ4nKp2L4EXcJWxvj5vyHr9dK28CyHImum1gLW2YE9aTz426PpLE7t/P
l7TUSxH5UW4lGDJtVtaDIdAt7xjYl2ZvmNoL1TjAT6DhBd0zU3tR0+zViiDP7bP07QXntWewoLtz
oULPx+QvmYQ7IVmymcPxOw/cUB5B0FPJlH/suk+0pkxDgiAfogt80/9LrXiSWFrI3wqI8N8JOX4h
irD5FFViyymeiVDDIRNjanTFp5ZBzk/RxDM45BpTmIIZSk/+y+0cILuz5sYZOG09URAD9c88drOL
1XQ6RfRkrkZwf9bSNVEV41qw46WfF+jCxprRiI/XXzV8jh56qtnXObReDxL7IG0TSVzD3jSgc9hi
LZZQDT9B5Yya9sd+ZshCkFwyKi4pRmijfXAPI5D5ZFaD74+0Ti8p1DFR2IV9Fa9zYwv3zLlH8pEj
asCQEHS4HUC4ROOXN9HIFO9JRyLh/ky7mOLHce/KO5Q8471OBFutFu4FFHuDQT0HyJ4lVDNHWXnH
+ehKm/QQ6phJcyvpu+ZtZAYFp7fGsLJ8MlDXJ1C1u8ayHT5dZPkaXVnV681PiXHVxmkvEv5OcrA6
XxeHMXvwsEPicXOk6LD4ZMnRDjJ6BPoKZLyDwu4kfyk73f1xHgWs3SOfTzdlloJyKqnvYbWZUqFc
oMQG2uHWBrUTZ4F6UtNn1ip7l2l1ZHrXARdLmadk0TvP7Kpb3r/NUaL8n/BihN26rnYpzM427xph
1m8R6SR3nkYEGtDIxyU9T+VKdc7OjR4TXRd8vf8a59TihL/UA1mFCinEg+TiOeOofNNdfa28Us8M
bVBULetKKZ8IXRmx/pwJPlku2y6Kq1INJGynH60eJw5pkBozpjq2yU3KF61J8mDUATw3fODePjD0
xG6HdHeyMRhzQQU+Hm/ioMYUhdg08GlLHa7I1l9l6TQH7g4tYXmRGbNzE55Lvnuv/SOxDVchiqND
eRCotl3alJcBtwxKDK43xnmLnIIlERtQP7mpNMIqrfyzeyvvoOMYUceDy0WoI7u+O1CUf7pd6GNK
t5InRp7K/TWzUajVww1LJYL3XKQExMKpmpXy5mJcp9stirp11e1cyB1YI0G2UB11tFO7WxG6GBYO
81Uzfkqo3G2Jr/gmERTls+IRXdijc0On7+TtVaQUKvYdy/bMWG+4lEXt4JaTQ+uL7aFUabbi9trz
1Sx0lXAEcMF5iUDeTWDF8uweYvN/glo0v7kbPRXXzx5TvWEpEtEUDMtn/Jm/7Wuwp1m5YlcOdRDm
M0G2dVPzQi8GMauOh5UeGKJ7ZJMrLr2S6c14vbBHp8VnfGQtc8pPhWCHwY+Q8FZLS9zIih48awYu
IjzZwWtWKohEmRjdl5Hb2jZ1rEZimQJ+MvfLgh2YlFfpmZLcG/vlkpYwaGdhozVC/XPtO48ZvDcT
2NmIKy1/2LqXtQ9cnD8V684Rf/MwLHjRNeB28LD6s1Mex3VsH+XrYLdnDfvEQ2Y0NajUHjE0g4EC
7uU4XYu1GHHQgVzdHMOOYSYGcCZhPClQQKBIxsMd2e1FxhWfaAoNAKCdB+xQ2en7WnF+sLQ4yDTT
m09BnnUP/cxpR7Dda8KwZOEMOLmi8fNXq+KVwzpFZb+AjMXSJ+5Pc1TXRQGFtg4OZITpQq8uJ1RP
ZrlcUZNqJQs6/j782OaPBw+AVFHQexRqyTSm5PhVeusN3LW+VKbbg+uqJr0TFwB9x8Ko9alwdUMt
EJXnV3CdMiqFwhIImyxjiXy6aGXgG/qSp7tUOrP/RrNnCcclbd0j4BGzcyNVs/Zkziv9M9tKO45z
55vXpkfva7tOU1nCDRHxwWykoVe6IJj6VwDRxTLJ57/OBhFVrrIXv+CZO71Z35fXW3O438w6TM3D
Q8G+QwhbAQfV/F8VfowAMPFk5tA7Qkxc5B0xdmjx3Vjm8jWI1n76G7pwywLYEOIo6jIQAgSicaI6
vp7nVSUPoCC0Vizgj2D76WiPyGqow4x0bgSwPWvw3d4ijVBA62nYj1tJX62z03uDMxdoBThlVXbi
56OBjBbHPScvRMb+NTKQ3EMG1mCQlk1EPdfKitPq3YV0L+RjBa8bSJf0zkfLoA6vmslvtitgh1j5
iy1ZFi3Ann47jmaEy42MUsdn/cS96Fs0dga2fH5RP0WrI/5XRw6mm7iw/7S1Ee05qO8hu67frMO/
BYFnrANaWvAKona/CenDhxCBCqaBp0sZ+/qE/ZP6KaU08Xir0X4I09g1cON1FntKJam8bERqdjVD
TfMrJPagUpE7cYQXD5w1ci/Wr28jkgInihpV+ulK6okaNxx2ypm+5vNIbqUAGBdI5Ttzb2pJvOuq
fGUAF9wkVdlqiO7dtz2e8q4Y7rT4k6hLx6KTTBudSNDIy+c8wJf9jT5La4O8APKW14Htw8c7vmlL
XswjMFsdbhV9q3IlLUEznyDuoCgbKMUXWhqEIOxfY+a8puK2oPrVTsv6ukqfjRNghVmGeRxmxfeg
CTIRkj45tR/ecAq2aS5ew+auf/DbcU4OENRbkC8ttWFcYwERsoGwkLcc7orPwMwlNgqOkETiW7rQ
b6grz38wl43sxiCuAU0kn1MQVkrDughoG23WKoAej7jjbASgr/OArYh8bHJ5hepE9iWrzvceiHNW
uSPoOJKpv97UtRla2HD0k3iGRE26b4I9GCYPontCaP2bM9pudp8rJIFid4tHlrX03y6X0LXkCVO9
S+3iliWQh/TUM4Cfdw/G+QgXTJqnF6ouZShUZ66kZTN+iw7c5YU1o4XYtJzycdwUgQwKxgtk/Gcf
F9AtM51e4E9nUCjL1aEuki3reKqzzoz3cZfotOUVEgl3Y29rvqKbYeujrdpQoeDjbUzc0dhpc+z8
DvjmwUuC7wh8O4PJwZz/0yjb98KjnzDK7xOgeCovwc1lWNTLn9RXy2NfIrm7GaYqGwCDfZlnTMMv
E0VKsLWhmZ59SGKnUSZpbYnO2WZYw/tsypZFbfZHmEIY8jelF7c4dtwbEsddKtPkyhTuPrQz7eKd
LxsEmeR5NDTYDuDn32Jy0itMH0PIzCIm8oPuoi0Q2w9go4IILTQ+HXjlTW4HclVYdEO44LrXy30y
6X+rna9z9GiXb1JnLL9yZZq+ec4mN8U3Q5k5b0T5vnal/OoEW2qeE1aEm6wtOa8dt+qgj4FMaWm8
wT5U3L3IT+TM2E24aDmWw9DLZpyv3AQvC0kArxqmKnP7uRUrr8MWQiVTa6gADFUuQ7u7h+fdPEfk
XYGF1PK39KzSHtpKKCTW5WPqfNQ1Vq9ESC5s1fq9JYQevN4qsytICJIdJVx2bkhXe+rcGxMxnTiy
HGPdnWE3S84MynweE17+0AzYdI+6+I2ZP2cnhoIFVDgkUDGkwo4OYCmsU3PEFsBbfMHYMP29M3CS
FTfdHlccGWCwpjt7vkL5dK0Ox1RZaXn4yyNHcuImgj7a6AXcCt2dWIX2kFxbeCNwJtSa/inkSDK3
4EChg8uAfT5p7KYUd6/gSh/hBIFiz3pehRwahnUe4QCCxglNHnXw8P39fsonxJrQbOOSSpc75YLI
5UPnv0eQ+h4lZlQhs7GwMHYSlFLjDl37aoThh70LtRLDUoblS5EU9lRxG0JukO5i7Ny8bFgxBKCD
6vdMPBDYpANlrujBFHYHdz159k6CSGIZOq6cfkOt9vuCdWilnDaYdwyt2pNG4UIxaMhw6/MMgbhf
nVV8o5uiuQY3AzWrKwgPtZ7lV+eLGcGaZGo1dEmo4z0lXJsGMJ7J/6S7UQmfBpouyJM8iEdMFM7y
At/MC+xzr8jpmUihocD4XUbk2zW4rCg8eO86psLVRrk4e/n8JC9BS19RJJDoq++4Wr1QkcrXidoB
9ed4ss0fJSMTEX0dZqt/57MTEIyXbnRDq5sRkWhfONmMeKSC87dATruIGWz6UDRjEKkfQPkNK5Vq
VjEyi1gXztfRwOXwjQDkNvC+Abg0EZztw9UbmUnNvVhjkE0YFqyFtGDoyn3KCyP4QRTPl045rg7h
7tWCN+tfCX9uEu+KvdM9Q8R7e4IGK7qJ38WzTjthw+CvUp0E/jvjWVLbyXrFWxr4uolZCZ6fmz42
eRnRdY1a48Z3Q1c1Nc6lz0hJIDRedZ8DsJBV/5YK/kDjOmXWwrDPFv0pthT9nYiXLwJjMbHm+tUS
E45vx63i8SGlI21sBPxppFZ04PmcYqJG0MJ9MOZ29be3NG3BcuxZ2zXYPzHQQhxHrupBIJ7C/b7p
/VYZmFncyeck+q4V6y6WoMEurnaPdPQzdsXm9l5K2LIPrapWW3Qg3xy0AqLfwtxGy7CG3zxxH/oV
6BGWtD5zFK11S2jyn9G1Ql+Qh59pjzFz7ZD+TH2/Ao70iFc2HUsi08F2Luourwe4K2JXwXAPEFdT
wUy1Br1a2OnfpEYp2cYqehkFJxHpMlDChx/GhiD49EerTc9UdoBmZyrqW+BUhhjHl6U5V3+OZaYx
rMbzvjzDemPrXL2OgaQxGtNGH42zqNEOZA0UGw8LX4nugB06XCVSTEV4vy3lGfLpmN5FJgpBlowb
aMHFKypzT1w1mfOHGYNkY1DXI2rq3YWntCs+TX8Wi3na7UbfGrSmaHVg1BRLmqcd0nWizucoMuI1
hdVWwkm+3YxmBQn2FrIWsNd6hpkvTJqx7XeUZ6A8tT8XftQucTOWLnzGLEngaANNOQqerabJPF58
xKqWqAFPSCx85JHh0FVHbRlf0b7uCXuF3IWFK4C8yGe7C/+AgfNj5rrFvdBt1QM8+DgHa4ExgcM0
WqDw9BLL4pgfDn8Qntdg1NmeS+8USqHIFBMbnP4E2d6V1ktsP/NGQyAbEtHSMnx1Kqcj5vTuUf3c
5CnzDwhUtVK569q4vUtEm2GD2Gml2AIjsLLkLrpEJGWpWreDWlmfFglMxNxhnpMkSkU/nvXpQqxQ
boX7zyjsIQM0IKv1BkuRr2L6owTh/BkCmzlqpNSsMM8XbADhoC4QemEHvPJIgaifbfwr54rydOzb
NuFqWiA7XHXHC0FezMJ3bVNd9PQ0cMx12LO//q8UUhTnVqiD5eqRIUhH5OUzSDZRuR1a0WuKXriy
pYUGKhBERq4B5MMsLq/Feu2y2fFduggQoaf1WQvlty3/gxCQrQHkoqivuTMjTBaiUk+ZGTmzBQom
3TlpYUdUeP8DQveySdQrLTEWL/LzrH6B/r7qjVINDKqTKuPg/HhUVx9892Of3X7VWjmw3BgFKm5k
gCxONQcjVw9p5Cfv3woJNCJz0O9/unzC3WMOD4sPnpIz4Bym1YY2/Z2Ky4rzhyzE4AbPx6IlLyI1
yf+xPQ8w+yePDl4zkuRld7FXY69IqsHLO8EfmhvKRcDrhwkp1Gayal/DFWeyPHwX39lWiDigAM05
9+5dIvhsQ78us6OlM/dZKlUekUa47m5t+ktsFS3hHt6sUEfGk1n0kbc9kCAzdtO+UXV5SnlOkxgy
+pPDvSlN8Vl+fQ0GkxPG5KmnfYex5A8aimm1oh1FdWY+Ihx6wnJ0TwZzm/+hd4J5Un5F48hoKa/P
CdBGXXdnmhdhhcCXgNXOcmJLwNfm2g64AwMzlxcKZuEF1F1A9GkhZRONCfVisetSro0L3/x3WlfT
dQbfgq3s9i+PWH5uvBsm3UmSjC14sOXDa1w8SVm9oFmXjw0QwhmNs99/+ELMkadI3+VYYCslMDh6
AFBrWHRH0pzwdyrNn0xqDfvV+d6MEqtnphaYtmHQjYSJN9v/9htsfqA2CtlHvOPhWncGEfGzy+UH
ckde25IpDGSj87KuVKw2a5vJ5lDCgpsfUThgxorKRfFMY3dnTmwJxo+NbE4gheelC+QgCrBgyzHZ
sksQqNYvB6mQ6ip/OLsANr3I16s7XawfqhTk0a9FzD+90kfvfn9FdBj6HJYDpZlAFhm/sAVhhQyn
x6mOV7jc4aPBckLl85Z8D+7gM9R/WQYXgjTYzlhkETDUBcG7nh3sD/3fXyJZIFjk9UAOH6f8EQS1
8JKDlazxPBWDrxvgvGKoZzcLhAa4uGHKZkNs4gAdIu+MF1xUUBIn6X3m0nZo4T9gSum0t3II1GSn
6Za5juXkMayKDcsBCG+mC6uMr5FfzYT+jj9e/zN0L24wX+d/2tmED1rHrtTMH/WnniCbcLbsz19d
oCR67xSz2NN630QHoZ5xq/+Kzj8bo3XlJYfRas7ju4JM09hCYQjxJaE1qVJM96yaRM/dDQD2V07I
LktMpJ3QBlCXDS24RaX6dVSLfTy+vb9SxCjopSQw/oD/b+bulzXPTxqkM8UBs1RzleTPPrjBgNW8
B8TVT8k2VdzCvcvZpOWIMBElNUTw9vil7QFzAe4f/ob7sRTw1UckhTHHmZkOvouAoa0KLWl0/p+9
SIdlGDwKjkR035ZXEcvIzCEt5efinU1o5obC9/am8Sj/jUH5SOJ17TxRxeFJKXS7wrxJRY0EiCTy
L1/IcSwygtrlgeQgb0gpsgNKfWyDBRhh9K2wrxAlC1D+MPTKFIJYdOWIl1vkKfvPL+jbCnn0Fdpm
cy0vTWCsuhuyzhpdgIhQUcHvbAGMsv0Y5foTpmRRZ061v/2EHlLy5s36z8eUqux6dXgu74k3Emak
Pi6ej/e2kcSKFLaIXjIs9cG+MguZ1gdCeGufNagCoFiNyj67o1WlDCTXrWfMKKxWun4f7NblAeBI
yOdNvzrEbbzqZtFPZz8Ga+tT+bsNzbNd9NrgmH2fcheX5tREjXBCoYgpGgfiPZu/9CfZ504ZijRh
JfFR5v/JJ5DrS7UM2GPjfky6HxWfWYtFK0TDILwRAs/aDgRl4S/b6zS46AeiP+3TCZX/mFavBJGY
Cch8L/Xwtrt5BgljgTgKLoJFsApEg3SLJMIrOrXsbd0t3JlkbCBgogtWKLN/ZwZ5DmevSF65HLZg
otRTaPELOyB5Cwq9HOz9IlAGzSZR30yj+nzRyxlJtCi5nQ3bV2nB1Ggy/BhbgbCBKduCnl3sA2Po
k9Jfh3IlbcTmFvrR7nFRtgdKDE3UnYWB9G9gCBNV/uvfUw83arb4A7pXDvyNuZ1jgpym3XdhWaIp
UtAddB6HiCgHxlzWvajCoQWvd2kq8ioKzvVdlevySJS/JONuARW8wpshCStaxD0AEHpWU2V32iPv
vTuCsjJstiP53NNIC6JcMTwRa0ejxIzBSGFSD7EH+JaSxf2IF6Ptyfh8B96o9vjw+YmY/oK7+7za
x0iwNeJs3DZqjkwDRlCul+4daC5sbzTe6uSy9ZNzfXjHfrd1MptrinhFuswTZv14dwYYpPOTx9Sm
pc8IGejZ8hkEv2okU6DpM3nP70VK1XLkEtDnT9SZVrnxf4/49Tyv1Kw5zmfuG9sr64BW1lFJN/+4
EE7p9bC55icoTHyIBIucM9Q0ZNl4y9qJvxvs2juCFTbf5aeKLpSCRmMN+Tdw6qgkVk7GUSIYscDl
8x1aoTMoDojWGFlittsm06VXUVwE+3Ok21rAFasxWBuVB5UL6DygewzvFVrNLLUo9QG+kVEwcCr2
/3GxfP+uz8Pn/eAi/eW1VEdTLRMQjU7hRxlKqsqX06EX8XxKt7bXKl/v27QFy28keU37bsVa1reG
rUGhlT0LPvY2OYCvm9PsRzWk6ULxPEdMdfm3nFaC1WOPrrzIsO/k/d6cfaqIn3fTfQbHG8Hjz4Ag
acaHBRZ7MBwYyhNpdBmVUB5TIYBU/Fkg93A/ZPsDjK5u0kCjnUPK8ykG0XuUAGeCM8OR1Rxyrntz
jfigivtx4dyvOlrtRYtNSgSTl2jECCnxJcmzd76i9BmMI2CSt7eXHnQ78OZS1NWBy/bkSybJCNXm
e6Y8r52pZtgnoIVP8LxoBNqNtKHjLOzeutk/CsoXHngFoi4d02xQ8ZnOEydLPGeExCwJPO+PY5J5
B69WCWWlKkFoW4uSYQF7AOZ7cxBEwK+2Hwkw1bKBPVVC0g7K2hz0H1SM8kz9Ebuf3eh5Rt8eupAB
FzuOFfdHSFiCvAtt8IaVwtJhIk0dVS50va1q8hxgZEnbem4J5Veix0l3YPEjSPFlznzQN+npW/tC
2avU6TV1zM3eJDveSxEFy2hV2cWLcaHaUltuIiJK/widT4tR8kWtd9q+RBtyMEZG9ixq7uwtmaXm
zqyAxsAzl9H8TA2Fm/AqZZy+LxBOXQjD6cPpAIgGrZ9R0s7WZ8N6CqXRLAuZJ9PG9ZLJqypqwqiB
2NSwPr7RNWv9heso+aa7Y775g6rgDmGrhFHwIgdEfxBGR1QPG9IOOC+p/Y9V5pSVieHv6oppLfV+
ZZxuTKR4OKNS5SANVt2ERazD1oYKbfRy9j+gTB/KeA4DC1hJ3L9oc0SqsFf5EmiQuPR/ecxBCYjU
0SXgqZ7qeKKfal5oVMtCcralnkNu3w9UNOwUpWj99I7iA4KfmNy1ft4FwFcf9cL1K1m7bc7AEY/u
MZDKyvcsegL/YG70BJQgUgKEFiMgTDzxAPXun5YTzlYAKmOAClI9NRr677j/KN0AkMmdC/c62TaT
tfyTyXXg0PEgNrk6e7G/boNRLYcUQnicwcxKJ94YlZa/U5VDJ8LuU5l6k5sIzaiKD0YMRuF3zk65
yHwCtmI8FligYYQBPCPhYT+Wol4KSFVYUGH0nlLzIC7VglUlWza7C+ysMB35GCtfyMLNlvjDBsnV
daDkP0XC6I6QtsyImn69I8wRUgnWRbGk4V9797X0RpahRS0EG3Cfn5FWux+ScjZzT0/CfXjjlF13
bWonF+V+D761SpwNeaYCOl5Mhf9TU/HmCb4ZCfZG2ys7olHRL/lx0mMs0bu6F3iV/QNEJQAiIpZT
pnDZRtsT1NkZwg9u8cJF7kEwxRN5J78X7X41VvKm/LsVxhVzS0s7ONGY7YuU5EedxUCENNGXiBxy
GZAvIpJsc0IWymYBlYX6QoIc3oGfEeyIE3kjtlOL1iWHPKG5YIeepvkUKPkBdlNMOC6c9+gqbivM
FSYccHYNEi4sd2ciAmCxY/e8eqxS8i8aiFo2SkuPknS2vN8tKtFU2qizxD+okSx+nXtZWNm6CtsH
NhiqapW+wMO3yewq9ZXJ8WjAzXWhPa9YSiswS/yVM4YMerXA9GjtCy+Fk9e/MgSjQGwAnGJXX6kD
uiwyzYWdE56kVDdn8ftcQuTiKFoTQoR7bxuy4J173LINon0TFpJclliRxF6kz3dDrHCth2k3p0Qb
zlpH4J6QRD0o6q5Y4cv8E1bESIjohi4/Eq7nHnd37L/v53+BT3kZXfVkD6l9ddAYe2QcQHExdWZY
knguAAdz3dB9ZIfuw6QYEkAfSPfoJ7DpC+nSilkAcvFOpoAuG131qDcM7hMp4Kap9a5Mk+6Od39u
DcrEr7J0Dqiv3z6AR6MXWvtAJ0o/+2BjIWdFadrN5U/oo41hoZftvHfOuUniM4/J5l992wYoxyHV
yT7CeVgpN5xBFYjvpoSEYyrSn0IYGu9vCkf0cWpjs0mSLjhN4zE1fby2WcAi8zUIIRATu9yyCM9S
lmb3VVEc3xszy1gQiDQNQHqdFjXYM2EXCo4LZzsDl5ocYRzrUQvT8ebQmpG5jPLWvSDtWgj35HK8
ok2vh9tomQcFe0ElbsYMctfnyuwbrmOqCNt6ei0b0fb57Ckufhhg+Sw2emlYqvcM29fe8nb1Sdna
L+A9tK8wl3cLiZap6dzaLOI2pbnUfUynRWrMB+BC/StVDuTI8qAtWOPyrOn0/4EX0y5m95PP3YGD
5Z5DuuqCOHut431kHP2m2xSayR1RSIfCwJ8qOl0Ga90naf2jQSSOxSRpl9xcGBnMZjviMWf0oC4z
hNuomxuI6oOGKk3ZKjm23KM02zI0jZchb5g3pQ+w2DZ42kfbx8kwUu/cJaMsofZcSrCtgPc7Mkje
nvkVzEv4Nb2SxlRWdZwIbC8eV5o1Z1E8MJubSQVQcWX8rqGVpx+sFZfns0QmOGZklJVIzhKXYmn6
PKrGYxcvoZ65J/6APf6StWfBw4vFO6UOwh4pV8KhaGXdnfSx8uB79cAE3k9l/NYTJ1vbxMQ/fPPl
4LIc1kxIWPoOZyMDMb2e9C4/ZZ0p3MQoeb+KAgFSmtKugZrIgUf7LKAYB5xNQLIKpPUk3rL8MKqm
nIvwUkMrf7nRy1T+e7/BjwSUfoXh57FUhL8c9awios2nomH5XVX8S7RX/c8db9O4CphJ9wIZQds7
PGpI1598+0gNEtmxBQBCdZbVepxzh4SIwyN+XGqbV1Q82YxgfzlcZu0lM5IZlhUW5bNBq4KDV/j6
TPrvb4YSBIj6Tx8r9f39wisIfaJhA1Umvli8927Q9x8BcId6tXwRSYpYTWm+rHQ9Vuofn+Pz8Eq0
rkO4U0h3Mvhvg5YeJCD7gJnaMTRwQFiYGSnDwlaBwExvY8nHdFiw0RMhL0vy7O8BzyO4iq5j9Yfq
xK8MStUdZNHkHEkxY+tEo3TNwCZUZnhkLJsaCinCDIjFGzlDJHeGvek+b4NRc30Jb1XqebIKRtRr
pEc49ZjO99VkY2LDt+ov0hCorCoWmW3J1SrOd4blS3Qqzkp0/syvonDAZZ7nEh7ZLClfMThmq3Qh
izr50e10tl9ynhiOI5kzz6JZNXtiqiq2mJ1zGpbzZPJrDOMijG4HNJ0fPjm//2mnS2qV8VSONqw9
0K4xyH42b0Zu1Dk0R4IDgVPISqf2mMwDw2Cb+ewjHdwfLcxNzZQWERAgMZXvbxI2r5P/ahX/1ct9
z/qWp1Weg4FcvlrRgDq622HZXtb1SBrRJorB/uvmSz32zaYxeliDne47n8C3r1Z5wwLwpnybxqwx
EcQmv52F49/GHOIazn8r9XOMeT/dL78iW9vkTBmpX6+LKaVOwWvUl3B3Y+vhOnceZl0kQDo3uKqJ
yzK68jL9UUb2iIdgI7dwapOKpFXEPIxsIetE3h+M6vOws3lSUiRAoBM6T8GXcnzffNEjkekNWQIw
l82pyQklm7/bBx9QrNqauhKzgse4/FqIYS7phHYQWJPue3z5a7U2zfFz7tiORuf8SB7fy0QxLyL5
tb3BNUWUo53kLASdGLtadq/HdX8HO7yQ/ZEsjkKLzpXMVtm8U0B42deDxN2itkOr5TliJvjnN70b
cIxU4c8IVlLwqx9XS0Q1YZRANkb2xyZpp4dkiQWMXuHCaiVRSoRti6gU5VOkJFrHhGGMv9acLqxC
zX06vLHk0o880ormCw2z10BK89hLCRN2oAcFk+4SgEDAFkGo2T3R3CpSQgZhGLl83f+BsWh2t7dq
nPIHo06qUjSgSXocDJj8qa7IsFWqqp+vuI0brA7e5vwpcwk+RVWMbZQ5Gal1wv52MlEwezNe1LaU
pvlYAcoidqfW4yAhk+iX8mHZb3DIMQV+6sKILXxzTe8jR0DGO/ZUwFP2kSgF/kl/NuYAg78rFjT2
1qiP+xWDylPw7PbAyvmq+RSPaCQwU19GT/XuU3gS5SDn/J8WduhbogIJR0zDnWGnFIGxji/CpKSb
EtwO3H9mFVH4HJFjGDsxEv8s33hIqXkiz93L/rATN/zkdIhHFS5nYlFuL8PUZb7VnV5KenEqv358
RwLMJtqZq3GTCuNitohE4n4p8iJ3kkBf308AlGfTWHOEu4lifoOlHtzcCYwSQnhwrwuD3PDMkXPd
ouXOPh9iTfM5O+cnQjsNdrNcOjjW56vpyAHfN7eZN3lwuHksuZoCD0KRP75LAJcj638LlakDyR8j
3VyK1Ldcuj5e9tINEWcAOgOaj2E56keur2PEIyfkBrEO95yJ+evjH5wg7FulSlAsEWa9Ykz6XasW
o8ZY1P1VFDVGP78XAFKcvSlCNmh9SFjBbekSvce34CTUz1QmOfDImtnuMCO/uoBOlVSwogGPEcsQ
BzlznU3VW41RNYOBcKxKF96cH+/lMIkr9PU82T6Fe8ejt+BHwGpQ3MKMQQacVPMIMtRXHKvwWx+I
n6e6v7IQwiJOzkUSdbEsLnk0PzYHrx1RKf78pdSSIpOTMsFa/PrLpEO4j69Kr1ISvYRBVcnonCAD
yiCZGxzbES7dEPFk9LHPhLhgv0qVEw+icHUEo8bUbb/Ne445DTqJYP10z24/uXn3qGw/CTpm6kHk
IqctvIspq5jKLxqu1oQNtrQ5pKV08cBUPn2JF+zft4MhPUf47aDzlaUo38AKopDnbiQM+8acpyvg
kmXRLx0fmpuZcgpd4JXZ82mEkncIU4AFnCFloRZCMQ/lwHV3sO510BsADW13/4mJlsHMDVLnp23j
EUSgcznnWEcYqtt8jnGzUZZXHasXq3/XOrUTL6M9p/LG/hfDsBp2dlVdGQllLIxLGRbVS6RI9sr3
Ta10vTW3fNQ26tQsb+uOfLpCnCYr9PgoHug9/X8e2lkhOzvnrR/Ji66DpxtyWxSbn/56X4Ad/kUL
BTbkPLse31RY86GI4hIWnoJwqEC2uglni4ZzP4/vhwBxQUtn6qL/D1+KWPP8Mu4XnDNxAuyYPGHW
ndRtgA0+OPMQxs+oZB53OoCsRFGXLrlmoyIePv3bwHIvg0SmyH7KVJKDtZkaGYHt5xfq1MXUxYyJ
VMu+aM/aW1f+7keYilk4qR2uIJstph8CR6EgTgFTlFGBLiXYxw/B2NCn5GwYDw63cfepgajTbOFi
9425ndHPG6L7ElR1CiKdJKYScM4vQ0U9/k2++TjwGx2RQZwB0oQBp4tZuIej5YOAdlDKRk0oC1wQ
DJvnttg6VyZbA9dO4e2nZrsAXxuscWxMsDjEvg+/QnCNtN7mYvCkX2Z/74zVeBVaty++Lb8N8mlC
KWgRkexQvV/InFvgHdn5QOuXTxNZFKxGdzP58caisDMzfZcGPnpvWYbT1mOI6F7yov9oiMdrjtqr
LujeXehuwD76YKeEb9TPPLX6PvTYWYyVBepyZjwPT0MtUQfv2/ix++Jsclz+qz2Rk+n5PHL77/FH
3iuxNGRPGSV+VMW6oNj8EzwmYBpMqGpzEAcTQiY+GxLFQjBOAgV+ky4iuDAtloSItSZamzvXFM/B
iHQT95hJWcegXDbUkJvMisQzJbE1Ktfbrz0t5D7h0V0FoPG0vy+NFQN29bxhe4GiUl7+WAXdl2sC
fZ/XsKogdfceR6XR9taBkce+fISOVWhhAGG7ie3PELCj8oVXola924E1WJ11x/Sb741c9LejkRbt
aSMYajJSYDg7C2RWoqBT4/G2F4bQqR2jsK2UpNSSmkiRAu4gceve1BW0RyOeQXtBqX3tU6LnCNNU
cObLpqiKQNOTxEuH9IsI2nd9x7aXswf+HZn0trZcGm1AkTlLOboc72zuBql2xVewLtaPLRE4mi7Y
FPoX7Ozo/2OqZSzYt5AcVnGvy/27frVHnhwrVOR1e9hnjADTzwcuM8w9ZwZnk0f3q+MSPc5WoS1W
8C9RgS4Z7uhXyLcV9Aczu+VK2yjsKSEC03/Co/V+eR/4MRpEy8ESKvRJgjteYR8rgoerB6nl1uLo
JuGLLTdttZ5ioz0L3n/HeK/sAbFkLc9/+tba5pboTXoiCefpgAveDIVIUdG5++WlwAUnV++aQtzd
Qn3Fvc/hpfSV57BuB23DCg3CPzB5lfg6BB97yZXGLBDRU1GQYfhOskrhvWalB1lgr/CZbFVboU5e
JEsf1Sy63sAMmpnc5Xt7jCi8dIKnCQAKRMJ0GK4y5ACCHHCIwnGa3lMgxnj5h5E30Qm7G1ON9iDd
GiwfryxkoFAV5Gl8PfIXyGsZk6ou9/ipV6K77LqYoOu1AMVzdTX4Er6w7WTPzPb7cwPL5fFQ5SdM
At4IfqlRnrqXfytlFUnOYIqrVOR8e3+wFtwPuDQtxVY26USKdoMkAMo2S5rBMvFwuLaffMoLqqCq
XXfa5PyiJ5LSyzbC1SpHDU0kd431iv9ZiLHh6exGcBx2uHoYKfomJ6CPBF1+ePMSi6496wty0kVV
fOHV32ceK1sEGU45y9dI3RS4jaLruWGWQiJ+Xd4LQhSau4W+ULAbFk85/BtekBrtBxGY3+1okh0k
Dp1cLpjYDqrMPvmgPPDg9u3fOX94jWFjmUoVidhELHct6abdMqHd+RuVAtYWovDtudiLbxiOKTGx
zLNUGmo/C1di/swk3ueEpgn9evmTOWiN+aTlUX4fziZRiaD+7wT3E20FthRRa0pwmkVt/XlBnR0x
pRLmICYfRNAAizkB/YQXtNrZaEiY3Wliy351cW+3iCT8clj5qnDM8nquBMI/a74MMFw73tZ3XLB9
jCPVQKqvkATxs9T0oTOKUMgNZmRu3I3aosAqyETqvq3qLFOWgtQBt46Va7rZT90FTTd1e/vwE4o+
FAGRkVEVD8Danw/9avNApIaASoGM9Mv7DiNlRQM+cY/NvtXuHgyeQSiiiU4WSye3wjQ008kVzxSJ
WZPGtFuRiwxo4qXQvoiBPGNeo4Y5V5p+XHBCo9rpsl/bk8qKIoMqybxy/VDGZovfifod6uzldosB
HNfob1wGPwSTbgBtQe8RMe7j6U3DW5nJ5crrnr2qFqRo5X2Q3+2r1L/5JlbK29Y+9zf5+ERuus3y
xYqWKJ9wVl+lWdRg4ZvUfKvYKeANIy/UeL+gmTdd2yk8KewFG2YKFiUO4n6HnJi2EfT0ADj8yWoq
EpZBObYVRf8+Pop5kuhzjtIznci6PTFIfy9+LzQ6hC7iBd/tqobY9OYrNCbzHQnbcAUHvucsUjA0
RkNO46JDOFMgtrUENMfWYln4I9bfPpnauKs7pcDVSqcZ+dJ19nFcUyR7FJLzcfx8PtjkBC8RGFGs
JCyQXxahNaitwpLlXWrVdRCEnlda7ch3c1vqjN0KdUS3qe1GofH/gCYzqJHHpb9mJzPYofFMlelZ
BPc3qgK4L1wNwTEA4pUQj2ER5SKKcLOp9mLOAJi0K90W59vgYvb1NjMWjqG5v16I5rttyOe+6oSt
yUA1bFYhIK7MaR9sslCsKKzTtnunMbX/A4bJlTMzwpTh50eLZ15yBhPrRJQ4esbNCigfhzc9ccAF
7I1XIZE60NE3/DF5FXwAas8OnQWPskKPSPIn9nN2nzusgoL/6dyMrjIrUlxF2YHZwAv+7XOOppBv
XO2JF/2PCeP3Ko7oWmYinODFldNGtyNAnmp89236UmCu/NlB7UtPRk0nycW1dC2PEI7f4/i9OG/7
ALnp96ha5ZuB5BCDbsIbWeVSmDV5hTyFCJO51uOkMBNbD9DOB09wSCXUp9chO3zZI7M0gvSyDc3M
16pfXN9DUb7XuC6ZrSxRVa+xWBWt3hjM771WBa3IdfwJ5iAadSjfoxl4q9HuRE4xeLwSNxK1mBur
5M+3vYnHYt6dHBYl2dQ5A6fwuW/N8ZXvwYBrv/8yoCRHOp4YrxnudBDvheI/0b9fJ7m6PGLFw5az
EiT2CHJU7AjGSFS0/q7aT5WMbk4zgmQGvwRSYKQFq1/wrMp8N6FS5PEUtvMdw6oy9o7jXJKKiCYS
vkE7gCK6Az9fRhPKtQLYASWh4YeX4UgOIRxJ7cHhPzK6jlpytuG3DumU7WswIgfMkzF5o7dV2fMY
Dp6UMRCN1/8CLqYjzzFsLr9CMRfLtATVTsnPCc425kzbEavewfQx3cssVAGpaKHBXY53kr+zUAQ4
H8pisGJkqh/2037Ura85V6tRFjq2SacfgyL3tm7L8HAZg6wEQg1qxXjavJu49ezGp70e9hgpQJht
Fw+UQk0PoGdDlOR+QiqLSsrs3wTX2yQdLnj+3YncPMjm7ln/7p8CyBtAvA4Qm/EpArn/lSGZpYEm
dp+vQ9WDbKHg157vvxs3NZrlOnCroxaFnPWFFCODMj4jwjSoQrDzDLZDHxxPPxnglmZLA8FAQtc/
mKInB/Vk40kN+IW6KMAwpL/n2Sw8sxJJAskwQVmImVFhcKv2dRG/N2//lFswh/MJjVMrCJRbJrVd
t866s63rJ8tJgSHRpKVB9HERLAf3RcrvvPglxFJRqcWPetbi+55MpV+VOt8Elk6n4irI1BTxYeQJ
xQWQLPguE58OfcaL81UNCKJlE47mbsXEJV4bPzvGR6gw1uCZbEYzdlUTwAK0fO5fZccCNCuK5FGm
K38pQ5j8jlJWxmcjQqoeNLToDqE6JGMmHttnXsrLmGA9Be2IL8i3p94OCnLjTzzx0xiLwRO2186H
hEcLzRl1RsaDJYFrcpLzTWxp7vTfUcIGmpuaIB+3UCd45jakm2TTFgtkwO7O6eg7EwCcQE85TXq/
gHm0wyE0bD804I68s885WNeHdKhT/+2dswBVlS2KJ2bYzI/AJKRRw5QMoFIwnKFastOb7dRiyEJR
hF/Q9mTabODscjZv3zi5GONpZqzEZHlsTTptOGHp8mk3hHGVYow1rdRwLjVF+DaBXRnDbJtMpRib
3e1FVhdqOLO9wp1ekyQR1gC8r1vbxKfHo2s+CqLvcAnOp5XByYkGTgl7KLAVwfkqtwkaNIa+9P8q
wmiMBo1I4xTx0VVeLH7lxOL5Uo6MREYZJ3Lx5qSdOy8ws8HHvgBCjx1XMXDWJ0KMY05ZprfcXFz/
Lfir80UsT5wwJwmPr1HFZlvqWdsCnUJT5beToV/4EycXCPnwWw26p3vV4p6XPKw/iBEF5aY2QsNr
ujwB1fdZUpwTv/Z05VwGfWo7oPaCXUtVqtKYVnjIbDmOfpf4j/ahjX+cd6g0K6nwCnzb20ywyJrB
G08ddg1hAs2kGAZ+dZzW2CujgccfJUBS3mrC8HVdMiDp7sNh1oAgXE+pD6oEsWniKFbQLPFdGeJI
p/ws9/3gDgErGqS5S+zdueKNdRa0ZljiA56GlHqKpsj8PECAwkH26JRGf58FU5ZlwY/zfcrJCMOw
f5EfCe4ijcoVgiaro78qsAQI8HcYLYZQP8XsziHyZHTrfxTK3E6bdtWUXzXHYfxEhVswzMb8LR9/
HHVhxu4HlCW/O/y0ZEAJDsyX4hoMmvNhzVrgLrFknhA9D/6u/KefNAUYmmrQboBQCIdTTBxR+fnl
HMlcE+HLU36SaO+yHjiMEnQdaeJVlhLUmpRkdSqZjzRHJaomTp4CCEs8XA21MJK/zDdOwd3ORZtw
U91wqPmD9Vtr/9RAudX6QiWRSGF7Zn/7BCLrEighZkYdvmbQ6t9jwnmk5MpxRItJS9e1fZpuZHKx
iGvAWYXKG0DDojKiQC8fBIail6xSEBsr17Uwhe0cId5XzHkqR6omj7m5j7IR2YZ/vXRd/F5n/y0P
t5J1RkKFtE5suY2SeS30LVOMYH5uoYc3Vts+UctPwjd/2yLXbKj6YhteSZ5nMn0lwFVmE+FTbijX
S35M7RC/Lid9ikPYddxmSECKNa8ltnmluc3Jwv2NRGNE/v77QPDsJpSQwG+6HHlj+C8T4IcvMpZz
UraasLt0b55ouUMrMC6bDKFdAOw8Wb1PRB1XXjNIMBnVFTPAvbBJK5bTl1U+dPgUy7vvhdyrCiLG
9UisaSR4jxcHfyszsl/Gy3BBb1ZNhXXBUuzisxOVZvDUVsh6soP5uklhzTu1I1uRVU7CEYh43CWq
Sfj/c0VakQjbOFH5HukyMlI725ceG1Sc24hTlZRlNwomM7sbji44kLa38zrh7/fCWQxS1BVq7qpF
t1o2GP0WWtBDAySMBuhtCVoQKB5hSIyMfSt6FDfUMv82EPb/A8V/RcNC5gU9FrxgW/JGyzcnafnO
cUGR5LycWyeHlm3//FrNGUQd0sVINX6GOhaOs6g6to9zAD0NlG3DE+rmKeua1vuGMemtOHivlRCA
4IoOGhGMnSNekOjiJ+nGX6YFQZmpQv9KPSEnpJAZDHi1/667r6tKFxrDCiLyoNd3zVOOaRFiCqu9
2ElMdLKE0lJTlMB7IfjPR2izvQ4IUauM97KKNtMca/IQPts1eyltJVlivKbm/1DOM+WMJwhvoyjS
QJDTLnMlKA+8jxaDGgHd2KuRuEq0btiPqY8PJ+hHmDxhKvJLpF/cHhEz8pMLWC+K/HWFcM9mhA3m
j+0/Xvn4r2T0RtJrAx+OtIurciNmxmaiHIXGCeof0WDgf6B0k0qy2Fdz4X/AW2UUxoXwnzMzXVDw
ighJ5SzqeBuzPNW9EcfCeuFHNXyWyXgSTkeCfKvYsWXXK5gAJl95kGuzCVOwZVUl/kRSkYirgrOd
1hJ0BP6CDIwxNqmDh8Z/4FDhs0iM7Q0jzsrxCAIapYO3U9X61VDplMfMIZhp5up+AhexuKVRWudW
p+lre1x1WKnal3hVi48n3yH42fEWUIwLTi97AOQbl0NF13PFC16DYPBhYs/bEyC5D5M2FeAa6l1E
E47OxFEdPNVKBzaS5s40jlFS6AZ7Ra0mJAiqDwcsHpQd5B5/cyDEi/V4Q+/hhaadMdM1txy/54TN
OzwU7Jz6ySBvVrzvUjcHJgQnu8a2cGe2kEJzxYQX/WF3Tgdj5FNL4t1jmutcETDZrE/gUXkmI49j
GJYd7B1QjF8rSgLw190KY6asL6QVDvL7I1dsDAZ6WrYhH4q7KQR0MvSm/je/lb8D/QfnMKVcuEig
pY9nrHXcKrqMpFgZFGSgkLncxzt0ARPi1AODLc8c5stSX3A8BmJc/pCqcxdt+CtQwS14rV4NiovP
VI2db4LCZMntLTXmO3VBHEMvY4K4MUPjKaQUKrGAXPtWDZM5SnRQ4jS2Q9ASn1Rr862tcI6A78Rc
y8IHoBVkI5TqjHHiAKV6oELBc4Y9dKZH6hiCTr+JmNmTAFq0EpO1pd69EGitCkBjdRalV7NBgudf
S2p0i81GX8rK9tmewyGx0+8Mjb2Poj3Rv5lrbWzLR4EszwsCuISQUdRbPCgBY41Emrxi8yxPiN8b
DHvVzShyTgvvVfVidocTCO2JJYGRXj6DuNm+5nKhXYYObrCggKP32Uv/FL+csyhx7EQF1C5xqCVs
rwqQifGZH7UVKMJPFNrrldzSXoyAOiX8NyiPMFDeIA2EQc86ngDw0QoZJ6xadzWaGJm2t56DCT6G
lL6gR//mHgMMKgygHehkz/XyRrknRQ1DqS1Zri54Y8olNOXuSbsZRePXPLe8U8e/GdYqDdcErTa8
pK5bPRDDh3UfFTs+qr/ZhOnd/lPMiuYgyM743LVUa4qnNP9pem96cwp7TYAJkaULmR+ftYf5uzaY
HEK+DCPDIu3YKTqrU4JsnqrEBTdMljiBWLuf1iGvHXrCk+xqgFiZHchZOU4/0sfOdRVmw3KpZin5
83BrIt89rwf+aZS/Z1NLWhfdvVF7JmwLpCm0VMl4sgRqYlBdVr8PPWFqEIYyzv2YenY1sYjmZSGc
1zJr/rOothq8IVc+MCJJgLeCwROdzETHMaauxegt5DrD8haQi1/LLE/g3nLFlSU4hDdDYcUTS6FO
PcrO0C4h/7be9As4S1bY7rht1/QBdLj6yCC3XLOc5URwbrj80vJ8fUSosg+a5SAvlIO4H4cZ4hk5
DI8KlciSV3rIQrImburlGHhjetEfuZ7r69GDC3dILK9E1PuZTrfz68Ng6DwYYq1f5ufCMryxWHkb
MenuP5cjKq+SZFXxvF6Vb33ZmKiMY2MeMQFcJzFvdnuHSy6rXO7wxAj0peTwlw3rAUOlfsXHsrCq
VcOiD7PAbyoQTrLgydfKbFLZrdg1FXPfTKAAJI0GBiz4h4IG5nU91XzHFAFxcGZBunaQ47an4ShA
bL/GsUPBN9dN1XuVJXkRz7HwfHNdFBGF42k6g7oPgKWLSqJLXnLE9J4S0L+NSV3+ocuVkk2GQQ7s
Fs05hfR56r7Mf2Gcj8j7JgCGyDZm8zLoy1d/mxzBJ1vVvIul8bd4qp6jNJ3X3R2WALER8jvWlMlR
5m8jT7yjDdcdq1C41E8vr+SX9LThpQK1eljMg1FsKVj6JMznQa0bAS4YUN7md/mgf4LvRmkRawRd
zOYx9GkBX5vrmS0XgT8LaWaHT++eTfEZEn+ld9nLJAV7WPaxS0lo4noW3f/Q4De8DUQ2P4Neavz3
w/35o3J5KJPAnnhm+jscm6NQXgX+BMuxoeNAaHE4tXJMr6XoI/Ok9v3Hl68QRAJtOen+krvL1PZw
oys6CxxjTIr+CSL4Hb6zw6aTe20W6ynPvbeCcCRfJzoGnC6fj5+Az/sFsl4BF2wh5vDdiCHc2HQz
GUP99eL7ZxzmAuOQOC0Cbdao2wd0ovhVVnSHUISPQvBh1Wj6Ruxl7ifB4BVb4DcDT/lSgvRp+HeQ
WsSZNYoavFU+udCXNeh0f6wa8Kced73rXZJ1TFSFHoOyCzF87n8E0ehlxHJEeIE5sjnQ2GNdyGrK
BCLH/lGL97jDXZg4pem9RXgLhftCTJRinvyeJeQWSJep6wJO39hFz5WaVyoIKm1GwhS7wInDT8d5
i+YMf6lrNVHVmPmwN+MHvnb36EqRlbIebFYHWrwREhEwmyB7VHzg1fHujjXITlRNIZSRSMo1dhsU
YL//TEo35g5l1W4cBK1kFb0cSwIF6atgsd7OsSJd/zaIYlY31HYebGeyIvKkB4NglKlU+y14e6uX
CSdXUX66s2wrT2Sl+a+Wio6DDwvzIG24EvIjS0KPExNX+09Hneau33Y02klHi4TSji+z0zIOLVLG
G7tE5X1+7kHrGGWQOynsFbEVDQKhx5biG6Rv/tMf9GuMOR3ANz1rrmcPyWO/igqT9YowfuDJWTtx
4Kd8gG/t2iv4EAVSfA2TsuVsiR1Cai2YVUb95Cqbrw9FuSE4PktKjG+tGTr3t3oYO3nRVnhSw3fK
kftwJCWiJy/Eyc4ZuQaFhziyXDgcI0xe2U6AJji69GW0GojVWIaIOJN+PQAu/xQiW5IxacTmJc8v
MzwyZoYiXnfvTvLdiHcvWinGyC0L0p1Zo9W/FrtbP06+UVgJj7ApmOEZFHxJyZ7/SAIXPhrC1SmQ
HQhpdRcgYY+CYVIHodZ6euTvoQck9YlQmlMUiVkTyTXlEb/jl8g/oVe/s9TEWP9ZXLbSblzZVXUF
IXR/lxmdBt1g1ih44W3n7nSI86jrElFesOAgJzK0+5cUISdZfPt+7xkHWsD5sgIHMM8Ejz1ZMOSF
BnnBoaEFoyqDB7Yq4zqm0FJSriYWTKseBQyZXDQUUD4dBFE3jCQt9S46FQa6wI9Alu+CNlbSBIgz
bRuTbC3wpUXcbX+/pmmmjkTzbYw2FeR2hKPDqfweogwMtreJINdIth48XAfpRS9uErDOA7lKObEi
SnLArkTkeCiQkV6k3RHyOVQBHn25f2bo1pKfqqf3w7jC0qmUg8fIUFMvqmhNg61c9KIGDfP+BMQP
wC3bgpjwy7juFFvT8KgwTG35ji5RWFXIz1/YD9oxsQUUXt86NWELybHYJTjpHGVzaGd0MUNB1M78
iLbB3IrDOkzhDINmRBESq6h0KN9hMHJxJVKzokFINRFRKbYrBdecfkAHPff1xdA2Y6cqOM/6MXV6
3swvjxTLp+k07CWsnvAZ0Kd58RQoAemluKkO9zqg8sTeCXxDqNPsCSxNTPGMmdqVUsbJXYgFeaJY
wIk+8+tiaIKNhpYZgorGj4nXZLVKgQSyDISEVxVmsgUnac/McQkrfce3QjMNbwLAXD8dRX+h6GwG
y210Vu4AZ72hj0qp4AmgTpkRzMkcSJQ6NrweUE/dtKQbMigQ+p1Q7cQYWEJG5zVO1eeHUGIWHEOa
yl2mQo7FxEaDg8b7bppyDtNEwUG8BMscSIq2nBuAG6sneuL0J3I5xXzYGgyaa3QyHwGeuv27asHW
7irVpDipxLYFdMRbNH1nQfb6Qrzn/vkuCqY5jFudGApLqRWYT0qsJ0UHSzP8Y0Kmz3j20BXesU63
cx4AbJYwNDzvqNoas8ft2U5ONPPsPi32dpjx3tj+RVLwVz2k2zOoGIDbFhuo2ffxmpQDvmR0mXzS
C5NboX/1vth0NLHOAWWOOGiJSKKteCkYes5PcrG+IqJ0xDQXhkiqquxGYmYUKafSVgBSrg7OV7cU
vQccXWBguUmyIh08t4WcUcFbq6iJaFkk7bbNJD3jH1Mbh8AOJmBXB4nAbGkKnH6PIsfH4ivTKaBp
yIAhHiCzHc6uA0MwQkzLhQBoxEiytEs2q/an8iG2Mb3Igxd2nvDWQ2YuY42vWVx2MB1S9D38YOFf
LVR+SqtCDAg2xYKpAkt8HHc5QTeOJMcWY7+ECyB8PIidqd2KD4gmBHNXG2ofvzzwcFzwJLq6gjLx
If/Mdp6rRxJKoqNvCXjz3NavVnw+3wnsJGDY7SDlD+mmrJA/EHZb778e/Tdn5JkeFqJaabW3Umhs
LDJWntSh1tgn4zXoNisM1Ql2Y8a+b/hD6YT5azFzeUnlp2MyfIJg5mxW2r/Ec4sd4/GKw2YjjAlW
/L0ZNK3L3uEb0AwOc3Jn7hKkh7dxurFFJs3VLLmI4YhGstJrI8E/elRP6vw91fmmO0GL7qO63byz
qLUKnEuBNLz+OiRzYXVTp3G5wCYn/d33FTJKKMiTkp8xl2Rkx686hg0qky4CIsmhUsW4q0vqjXq6
7tPNqWaTh2RLAjPzL5yKzUKoeBnjSv22vFyGTgTj+sQkGZ03Y/TJCpjw0ij056q1zRMMOZVhJub5
vyhcLeWzNwedpXwHVmW47tcY07m4nxccOTdpmnLO/xQG9IIGFNvhTP5lpUzMRB2sr3kOl8zHJ3cq
Q9hFganLi0XC+yE5D5fmRQKxkr1fV5d7dzH+Ma4YYNwwOybg8HAiEdkNzk7TzwQcQz7JYgO6exeq
g0Geq5RR7F0zPXHs2r+FLbwd7iaSl36DBp92ljGFQj03ApSSoUt2laBFJZkFUPnrrrJRSChglJvb
a0rTfxmRHGCLNbvZ4mF4crk2h88eYFlzBF1G3zeBcbzn1MXmMxaz41nzmRPCf298fBWVDGnULKye
4dFRkBliMXsQU3bRwUo06r8wNIPjLP2AyeNB7zqtDLETjK8fo1GxElnSITzU4HwvMNZodcfNV7Bv
CJqob6zcz8dx1K8thUx0jM+tI8R/MfPkz/Q0Wxgy0DiLzAd2QBJr3utFSxsCgWhreCYfegSVvV1H
Ru6muF2CEay4oQ093GMhr/SztjP8dl12HYycdZUmoqLXpM++bDJd6P66CnaoTt67I+pQfNzKwWHg
9cLQYQU/ca8eJ0EGduGOZ+uCeO7DOhUPgLQCyzoYUob8dRwtDB9sa0UktBAeMWaLm+TSTu0zi+de
bu6k9pr19k2DTTQ/Dx6q8szs5X+Xe2cWCdJ0tzc8XHeoXD/+shqrb3vNdX3cd/I/pzJLO/OOA01m
oF//vP70XbNR/b1UtOLgUCosqnaW4E76c4hfoyI68wEfZ8MqyBf+7JcB7Cg3lhTyNutaa3VjFfqo
HGYeZYoGl/hWhpd0s4NVWeTYChvvyhO6iW0zCPaX/L1ABM0sHYmFxrr0msk/slOK+n388vw3SWdK
xXJSL0d8D80EpEJTRu1J70HvjzRmx3vK6zcp9sm0QhqACHhuOIQo7wsGktUbUhtfDGTITB2SBUUf
4v1veQ8JotCdmZ1rxDsfjW35bzLDjY9o5SfKZAP32CVQp7cHjrdfcRYjB3VjR+zLFlxLLWhc+PoD
nWsUbQETdJzb6AY7oczLPRnVGkj2z3xtgZ5ez8nV4ivO4sg7ymQZ1zNQPFelu0e38DUYngdhuZ1k
9UuxnI2bb280LvfWBfg8sVKh4Tcj+T4G122q6pg3i5owhOhOUqylpBEsRIQlol1OHuUMeqJZAuE5
KTlvH7LdubnIDxu2KjVKIopTQncIVYpKrjJ2N2BmFwEo1/F7TqWDjuaL+37GT0m4ksvkA25QJ0Pm
S+/7UKtwKE0LR1HjNfUs6G4ZY9g7uRxVByI8ILZZ04QONovdykd4K1a6MKtnPXXG9pyaAQfMOM5g
uRZrTKa8zMd/izPe6zapNQXdT6S6APgvtk+t+aHGNSxXT5xDwTW9cSwzu6sXIjiph5DQ6SkBcMNy
qWukpoXjW245omjUFxQ05LAdTduow5WDCvFkMIKl333dNaLlBTItgSbvJX+SQXZPopJU7jRDutvR
N4WN0os5ShbFXZb30ihgs37q+MmsBxzbKQEuH3GFJjyt8chhXKcYf0UVC6lK9Tw9vKXtgVfCRIT7
cX3WRRGcgfwtV4Hg0FKiBuBfD+h4yc8zYR0CHsfcAt3Jj827KoLhjk1NNg9dhlx/F/JdwmDlWeOO
13g/NHi9AXBWHBpLbiXy24unEk6YkFuXpUOBA9wyxoNcQn5H+tVYqvCMAAIX1TzNi/OcGpZpwdbh
00hCbknTNWTbtJ/kWpAViSL0Jxlar79prlCB/xQ5wS3F2fP4xA3YEguCleI4xZWS/1FnjyjAI8sI
HRuBTtQS+/zNVAim+PIuWtNiuRbsfclZFluKZyj0wYw9kaR7WVaImO/Wqk/Af8SWCPHAISQGUSov
Q+cDSRFPuIC1/9DCM9WaHuJr1/JfrqiTNgXCvmtYAQASB1Bj7ewFdzM/S/PyRwmN0EOVPFL7nPH/
1+IrnHdHfHidcbsWNv+PLryYyEP/i2wsrarPtp5zQHSxS5j0I6hzyggD5RoPGsohiWPHB/HmbzXR
ZJPhiy2ALE5S79tR03wAWvuW7gEHlccrOnJoJNvF5O8rlYFk2Xs+CMrgEBPdIUt1feRzQdRXrzWu
yV23THHTGvlGnebIE4CWBhRAs7S5JgPCtCY1dmR3HxRKwwLORIPC58w1YKpPfdvXdore3c09MuVo
1x1zG5t3SrXtXRrzPYx9w6MUb61OydQiyJycQ5Ae6/SIe8AhWbSOCbiNkQWG4bcV8+dgfQQ01dzO
awxrsIPW5dMdd+aJHW4GIdgicnbx13krFZMBWSGqFcZFj6GhBzLbVRDp47/i1qjX5kH22mNu29Ej
/J5a+sxFB9LVmvi0WrHqL5g5gzojwa8TL0Mr+dVUHTdNucJ0QeByONOdT4c9e8fDhLtHFHcb0yRp
HKYTUbnD4b0yXtStcQ1tNPLHHI32AMNWTtCgkGaEv0WQ7kvNbWpwYaXwLrTKf67Sjfm4abNIo+61
QnZtHzDu9n/gA8deyytPZ/E6bwAv8Bpo+wAb56rsqyvhNeEFZfmmFT1F4VEqf5FeYI6KzJE7wTDv
M2qGEsW2k+D3vAaAA08pp+sfB14gQt3iPGwdJkmi67J/sK35q/F1JjFu+cLGbK3ZG6zG0w+sfQjs
/Ii2ejjFcN/34ejnDBWYTDYUriWE+n8EwrhHoylPhX2vEm96KxPPUpnlnUnb0HPCV4WAfCOhpini
zIOSoGsIY6Y+D8zJhusWQ+dZYaB7UUDPS5cUWr9EMcJNkTqJlgUI1r+sBd+KcM3CA5zGUoX1VxZ7
OzX7QXmJlJt5m/Vqw8Y/iKARPGlkeTrBTOHIMguCcVmG76VBnl8hlVl1KF9ll5jXDvjsRSuBDWbZ
zMiXpTBPwUcZYjXBuW3BabGoxqZUh+Jw/c1uazrsCOy86EYy8FFL2eu0m7w4TX51U5az2vYmNQyx
KoX83el+Zuc/wD55fBsazwCEEdx/RjeTUU4KJLoHxVSMxsoOYJ1YjlpSezkBpZHzR4Ud6O5twn1B
Lt2OuaODSQc4YVdf16/Ghhlf5N8UPp4eXyrpydjGs9qDO0ARRt5PLOiayfkwVgBJQgW1R5CrB6hA
r8rNIkm6DaXN1ZsiD4tGM+n0WF2OFpVopQJX1vGKvJ7TJyjeX2Do4H/X1HNhAZt0S/hl/uuzOeDO
ALWkz2EqObfZLeYoOHvcmixPaR/Q4/M9Q1wNONde+QnywsYBIqAY0NTpxKFwsVA8RODoXBNLiEe5
ZvQfbPs/a/Nldm4Qrp6GbVn7x8VA6HOp23ubDtrNh2D2KePnCGM5b3uVU3DACElYfwCjwQThAX9a
n423N06jQtIIO93/IX/YfZyu4MqvD5q7y0+HbWUMd7TXRaZihB/26uPo4KFZFQGyMWPJ2if7hG3i
DOjv3qrb/68EKtaelm7VYX1WZy2T2idoVgp0iCgz4Tp64/zCw4exKr44jWAiX++wdHo+Bh7I7kbw
dLhesf4h9cBtl+vBMiAXFuoNf4I9PV8f0VqpqpnmyIzxEUPoAz3ygNaJcjYFnFwmt7QwhIbtMR+U
5SaEExGrRrhvoawzL9OMrvXZqqmN656V6WT7/vcXaWCpwL5+VsRwpf/HulBATPkkmGyTQZOrIEY7
+T0Q3EPrEmczsRpmFvwoPzCrdyyjUPTBKbRv8k0QNukT6taQ2DMeIK+falksI6sAavtMdVgnBTQX
j/x/Z0YLOOGy4SrqbG7b2TRXFJnR5LAywPb/LtPswO9SpLpKP1jBGO3TpwWl/PUZ/SDmidHOPf+M
eNxXMOEP3M/36jxz3yiZJ52itE5B13PfXb2X8g1S8ofzPBnF3zg+JpkCoFi6cg9MzVrRBHjZqraq
3yJgMJNR7fKOxlZ6vgZcG9155ZQPe5XO2W/Gnia6qKnlA5SImJWkXuqnwuwMxxnpP5NsczNf5Ai6
/unYoWJ0iQ4tIHQjLy/Yy7CVxb4HT0PStkdfsHxxjtz0QEPhN3Aba+SJIsUN/nBi1zWHUJHv8EP7
RlQsgwVYE2sR7xGmjEuCzotyHzK11zmTBJsNvMPYqJs3+wjOkA6n6E9gwfreDjrfkq/+OV31uQyo
w1kf7vxigGjn6ZIQZjCZdmciQBn6LCr+xQV/DmtC4DqB+cM77sm+BhjudaarlYFUuOCUaPgz87n+
LYFsGTS2exAWkKWj4GewmrEhw7b/F6nqdIGzXFIYAa+JzsEXsnzjZregxW/gplWZ4XNwcqFVGoFY
fTcpyHRBL5vsfd5RSiFi/qbIvYLUoPWelGpobYXXUPHhIG4Ib0pW6dp5KZ3LvDQSnl5yJMF2MM5+
hIlOTNnEK5CxPnLm4RWSf4q1lAwUdK+CLS6VvHqwGVa4FbP8JuFUqjTxDasA4dMEc8xughxVLX2X
BgNSUAlbu+cz1pdKkS8VM/LJzD5HyKOptFQQZmFev+Fgzt+JHniXoyW5lhNCCr2e5ur+SI6QkWN6
MF+GRRmbEZGQPBmjsxInSx8ufXSIxegH6/UiWglqCF2GSkt4WAVO7rDTGyaxz2eDWYWSAWjM5IpW
7xWofE8fiZyC9SSjGNOAnnoZHQxU9eF0G76n4xn+MIEm+BW0Q1i50xdonqZlsr6Nd6seP9+Pd9tl
4/lmQEZBhKuKgSQaHP83rKxlkJ0jARbTVJeaeO0RxqiusXSLIr0D8kiqlWdQ/0GZHQ8rmM6g7GPa
dB5yg45rRIwGZPyR55gofwfXeUsWZOC1c4mTqY1zGcSW7QUVn1PmXfu2w1Y3Undxpg4dddOgh5hH
p5sCCydZTSzSphIByJp/lAwbzuwOSL3kI8TrMyhSVCAH6RTFNIa+2MHxLRpSQK9FiJw10CCqzqYo
bekD3k6eQ+vDBGd1TwG1+HQ1IVyl/qNs2ryQrNK28tV84wMQVJbtMGbA+qNT7/L7KQUvtjX/IBNA
axP9e1Zrwb+E1c2TPLU2/ZMBpkOonWGLswKVMkLsUtpeN4GL2MmWvxi+meAvs2W5FTEqfOf/8CfK
IyablJLCjRsiaauuDMkYNXFpi4aehKu8HPXlDStoanDdELatRy6b8K6aDOB5FYO23h4NUR4b0eDV
JCcZdMXVgg53fWPz1diDhgtPRSJPWlwi+PGQn0dfAyKS7Vqrwbh6XT8Wf0D7wwRdd2Hd5jsJbUf8
nrHGgPstONEcEwvyZCNa0vn88NQQCtXRtOEn+6r3ecqcqe0FpO+LD3BDDoAiGisb/AbVljMyqhTC
3efShQD+1rPMl4dnwIszfNQybaORZkCele84kMdOpGeClUDf9RJGPWqSJ/W9wF2j3jALiUnut93k
qHLhPpp9Ku/tBMRWksJ8hzwufcL88JPAGTQ7Szb+YoNLx+8MBr0yG90prYUzI8EMpk1WAjVIrC78
CxLqlVrRSIVLB0nVbOfjbBHgpcb1rc8qNOSgxvi+d/LNA9mRjJXzJ/fD7N/oKAMmN+nN52xePihs
EPJnYLN3TiAHI1oRtU301IO+Ninu2gY2uV+WNbUTthTLhpjneimfK6H/9OGiuagK7g7tUbC7qx9E
fcg9MJ1rzgeslMA24GifQC51XDZMxAbFrG5WuY5ejjKy1uPJJkAZlVDND+1v7Z+tpzrkh23LYHQd
nJQkVHR1yowlIpTxfBXGznade1pt8wE5DU+md8uAagfxd1dgUVTxuL3ODVUQOnS2pTXMPDCDfqMg
JtXVYpS6oXAv10mq5Wz2LrkP7v/9l9+anDR6IGNyOTibFNRRbfBpfv43+sLzi8u5bniFasmc4kRB
B4Mr1K6B/F17h9m+dD/iIC4Jv1DKm1ZU19nu1Y84KmnNo1kFVJGug/ggGKLgS8DG7SB+t1W9feOo
4/2JXr0WoX3XXyjKRFvPwgZXFyHUeUvXimPmTSbnYCqyGqpgUzXeVh22IAizcoraI/xDVybzcDIA
uKSV0lqAWYQ8hb+OB0mjT9d0Cqohzn9+WcHuQpLRZ/7MWq4VX1p1otYj142Pw0DcKuZlPS3nvxem
0H2ksWJRGImTS0o3OOwbzsFuzH6W72tXfttL9bbx6xTiUDeYU7YHOjwDb+u9tAt09hwYySww6BwD
AcUDQGuz/XKT7mIRY59kI/Q9I2VXMbMKBmRS+Yesn8nXchcXovEgBkp0kDER7kPw9BcrOMthNVgu
I1Gt6s01C/I4kRRsDhfhCv8mjcfMmJu+w8lIWKLpKcMCQ/+6TxkFz9YDgtUpYMFcwDkb+NUtRg9y
5x589dFPwE0d9Lq76w58Kfap1uojEVvBBR/fVt8x2Z6zecSaDxGQzijmZskXjPuQTMl97ZMBxWU+
7kBrrQNy3D6cOKvEBqy5XNgvwJbiUMGv2vBZ2pbZmJCEGaVZAIBdu3oH9Cu+0rHFZMPXIQmkQTsu
kuVpiCJcLWnHBCSWc16H8k0QzqRwG5y4xBXkJ9JfK0ip7LVKCww0t+Df1UI2puQ3dbE+ASJBGXRd
C5eGhw2/3Pn1eI05kS0UenDZdohs7HACTdy2WHnFJelT5T3sWSY2xMkGFgkw1J+ntQip98dDNWOc
8ajQ3rSh2DL4Umu+u+0GzY0IZzGWyRV/TfEXwkIiA9ZWEXAcRjQHG6CHP5Ado1CS/I9TcIqHN3qd
JU6sLy8x/bjsz1VIqiO49VNUsBDyooSbPg1QDL1ZRsX+D0xLQkJGhRnXzNCaVf5q3RWA7jIg6CVk
hteL+cmw1WAnGNo16ePxKGmtbKRe9HevNpNYk3quKUK/zK/NkgySIMgwOgTGC3iDr3tAn/S5pMNi
SQZSpJ/4/rBPzVg2MtqpToCvTRCIlyhlNnjfexV/gijmhd5w6wH3xI/kAR9F9+f4oERFiwKnG3Gn
5OQmbuH+gbVxzm45pKJWCdBVFVSgbH37RBF4qVzVusyuxhOJGbxqZbJM/eZQ6njmyyOs7ukjwSeM
ohGrgwUL3X+OEnEhLVUkp9TAROJpteIqXM0H9YFSwsCCiCqyxnyhEzXxz629Wd3sAjBwIn3FheSt
cPavtAj41KGtO9s2nHtiAZZ2ZuWbgjZkCzs+mwhTDiTAI7uhhmL+MWEuDf7J5Zt6vNMKV6ehaYsE
WtDuk5EL6ZHNRDWaI0/rbaOIvyumAH/zioGEz/v2lFI3adSQ4aNVYC1vrQHs1s9SK8HfVJNiYMig
aoWkCJWQK7PBswUj73BZXT8k4TMBFij1UBYstyjnMrU9GPi9G4heRRzX3wuZgcbfZBcQX3t5LgW4
etbk3ExENp7i3W1J3CEg1rnq81lLWakZ9Pq0+1yJuc/wsHMICR5y5TW320lKxVMc5qAAzVbjO0pE
/yLrJhkBXpz2TzkG2VuwXsGGeYS6+FMS4q3nqJjN8uTrQAtmef6qTeI8nShJ08DzhwZUq3Ykydjn
b88yR3z/60DmzpuCQjC15WVaI6325NgnNW5NRBWmBqi9/y3Rbq4QfcTZ1oMp6TXeUv4YoBmA1Y/g
Nvesbz//huRiCcg/X4FS8GbWgLVaZLOtZRtdgHA4F4brbbH1vCJn0SUfrjfEtE1776wh/Tf5fy55
2tAn5KoBUDmDqkYY/L/24Hm379vCGD+lnvrj0k3TPJVjqggCiM7nyaT7hZFFeQb7HstH3MqWimQw
g6zbGGk3SyBDa2Ud9HeZ84RZURVchkl510bku+MaBKY37ew1fArDIcR0GmTx0Qz/2bm5x93QuEIT
5auFmITy0KQ0sh8HlhcxS0sM1D37EKyqzitCvFyFsDruaMk9kspLuPn0LxF4JJ3wCfNDI0NqcDik
hz5EY7qcdL+iggh2IdOJ9cR68//qZJhgZ3onKqukWhUz5kYQMHcEBbcJTQxjeAsiblCWDyBirJg+
xNVNMWUNVAouaQPw+NusHUd5A9VapF0wqpDH4cgdizjq28CdP+zywdzNsUstW/l2SWe57IMOc5xR
u9k77ZbW4Gc/tpuMT3VRZSm9fZ9tdPp4wIVL5JXt1cUyOyqa6lnSlv62eb4DirgpoeqVatQ5ynaq
4sX+P6rkz+5vhDSFBqEOyCPIECGbeUGYN1fKWau/snyThgjCWQ72OGYtmY87k4wYWPO1PRCRg3/9
fNSHWwak/aTYggsjWHbk6byteByTzD9Mh82u99OSA0vpRA7Qttmi88Py1uBlkeHbC0qMBKrgBCm9
yHXWzmPhrNVcvePWqP1SrW1dhiKJS0PTmOXw70xnzmX9s3qwpKEwItOe0MUqvGDQB0fm4ikPYcoQ
G9jDIkocDu3yCoLuVdP1DL/Fd1xByPm45dSP7DZ5mAC9xIRxy0WDcJ9gvxFqMaMVVjygOdAG3Uds
C0o0KpzW0AG4V+oFGKgowtBuAEGT98/uNpUldQjhKKWMCZFMfYb2K+13L7Jn3OYw4CYw9F+rVD7O
7jwzoAbREYk92FookyahudBwUf2C803nsf3OoDSX061iZ1VbUPBF8ESANFq8+h+Xr4y35QlMsBlh
So9qzRN8RJ1LqIcZHONdxgyMHSYi3pK/QzWD7uO6O7FCkA6V1udhSQ5k779cEynLV4Ja9UpMhM4w
SsdeH5pMt3MXd9MqOsbxjV77iySl+MtGKFSYctQeWqxr+qkqVFhEjABE9Sb8nJLDJaeph2uo2qyH
Pz9lHCA396kmnZ9bsbxmV+0S4ppN+mX8My+E1M/n3oSzGDnXIkJoAxLp8oNYt962DjSNAfshtXwg
LMtnwrP6xgHhR/gXr2CPaQZET77djIwtxARpNu+Q6J3sB7XGJW2agWWDbOC0VMNGOFE2l7UFb94J
NRgSu1XOwn0F/J8JDVz/+2koqCmSUEC4vvF37uiQofTX6+cGXE6tdAZkcxyL4sztuav9/DTwLbJB
TS9Aij2RvY567ERpst7abA6eeQ2uaiCRML9vTZ1jOS1uE1pcY/cI5WltHIeXQFqN3XpzrfOVXzFp
Q4RY94V8Iq90cG459aF1wXzGbVNNhGWn1xG6TOBXNQkum/SERWpWhJxbfNf+snDGW+Hr163Q4dm/
hGpSYryvXXLVku66plbP7FW4aGTjiIpFumX70bAOAh4++4ZIiosYImmOpyBAAk1kfIKgngxkA4As
LoHB4YdZUiCvELH1UwMOdw4EpbUAUxfPwEEFVVnFz62jbjEVEZCuA4fMMti3KwEY/GFK36dF/HOH
3eM+FIat92065b4x9j6IsoBzGqYYPtzzBt2wlzP/H1JQjmObBnlBBZfPdoQ+UAvfH6rg0IAbSXBu
rICEK6sVAI+2JAleBGrtCxS2aKaM/J+PgTMpY0oj+iddCfSog/a7q7P9ViEDFRUn3JnGOvPKbu9u
G/s+q9JIbX4VSc7OkgXwTXHoE8uQFMee58NhY9tfGZr3PYfVmiWoiqAPXZHMGnwWW9j8LIX9c+kf
zPGS+0ZIoIlPsRh11YCUDCCRK92E4shusO1hG9rpcdhmiDxenzWrmig+zh0/HB1+AgRbfBIk9W3W
s0PUktnbGEh/PUBbNB/63l5D/QHEDHhL6CQnufxUObKpUP2bNx8dvzfn0DAtT7d4C82p3WcPA+S3
A0Sw7AfnnOYqfIYznryIuRnAM9jspQNupHX+Is7e8M/7OeMPSbYkz2WjR0uxGtPQgXdBXdf2KfKn
SayAZG5mdoohRc1vofke/I4eQzCsSFHm3MEFMUTwrmnCyVW7enHtB8rhTEAzOqnn4NUKj/RMeE7G
PVgX0+GBPL6px9k7tYCHYMrPmOsd/bCljla2DLDOjEyM4ewLxtCknhGVXrPNKClc8iuDt3StC5k8
kj1Ze6vbbLNBopJbs3wzIwJzdP9VMJ1V5K5pqCP/Tc4GLrbxwmvvs2zFL2722+i4OALXEhHMKeMt
hQa/Z5btpRRmPpMjf71lVJ0i5fAwYQuMXBStlR+Hr5oNJhBim1IPZ/ytiQR6zFfZzBzOSTLuGoUJ
moixwpcz0SwA+wqlDfjz4Hx0ODw/SeRN/7EAU6Xj/RLB3QuyfFeI8rWGLUGz5rElcfOVILH4Z8Dg
AsppV42Mz/vm89xaH383qpDzJCe/dGW4zXk/otiVWr/XqkN8ECJFlJKW1oWea539aOf9w5rc4A/5
lP7tUInMVt65RxJ01U5wWt/zm0C89Wz11jFUR7fWfrEfGkoh6rwmlRdn6XUBXoa7StWTdDw6wl4z
wFL1vTGkwE5+4q4fZ3IQNUoQ+lDC5ArTjj2w9MJSd1lKHBTqJVhfzIKS39gekBl8J0FsaE8i/t5R
zsNlEYrXq12lSR9nll3+5qhEeLjVtpkwdsXT/FSDRhd8hy4/muQqhzBLUB7mTZNNj7PdP++FDmgp
YSWYxAOmYgFfuLNGNJqvQ1egzYlOjpkkzOZ2JJRJ6odsG8tN8Ot9yD5lXrLuCo/ttHcSqE+nB/nT
DBL4k3wjrg817dgffCRkm1tdGa19sBgjZUB+wwfKA+GvsOFRzSmYOK4VouOS1s9SGVYec3hbIzS4
+KE1NvaFpBecvamogTD1WI2wyTufoZaZv/O6YIKKydmbm2jelgoTWjsZN08uXNA7PvKnCYr6EQxX
k1b9Jb/mFY3Mq1Mztvzq9GTcAQO2HxMHo0WlU7QS8gIXpr4IKmBsISCpI/rVK/Uv17WKWmUaxEgh
IKr3V3CpMjT2glLKbWl0DpWjmeWJyBeu0E/aYVcl0MLm2l7NbY3kvPQYZF1bYy7DasHs2NDPOijA
zpyITdY8U6v4IO90V0K3IRokMOMvqx3GHp/4acid8xYYl+XtfRtkJ/7HBQpBsb1XonSc6Qjxbp/4
uUUyW+AdZBxTv8CNSxZB9FMdPXUmvE5VdvETddwEu3FwEUnO3JQ9AkuQEgoTs9bjZAEsVRZNby3F
qROh/Chyq1nmm3PVHWFpsUDbVCM55GLRUkRWeRxaoJ5SKzXv6AGcm3s+ZLNBfqX9VrKrKALzqzeV
CZ/PvuxeF/W4ZY8ccz9Rle1RAQ+UJNBo2y6jjp0QbHLJ1OZ9AvNM3ZQp2Ly5n2CztMAJy8sX7wp0
qY6fX9ZhCIKplmzSxfFdtaQzaf4DQOeCt8MnkxFk8l7CC7y+tsbaAyPzphUuyuoI8kUT+AJLm5Al
Rbd0fuuRzC/kPzgPzaoIw9B5TxxkP7zRr0EDsQbvqZZDkRj2IUNCvzbDMzbeFGTAlyX4EJmRxpnE
sl/6BWuV/WXSUVDn9/QppSy8adDTCy+y6i57tMkn01B/TkjhqgVWZWV3et0YOK5gemlpx1Egu1sh
/hmsFKZTEHvhY+llQe6Xnq+l1WEAvBqCnI8WykAVRMAVOlWfjgc/APSokmMTZshnoKEPR1BY31MS
gJA/uuoSj75beXcW42msbEeTnMnlHxs8tMSopHkxetLpizJADdEdR4ceZlXgP+mwpK9oaHD3X0Og
RsDj3xOm+ZEImDK0sLHqx7/+KjDAbUn34NqJquIcs0wS1Kzb+6ujpwKMPqHBK/O+dqudgwEVtcTt
DwoQ3HJ8cmbdaFOLi9grbHBNNo6sc/pe6TSz6mZCqRMq69Evjfe1Hdu8+q5m5VJr/STJDnsQRFnH
ZLc1/DH6Ub1tVP0H0n4pwaKx3lO4OCe5NmvjekOY7yN2Kqj08A6SBVK5GLi+3KottL6TUfCDq2Ux
2ghXuGQc0yCWWHGjmfiqZNNUYsyjCGFEmVhz1I2vQdu5a0Aii/iNSYlc71Hf2agLUqYn+C/jAnuZ
EclfiihN2WTLzhGSlmJfYFhEhglQq4v0otnNsX18ApmqwEwaX6G58rClfaVh92pMJ1roy/SuFvrc
qSLXpyS567+Ahdzh3dKUzkwWTE6iDVh8seIPW7GxXy21D+/JD5xVlBoUtluGQ90Te/YwOHGo+/hX
KIJAUONk+tnBi++mORIGV0fBojKd591kbQHSrSsn+2EBhUCxiZhtt4mn2dJ9vGe+Xd1tllsIGoFK
FYImVPiOAfU0/zNu5bOC9Du4MbkauuEmMZS/6+ljBMlzPMI4or58eMwQfCiwCyIjkWiaPc9r0yKo
H3mENvRfb8tuNfO09E/Qps0ncIhZBhYR2pUYA7E9Mxylnl/oUa5UPgIhA7Voe8ogE++PzRoz0Wj7
I1Qg/nUP1w3Np6+DR1RvgEGn7dAFRU1Tt9bHE/jvqkDYFdXGBcz8gRQmD0+Y6nNEcDkObCIqQRau
BzEyYLnMP+OZIy7vaKkX4Nuq9M4XZ8K07BHX13qdeg2IG71xMiCiUglsbDOvpqrVUU4ojhDNCqJN
lgTUfFg6uSrG1AhZZFTJ5meaed3mB3Hk4CeWYzhIECONI78pfj0fEM7L55BzRjzCpXMKHX7GOwJX
ukYgUFPw0wdXbDvbVPpY05LoiKFjZDX8k3PGhS61RAemdeSf077t9tZ7cxS1ceLIgd2PDnOIc7ql
ssBoly/tDW3AOQIq0gfSIhGpYEzOXBv4a/T1ivfXgVjU6zVRVx4Dnol1jPhxTlkY0KOgEEtlk7bB
4JNPXUdabTd9kKty0afUJp9IR1mO2ZF/I9GnXFi+YaQckF3i5mxfDMAr1sPDGdU6oI5vCZRfCnuW
c4R3SLJJ2aRb4nFhvJknSkWc39+cfvrMtRnYM8hKXi7j/QY/VzRBkiRbaXT+75pTNzBevxb6wA9D
b+ifsg7nLh4lm+YrFp24EWMI0oDXkObk4YtpViinODym8TaHGh4xh4m3Ywhb50aFu7JUmoQISajq
uBpQUNSlzzM1m1HYdKzzgWaGNWY2D5oTP545Cf2hLrXDOIzwsk/FLNry00JTxEN+TgQtOYMfyjEr
lno0GH/XgrlO/RJnoUePN6wnRgAxpXJ5Xx4LwZxTBSjbffS9tdoiZXtiHAPhb047Nw6P9ygZ2gMI
mOHv3s0DGeHhi6Et4UFo0Kd5lpChGpOsy468MRFtuFFYTa/yHQI8qAVK8qnuangO8u4hn7U3D8qn
1iLTbeuSMjI7jBz0106/tqZJOhglSpJ2xzuqXfwk+3+LJ7wWB2rbjp0BVBH+jio2RprM9lyPWlZX
AY+vbTkQWoijaKPyPZFBP9/9tRH8QSN3n8nfjhzM+RDCBNF1BcuoWKR7DhEjKpJfURzb4+iFWkO4
x0oh+CSiB6gvQJrOn+7kx1Fhs5L5h2TYixjp66rc+rudIpzHLMW26o9vaFjYeBA4OT8/kolZkrx3
I0T0vj3fR4rAdRnOIwLxq0X/dj3yGoQb5nwf6FzvYMEwYto3Oo6SMaoi95tl6udIHP4KuzMyqLoJ
Og24cx/XnAWeGBkINNZPjL6MG+M43rRCgGSY4ruLJkJRY0sAgSsTvJYeUWjyjuUnLrjJheVQEJIK
g+se2qNroIHRNlYfza52oSr603I3rSI3QHnimPUQUPpIkj/+8HmEcqiGobmK/cB2/GpPSV70k8Ma
zc1yblpWaFOljCGjF/UgfO+rOjKRW+jawR5uoLlvdgmZzfM+esdqLAnyahLKUY9ZuKekaAV7Z8QP
Q5KgO5sAuQ5Odb8btRk4XtqWAmw4hPlsKd5IBTBR293jAS3vVC9q3qc0dqzOoDVnzHLVO+tQvgQ6
7tvyI0MNoI/NOFMnvx319iQ/fq/sSqegEHZqnefzwDJUk1HO9jvvjKGYNJ5KuicJ4Xcych5SuC/B
uSiMed6CM6fo0Z9FMZCNwJSuIKmIQEm3SEPZobToDYXhNyr9T9IHmmyNttCbgpYWUaJRVrAwkUzI
+n73ePbJwLxVUc+ho1yChRrb7ftZu/Slv6I5ii2zQ8ItRuyZMpLBzP4bU+I8ubOA1CDCXZHGPgG8
7I0kpe3+MPz4w9F3BYPf7DK3KqeqT50Sc1k7R/asRWCFCqlIglGsluaiY3GE/nAFRtYpw1u4/6+j
zz+7SBJkRKihb9Ppo18jitZu7eI+baQJB2VLeqvdvmKRpT+JpE11IB1j7wnNsPoUibvgUAGGvaPn
/yXVj2KQdSygDWFBwuE/5tvh8UWXTK83eXoZjdHjBn7ENr6VrBfaRMXkw6HsyzeR9uK6sK7Mbbxd
yoZJSpx4hsOwiFyOJVBfIVLSw7gO6vnIWFJApKVqCadoDjmYcerAhxXUgYfZUzUPJQKqmV4AKdrO
2GNnPBBJINHxmY85YYU80FeLgVqZNYqk5Wdjm8kCHP21CVpmM6q4XlW65Uim68ZzGiLIL0vjU6R3
n9RFLK0M2OitoZRwdotecH0b5ID6FRUqOvjecEfC1ZdQ1C5vEWhaH6ES61bBTXrz0VieAgEeLw+R
KUkp+HyKGJVsjFu94xRiF8RJi7hK3iUU/9q22iwYf+AK7P5JbrZxYqXuQtqEzcHJ9feHxQkkc2+M
QJjcEcCawOkqf/BxGw+nBI7c2HDxaMUePb7xuL8u3S0OwuLGIH8gkJK7E9q3l4u9G3lvcqulHbJF
3d4Pc27g+y2hre20iOndLBF+TUN1ajLlXV6WwpVIVuJzHyQ09j/ThD7vMKqnpnELSxKDerLpJKHb
PfeAUPH2A3JEfayMkr9fHlWlWAVxK02AIrpypbFYXJmSQ1qIJRMHtQJK3jJTSpywD8LEeoBAP65r
+4z7jICWijxHjApiLjGZrMUQikKs8nWByv+014WTqjQ6UkgsR/OYKf/7GXaRCqxypaSoIAkLc+a8
RJpYpt92AhUalLpVq7Bvst/RJLGz9vu+MAkgOTYEKbyCHVhjK7ysDiOP1NQONAgXtHnyOCEsKZXe
r2JHUCxi6WInGArA9SC6Me6OECI7p4D5edNwXPuZYQ/TF32EOMlZ+gyHVuq7TXhlu0ijgCst6iTK
/XhYMaLoz3f2+eTfgSKF18Cq3dInuK9RYztPBT9Yu97PbhZLI+CuH6xQ/rehOd/fR+5g+oVpNc/d
SKqDrjzuMK5veqiAs327c0SXI8tljAxj4zDrhA4YojhuvPgoHe4TTI800b+W9sG5x+WcYtAdiAeU
02b8VVnmhOH9EI5uG+NHEQaWj7cL3KbfiQ1IGt2FoVhNkoeeUvXLQ+bTImayVN3LAd63SSYk6PwN
vN/NGx5tcQIr7cR4Va5KjGH4WYXGz8VyCj/XP9micuTmposp/NeP19s4w7bCymVoM+6prNA1eaTu
DK/YGMQSBs3SwB3IKkBFe5Ye4T2zwJ3tWsQPx76jfOP+hs8ORMyCq2EOxVvDLIMVn0zc/8CarT1R
X8fXyiIRMH3mZsokeLi+iZvo07J/faHnhYBKSa2E0WCgAdGHQVEfZnvCf2cNRPssz5Qo2WjSSCgN
iATtjoVCfROcD5KqS9t1xVQOQrXLwXzpWFplB38Gb/bXv7qX6+EHPaMXGB5D9pTwxwsd6ECnqVqz
JvrgK6JOqEZpfTCpv9XVGUm0WF45UH0DyY+P0+CYuOVBJdOtavqlIu8PRYLfbGfreU31I9NBx8rc
vQRRpefM5rJyXn71HcDDIBb1nseYUNSLUzMkGjE8N6JgB+Mrhdf3or+VdEDFr2nqjmuN8J0YeI6a
khTNG1tnzNRhQpS/ksvUCXByKmyGSiemcOoLYozcdDAgLHSmHInaCwW3pGIupVsEFkyZ7philUkA
/bRn3A8Jw4JZc9cvs3/UVRFYAbpn/LwopauO6JYBnMqRqH36LmOnWxHr0MWdyiz5CM0lpmxMZ6MQ
I8hR0NJq1raiJca1oxQz+EtgRqYOAdMaKsWV68m8Llg053KQGF1MzZI6XO2UGyIYtdcT+Fl8ksHV
OSlaVjFFeQSV8JGfFkAQiInZDoOaklXR97dU4Hs+zUvWbZCh2sD4ee70etOVCh4PlM2pYgP4PgBT
5eidxvT0dBimErZi7XZ0pX3G7RW9WvkAVmZDRZEmfzZ7bRI50Jod9KDG3voywrRfX1hs1DrDMnmF
XFc62X8r9epcN6N4kro+Xm7EM9P1uywTXC1sJ2wO03h6NSUZFtGC5NlUwsU+C4scbRUPyS3Fentw
pLH+PaLBfvYCX6eT9QptkWE4BpfiMLMnDfzS+6QlQ8qXI9ChX6x5y0J43agCaz8nOpQJVrEnCoPS
iKV67pPO/sumA7uUXSvjeSm5jPjCfVWD4jbMSTY0WkmjLiqCFydOfJQtYqPJ8yZ9LUrHHaw4R49/
HZFvxULwYnsHE7dw/q2qONySG8iVh7KbBvdEZI4QuHXftBVBgzLqncCWg6LsJ4b7e+YX1V/Gfnj+
NsSxTIB4LC0IAR/xtnCxDcNR0giLIyotqjtBgQC2O0qNvfmFZq/xx/nuCjN7QyFsQVbSMeNWEgZ0
cQcU8O5Jpy4R4yrBn9dNnHWJH6mPFZpamF+RyYvvfOAkxSxT+RpQO2pcENQL7At1uM2QoQlqV/Pk
qZCYPJesbLSaDh7LmR2gZ+8sM6yplLPByPwNJyLFT1DYygurGNIw2qHnzw1kOM4wviSPFqqDSKTH
wdSJjl35EoW/2GZ8V9l7vF4gsfcy4iWaeEGwSAqhm1sfya1fWdjsTMcvNib2TGDpHdQyRfeo2Qsu
C103iIzStf50IioXCZ/fSjnPI8p4kp0uSalSxfLnotjF2ch/yOqFzq89H4gsfnpLgr/NqH6q8sdc
IRhWETyCxhUoWPob0xcRqpanRN3pAeKwjZgT91ig22fY1wecVaPutNV2S7LqcVthJ2z34au8cDPN
raeHuTcnKcKN0xQ5MkBMRaYLsjb8AyeWKwaxjPr5bvXAV6ZM83ezpIacWRqDKumcVtcKpmF7LQvR
tlxVpGx+o66LP443dfOygWCUuUAoIWPO5ogfBptDRnvC72xTC5Ku3Lo6YQm2SI1WGVLXYejKZwD7
8/g6uN0V/skDZYWS2IMjDvWtt9wJKBo6hP+f3gRILeSh6b1OIpv6BmNQ4A72LtBAmKs9kChizqsz
nbPil4mMlMjAL6AZwBz6+D8TwZMRJOvAXSSkkZsJCXi/Fcq4mn6/K2V5kZiQO+ixX3z84PN3Q5eF
aVprgtqHbGF7HV3PPv9WbsgJ0kyDSnJXOY2jQGpyCThKvc+6/elZBetpKtsFimAt5g8iMYd7MZCX
m61B0UpRv26wa5YHQcxAMcwA8vyO2nA2tPEFZ5DtUk2yyjOCB91e33WmJQAMNuMp3bkf4/XlT59Y
XudI7w+6eHiDWV6FsAx3P2qqDMALaFoOQLVt/C8FYy+xjPeD57i9ILYQ6aRMR0zknvxAWXm+GZpg
wquZz+7iVo27ZvPAvA4RpHblpd+Ki4nvPxCGqkMpACt84I7IL9vOvZHbonwx4QqTi/3kzgy2GoRY
oHTNMBVW6rpUpr5JDbUmSiqQrynjqb9Kct/JbHiQXwmo2FsRzOSlXtHv47CwXRRavaAG7PNZ8JYl
nTt+t/VQ3j0No/Hezzlyvv4FmjZ9mAAGb1WFMj0o0A0gCmttNljC3WrStwmGCJS6zc1faps39U6V
rSCsT/ss5uEYirrTFT/6AnZxHQGN3z+rhV1qq2phKIZAwkotrKSdq89gsw7Y4d51vkTjyu21rKlY
9WkP6gFaFIUZEyk8heWBAOGJHlLW6bImvQP0aIGXCIZWQyvL3avVBuC9NCFHxPZ1WNrXHIE8qWUp
SaitCEjd1n6jmgewIe6U5IJcKcq93VhgQe4ard9xg0crRTGFZWno0VnU6KmJSd/YyDl6Tef3NW/7
dHI9qd5ToppvCLBBGocacv4QYe+bpv3Nu1Ofsq8JWYMopNwUHG0JO7MjtUHPByHNGhyyBLPj9xBg
potEa/P5CBhvR9qfcFKTlreYCmLGPDfVkoMQ7A17b0CN5DBDU/30hmvWzzL/smbFekp5cCgVuS9v
fSbQq5KDgWp1FhfhwJKwxJmjYXN/0IS8VQu7FpW4Kn2dkeuFXebU8oqO4BCI4hyyNoWA3bsyDaNT
s/mouKvN5U1y+ecm4B8tOJ6+Yuq4Xm3RwO85kieBZtIQzjm+o4v3O/FSwTn/sbcjpR0dI8osgOAD
fAc+jPM+sA/oPM8tO4hgus2sWNxOldoGnr+GRwev/Hgjp+wVIsAM4Brs1WK6Kc2lVT9Bt/bb9SNw
JtLXfxzsNUJqeoXZFFmTysMYc11V1LVLymaiOl/p9DK5ctnFZqGE0ZVzM4TAQh2sXZm3y6MFhgR2
kKtJW0qNclZrddbTySA1m09vDJODuF+/vB5iyqDHYxl+8laghz6NWM7rPVwczuTO7jNNDn24BavY
d7TasGcSBCmsb8HoUg39EaJo5Un+L93eUVtaZJVNygrFZsaNiUvMIld0t+aDIw8Z41InRnM/hFmW
iDY0YCXBchOxQSa3j53fF4r8t8Q9lZHBF7jOdIkbkz3sF1mLVwV2jo/KXveYCf+luJNVGqWwPZNg
wWzQRSXl8zwZ0DveGAxflXz2AOT3UQhSRKF/Hh1pPH87/80vgB9FaYH6UYsYL/flXs7sQAiAr4Wq
KCzKzQt3LnEOlCEQTGR+AhNgWEXdksQKzaxt/R1uM7RWqEfEeDD/G5v5gJBX04Ui9XwMF3ilI1y9
J6fDa9njPPqatsi5E5YW2Qv/SnFxLVRZe+5rvlGJnRjpi+tGcQcTgBXauHJnlUzq2Ab8hcOiV/bJ
ejnYqlkfNHuEKmXi+3zXBCT/X546+LezGmqJrLQVfUpXleFRH6rKt4LD04KqpLwp4hbBMIfQmkjq
nc+1tqTFMB8EkQvNVZtPUaneNkg9BhVR0c5KNCTIJ/MJcYw95zzBlNB4+2Ixr0CMCt3RycasCZgs
7xLQkviwqv0U43dAB+hbJGBglrDYnzTi+N/nad7e4GQa/XLJ7Y2yLuT1QQVQ46g2HfWsIzBIzpk9
/++5FTTOY6n18ygL6lNRg9ugKKjEIekCatfys/XDG4rnYpfZJScwbM1ooY0hv2T8L1s2u8vOU8I4
o5CeMeC1x+XWrhSr8Xw3g0bb8Inyxvp+CgopZ6IQO8C+cRcZ21vgRiZtcjD9iS8i1hLhNrAXdXH+
5vlftShgIpJfNjDTOKhNd61JRQbINAGIm9Ec65EZLSUzJa4c5bhSGidJMQaL3xwBs3lGWbplTPYw
yL5vzhqQ6fzACRLZ7PKtVX+kiZSqwTQQYIjs5rqmWqtYH7RJ5+o0zRjY/2TDJqKeaMCyr0Apd2Tl
cCduU9GXnugkYPm45nT+qU6BfqCj6xBBZFKw022PsA3/Q8wCyL61Bk8TOLN6UKY3t5UHnTveLBY+
lpTG2lzCJOoipzgJ0psixjxwgv2fv3cbF2r5AF/9XqppZ81UFigfKaTWziYAvv7L9aWm5gRbvkL6
jAWV+HMdkOcdLWJGpZFM5DOqbyiIfYg0dtVlPJOfuMQm3Spmuz1j5xqfOXOrIXAZhqF5wxl5EGI/
rTi1xHTDXfN20RCA8k9yEUsjAjbvhccXbhJfBulTzktREyF09PKAeoZO0mfmcMchFCukqCZjIccQ
cFYdsk6vGH2jNgvMALdEbx5UmasIMiG6RX9dGWW3W5YJX90L2MFsPl7e7xWRq4fPEg3DqczERjBL
qvdRXH1R+zJ9j40d1EKVwnLNg3xV+UAlx5W/+eMqAyP01GrXeEqVcQt4MvOrJsYvUQOs3FaKKkqx
TQ2bc5BLfLtL9eNVSmxScfZuKh3sDopJbSQDpzxYhLopncxgv52OUgSypD9zouJ/3nQIx6CRSUKS
CLxnwmj25hBCtF1+PWxOzQaDHP18hDvm9zWbH05WtRx8TyRhIW2nr8j9R8V4Ll1y7YmvC5glgp6u
BDxcCPuk7MDrUMGub0JxnFF92OprMksw6dKtDimADrxOe2DXawQf6u9Gc7zmWl1sqiumRWXMV0AD
GUilGB0gpgzZn37ZmUauI1emvVZIExxc9J8acUH1sRhnrbUi3FeP2Jcp7/6+T+pRXSbLTXrS1zf8
kETtPJbY/9DejJSQkMk+RTCGXwWPaEfM3lYJknEtfHRlIeWIOR8ko4cJHtPiBIpHcru2RnBVTXT+
zrqlXtGkXUSM2E6nbQ0XOyxCQWZoBwVMJPJ6hjY4aYUkzPY7LQ4nSnvAi5YOP3+Vdg5P804I4CyM
PIedFVbaWAZY1vmuGixh3k7EgSPEVWxg/tbRZS6gQ9I7W25mLnV3p7//a1E/83HV40CxHgwGeGQs
rgPKA083xV1gYNY+tM93CXsntPnnroRmbQjYQ8HaduicYlmtSVfikK+lFIOd+CRUPw4ZsLbzvb4O
3UQFXKNLG1J1dJr2DraQDOHZqVeubLJ1/rAuPrGrBn+kB5Qafyp14vcGByDtVW2fmueCAOA2ShaT
/oxW6PoD79QwfCrIl4gNpQcr04bFqy35d/JJStUJBuqg0TdOFyMePf2ZwM8LmEkw/LF5EGpvYi63
M8e1jatkxSk6Z5g0g3BVKI/FtEuI9eTa+3jqoKg8rWIC9SYnFww+Q70SynXtEt0BBIqErzIDopfG
A+f2GiGmu8B6sgljSuetmTCdqYJoEQfrVBHvR2j5ZTXexXmpLcKEPGbJsD3JjUKJBoj042korr0U
YM/ZFTCiFvq9lXFXVWdPfmjWdeMVx/hDv+NTiz4EeIi+joXlvsjqv8HGC1WBWiFsJmNvF7DHA1sZ
iAdyabPA/UhGeFdcnuN18LorXl18tWYVcsk+1ykW960lBq1J8hW/VSPP9gzIph2KFIxhFET99Ll/
L91Pf//w1dSnAwjdxqx+lR5M9HeeVomr01d8cyX8lATeDE0mz8/Um0/v/nMIeMQsbvBkjcH0/ooU
Pb97qv5AAK8eAfiF9lmSveIM3R5XvAoWpnewTrmiT4fFoGd6jCYUBqBlLcCA6yjFMadm8sMxIh4I
PvwrP/0kAVO9oIxkDwbOj0I4TBId8FYk8aUYKzOP02PJ0g/g+sHGopZV16SGptkng8RrlLvit0KI
187EpNPi9oZb6e36ck507qsDmaYigFUB4szhGn6j0vbsTlbevzuEa/BsJ/P1qKqW5O3KLj5yv88s
/1tlA0TGVAPp+JEqiSgEqJXsbWppyWQh0eZhdW3N5euzp7Hu5UsORYNIRrlMZeTfCpES/c9GfBxZ
y2e/nsdkL58pVh1Ut47dUXGMjSnuOAPQjuuk3Y+O2usjiIYEDPNqjNEPuyF2vj03esDqaoCBTuug
0+sGv11FVkNRqopfSsDUMX2mAKLn6gsKFIWtrCocOqzypCe1Q6kzpx2XrwbrmZdN5ku2PZzS7qLQ
s1zHoDblsIokcDSJZjVy1uEf1Z5HlObSC1sUEvS+2wpQuvH1dEAE3S+/Kbayf53QZ7RTKuuYfBjT
z2+11fNEtu6OTJypwzOnb6Lduyu6+inLl5kDfkDVTsUyUby9DhMUq1l5WmL6VDXWcEjK8/yQlPmN
7rKkzzTGGF5kDVkA3jWO3+Xi7ypMXoP87NNSn8OHVZR4GPvkKXhWZcjOCR29m5i+eHps8MemVjBN
6MfSVC1ZcbudjuJkTZFH/3EuUGwT4NYSnyoMrEOydbEQisKJp/q1UGphwWmhkQRRUu50s+y9LMER
4hevNMya2e1fWgYU792uor0Sgm+ZHdnWhx+BU/PLzym7Q2vb3iopzztb2+ugdUAFaRvBdXyUqlkC
xp+6bTYPw0eJNfxvZ5CmVQ1Kur5d9rXSu3IPfqS5cxUKmsVyc5W388SlqCa2SPTHX2lJstMMAE5B
i8sx8h1KTrY4dFssrQDI106bUDpZl2EHUjJ9v4GaXeMB49q9e+I+P0e3GjSVbKZ05+Ra3wliBCO5
dwX+auFkXug1MlUXYr1CbZiRyO/2Ansz2sfed1JXShgpeDRm+nKo2xjh/CJbYGcvS8v4Fc8vKy2k
sBYHhrGH1UmrS6e2GONMti6Neevl9GuQl+9fKZmQ4/khbhtM+jCLllTetN5PwZGDt3oDmYR5TH9R
EQkUfqvfS57c1iBRXoPULI90x3pzw5Gt7PUCm7Y0f6v1+ebd6LtoI1p+7T41kxN6WtHFErjcCQ9k
h8MtjWPyNU57cmCR83GJe5ZDip2B2LnNRt8DIPRcuNZqxxWKUk/kPD9rLyGOURFf007MNiZrggZf
BA4ptnBC3d7VbreJX5Xnhphx2/1BOvNSMUnK6QtEz+KdhzBeOV/wXQv+PMyEpM3b3MmqGl1tm++J
MBDvH7t67tRmWf1vy95WXJBjkjA5tj6SO7g6HR+2Jx4nhqIwkQ4W5bYm5zwsEG1gaYONV1i0264x
38fIfGBPADZM71a7rivxb0K1pFrfxaZm7xo3Axsg4w4i1FIF3rZCFQTfAqAFBzMDkcz7eFL3M860
3x4G5yy37+7mZoEVMc1B3G4Hu0Y+kiz5er87m2kdjxsL+H5ks3dIfZqMAepXfd490V28qgP6xU0C
OhpQJNr8TtJJEavjoY8x1IJnp/ajuCxTwt6XAq9JOAbKHkfrKfmRRYfCiCIdO919srAKxu9WtIeZ
aNf16dejY0jfMd3MjXsTqargGtLHfq8Pmo26JIDV+nso3HaEp/eBSJGipkSFroCWBmguNuVvoTmF
tRDBBmdua+Hx/woM9rkTp51VX+N/GxUMMxaOpq3yOz7kt0SLHQdznVVb43RnzmXfgagKMPbg34F1
4rMFOv8a9qNx1uaZ+C87UYch7PINYyoEvYNhuWzac0/J+PnL2sJ1ImbMCanl1MKpJddtqkCGl5Gu
ATMeJDDNhfLdcgRoVaw9seYv+F/KIhfr3C+AFe2gE1yCxWxgVsSSA8dcQn6pqwqUCJ8kEwckJWNT
rgdR0ycbBccXzFCR/tM7TsTrwBUDz9MRAARiAUYrMdOwxJgpRq7QUfNs63jMB/8MddAwLajsFVYy
eFDxZXYBotdbZ40OyqLwQeG+ladhXm4MD/S3A2iYhKt6nxzIWw0/CXAObA399nrbmbqaJz1/u4ik
Ss8f6JBdxwf1F5xxPE/QVwZ8zYsNOUVSTiCIz7DI3kM2vv9BepvTGu6OLVhownQ33H4++HbR2OSc
6GCtRzogQVRUXLtrInrB5Dai+IFQsFG36iR6UcQKSs0jRh7ecFIZVCtZ/DROycfIyAqAsV3ISB28
ugp1ct0WI8sIlpfqnyTGj2aXWCWOYYolkbxRNdx+bZEOXvKt8mAcRn1HDdvgwnqn21HS6kGXavWJ
qkMSp4WwzDFXi4qLwBA8jz8VpAzo2PPwmeLljBgrngbzNJd8JWlohj48ycbLARG5U8pzs0ankZ/U
tzxPbbCtuhyN171tR0m8wrcQAAbM8WPCDz48+RwCwo2UiLS9yDvyDTHB2nM0YGDiA8Q8WxTD/b7M
AWQ1Av8MVlZYeGgzSeIgXXiaK8I0GRXV6pyc7uwY3tUGg7EngJ2WeDaldDRYvdBquhKFTE/hUGdv
Yy6NmJcZrYROMaKenB6zB9IhkLOghydecRZC+KTYNKm3GI2M+2okPUVBSK2x91AVK3SY9qsG1Oy5
ExB4Rr7AWmvq7JZmP+yT0j3LhO6q+khGJ0N1ikQ0/rFHNOKjKhca79FuTsufec3JxAQVfO24WrRb
vJd/zw6WlpWCxtFRe5aFLy6Nl/rNOukixJR54TKMvogAeqTFQyulmj5sYFbyStlzVbVzTeEzzXgQ
w6Zmz0TS5KFNGDP29ajLc/Rhz45euiFBBBHknEvdazxPi+5bgeJgsE1+v4ffM/9L2XUUJWTYCChI
iPJD/m+vvvou2vi7VOpmycKC+uRJIAUoHb+G8MCwF458OQ6ODKgHuF0soV8pFGUlBSy3nU24KkLa
jzuCPzmiEA71XjXy5v1dO4LTD/flG+NWcMryI8ToTCVIFP3h9OA0BsOKYCc84rfkxDB+EKRWak03
UEZ2yKKttRpaoNl3b/8cJG4M/GRsc+IUhIvFR77jR0eJPYB3c1lNcP08v0ImdAb6mb31xuD3JFas
A97QWUhLwtgMVMeR8qPPouMZf4Y9zPq7nVNHIdCUgiakUbm9CgMGKF+HdO33c9wApcM9oTq2SKhW
lSTo5D4zNByXsRCOuskBzdSshWXxGLm4r6U+Ju6u4u2mLcMCvvlV7RlGANiJFEGqihEMRkF2OE8Q
dhCKZVAZp59FqMUnMPg+IdssNdlcMUU0mnUo9cgfDSJp+CnY0+QXG+AfkylLTd6tBO5uDVWlTf2E
A4kt5Onsez9ct8uEHnJxTkKtqfZXz2fDfqDFCM9njhuPj+oWNzZa1owrZek34ZacM0bMHjYHTcOw
5Pb+EExpzFbKjlPumVXgmu14RczJRkTnCVOSqGhsZJFS/4YBp914RxU5yESvdnuEuJGQeeuGEamp
OjKDI4vLemnNxfdDnli+cvEb4MBX+7aa3lXhaIMlGpm6/UnUbjWFs01unZLNXBqfOG/7jd9U06e0
pQM/V7Zz7YW7jsVzsDFaa/laUFzj1KZIr/K29FVolqtd59FDwPH5AjVgtbvKycWcrdrL5MbrJvK7
NMrv1P6V9nL+fT+HzhJh1o4UaPd49ZXMgT78DdHl0xcnYCQiD8ngCDu21YURRpploCyGUXc6WQA7
yF9eSgkvsMJtBa6J9YqtOkAueyncYYUKx+FsQOloRVbsOchhoxcMSjJdXk3VghV9gANnknee7sbs
Pg4ogMMXt9Rofc+6xDC/mdXQyw5fxgwpABAKTwQCn7xH3B+Ckd90A2RhonJsklrxlbbPVD03iZUh
tAuLcRxOSZKrdq8tt/4HkUa5KPSgSWxv7qj0G1m6VIeQH+8iOakBx4XCpYdn4ohlhNFvKYiUJaZa
iLrKtvVq5Qj9hpKoE4RsoCCVo7qKsNyD9FWFg0UkC90fdl3A9v/G3SxOjEIN3cgU9VXO3uNWADOj
m+rwFzLSfE1EbihB9nF96bNnZRqUXFuT2KzDVuxJurm7sXZTE2ZEiUhivpzCpaZ8C6RvdS51Wk9f
ThwhtG5cUw48TkM5ZTr20uN+vue8kCMaaKbuHTNPLCqOvk3ctb4bO61fQlv9H2rw9pMJLLmA//0A
OzX4V5nAqJHDKMo/okEDX8d4l/xvzo8oXUHIYu5nk40CENQdZAgbmvtH5NNxHNjJWqFeH/r4OIzA
5zAk0FQVXfsGmciTByBIsZGHm8fhwlz53DFL4dTYsXQ9rkHbzMyWQJcl9LbrgZAmkwva08jYsVAV
tkpQ+PPNt2BaKKYHp2ipQYqPI5LoIkv+qpXQBESy6Xn1BAJLAbUsu9sGcAYhdX1Kc/jC5m2Wq5Jv
QRrYjzcDk9HIGzrESYGYvoQqyKRj98PsBA7xf/P+r5UoA4XQGBfsj6nsvI1iXbbuvZfCb9hakyYP
94y2/vUoZkY0t2S8GfoeJIXZxFIJ2+VZj2Eb+dNvwowktq41AdFLFUnCAituh5VLs/AB59O0MFus
BuBIXZnF/znNV7dReKuR2/04EFFk90rEHItNgmCtvFETsw6MZtinYO7S4ljLiv+mNDHpdVa2uW3C
ZWj/f9nKeyjsdWt/BzudZ2lvJIS9O/GjlwezG/4wcjBEgw4jOVuN8bpGP3cbrg0vMGgcLe3bXHBx
Cyzb4B/Li8FCb2iymV3lLfiiogHK8ShyAMepEltatWp4xszNmpaHY5zJBGs5behT8u0wIPoo6aji
WcWF2fE05acA6kf5uazDleYNtP16njGTc8jAqXkc+RARLgivZnH3C19F1r/7JkWEfzBSrnWr01Yy
ChHh4DcdQGfGozqgLpNfmFXYwjCDk5L5piDFaWd+xi26mJ2gx+MCAAtS9r2k7wbJL22XOcm1PrNF
tAwA3ZvAdMjR4IaL5pdlkCKxPt1JsYLkxVTig0lKF4ens/gak+f/d4ZcjSBmpEMqCz57DyCJgnnb
94cLMLOBgo1hzuOb0unqxql86KjQ0U4J8TCyZca3h+N8tKmT7NacmVSMNWlOihphGp+XquR5v9MX
h+M1pMs/xRYeeX9dcN1OKPNMf5gE4vttGdRQZjguj4OV+5Wl9fv0pOC5FDdr/BidkPW2lJhxLUgb
SnUcY7eDHjZ4b7F062liOvZEfLjIoyva/2kP2moaJPcuoec1WYnIOlsUyuauyx2GVYd3sqm5diZ+
MqC0WebPEr2COkdlCd/tda/ieY3QYTb2QLCfc3LnpVk5CsC0ZWLQ1xc7eOIbsYXuYKMWHnZym9HS
uwShZrbpTyVkKDyMvy5L2DX+N+S/IZbL35QXBXbW1GfN6j2NSpKeRUdccytCiB+uOLTvugtZi3uS
rluPcaEkdXnQQjaVVrgkoyIYKrNzj31Xj9BeVLuIdlHZPaSTKcqfY5Nj9hS20hsJ8ZEXnpeVmCVg
9sx8a9h8/3y5C5IdSmMp+lfQmrz6So2UBRtJO9wIb/rNNWeu7hdY6Z8eKbEkK5W6f1X2eG642eru
zmZOgynHUO4+pW85j7STPYARgN4ywvnt2gFCB6nTVM0NeMv1/TVwEuV1kTQWBUBxz1J7GUuT4vhf
5qbE9pZY0m/47++himl+WHfQ53Zdk1etlQa6LeUINnKIdDVdxIr32W4lMp4L6J3YxluYZDl0D7L0
0g8rCinjhCunGAqV0sqJGnAJJOywCbZSROwt18UYEGPUzYvqMzCFIRhlANZ+kOtY/xEA8tfLv9qk
NVqaQOVyD6od3InqGrRjsH64qzclwmYuKKvrt4tqnsi3PTJsBfd7eCgU6/4HlPFB8QJBHJlXpvjm
zTK7mJrCgqiFufcwLgcSv0MDEXSceWF9Oxif6S8MWXJ6wTitRWywL8OZaW+Qy33Yp3Mxs78al1cC
CvqbSoAFkymAGZB/N6RXdZFwKGT0OjmQ0NWOg2u2EUydn2XwEJxn+uBNTOfsDBNyBPOkr4k+tclX
TiZ6FP3SN93YTV5JddruOXT8pHv0GXM+ZBh0/f9AwFqd0DqgJwhP8k3vSJmazVbYPLXx+EVK+yWM
b56Ty1B0hRS2/9VDzTq1JT9N/6OQg9uX8nUKXPRyDBglIaLJ3N2M8Q8ryoPfX1TAA+ICr7SwH3Ye
ZP2Hrk5+IZxhcnBKn1xBC9EEmdvVMdIeETeaVXBZPlV5v4rKVc69MuKIoMk3jbzkwEhL/KIL5exi
0UBV10MueMZPFOuQGjwNPW6MdoZYh+rlEj3yC5PUuXYYFtCjcBnGRiWn6nv/0BK/Vw6V3NwBASIp
pJTj5lt4YNcZA6kFhODFaQj67mX5P2s9xkuGCRc9xqvimeT5E5nIDNCXPtmWFb+i19CzxuLU/Nx9
Y+kOw+CLDBgs51VH8PnMcNqnmBtbkdNmeg7PCcnzgD76dGvWWEasIxZ21QzNumWHvOKnvMYtL56N
SrwWNChj6oUzbYGV4YyFVget8AtX9S4ksluaapJ7CHwC5BnlGnqDSjw5+66FrFskfRAC8TNaxuLF
yx9rAkcurIg8CS6PiyQSOIUY1xfKjPD4J5GUJJrK95raSqWuOu3aD8PhnkmW3jBNWI3B7b2S+BJ2
mg9YsZPiJYcMiQoq+pknJJFCfawxdJwBVttinWH0+38Zvsi3w8lXwJYvmpqAjYjS0mzTMG107Kk5
afuUKXuJ95gOhrRcWywnDi/GJEF9MliyaIOXD7xJkTkaqeE8oocOGPrJr+aIx5eKRHknAqUjbQhI
+Md5PlP+G84fZrMSl0PxmNFsccbCLRF73l24auOpVUZFXgPmXJPY30VKw+uDHEj8O4CJiXFruysh
DAXs1yskHqLf8lCHf2323b3cUyx5H8gzJFDhU5UiJoZVPet6kYfIb3FyefDg1vbHGg9nSqHOTBMg
7NfJEQLOqwRYKD6Sr0KVjX3Euj6Vg5AfIa0+Jyo0I628qGeWlN6QKgA4Ra9crkHLA0cstQZWPCZa
D12BpNwNLeB/mzm0UbYUvwqXwbOouqZeUTE2AiCDGU9M3oa1WL/kq+9KuVjv8heA9WtvOCLsLOW0
ZLxAUMpjVTu2BqVLmEMgWCs/qvIOeHfzjeZV6SfuACWxCL+naJgNwsbT6x5GUdxiW/B5pubOodb3
WrjYE66aAiQNpAo8yw4h2jrs6gRgwZ5DqEak3gkIkIVtr6NPhnts4GT456hiBVnC+obs8g78bNwV
ALGaMFAMtS0jooCXlixcnSLhu9s6okOEHXYr1L2zUXNdDrzPl2Z6lfPt6oX3SQZXGKbnVUqwdXT/
MwIipiGExWPGhtktOX6mtslGShvn9So0xCYkIQhAogjf+nC5YVwgvC5dqgz1Ya7buA5IBxZasaYa
Iu6FNoDqo1PAwDJEGhZiElDV6qMPFuGraX7CSms/IdeY5eERrm1FHKhNzz7tfIZdJY3jZBVJyVeC
WDGQJdoPZKMGfZVgeNqtLF1+y6ajqIKnpUPFk3bcU63ZFWuhlOkzIqFC/i23Tv3eksQ6fVODVgo1
NdLSXuLH0V9MN0AH5NNx6KIpyVMsRmrYKIoxXyaurf6Oi3sI7t3P+gek2Ho+5dZlfk8xB9IicXKu
E50A/2fBOoI0VuU9IuNItbB4DgLaD8W5CRjIsjJ+Wmrl1Ktu0V/RCsbQ9q3bmt66n8KBY3QK/8EC
0WChvtj34fzmKffRXLo4+NlJ4/S7ZEps6O9r25OCq/GoS0ufVS/bkUuvKOYAbezAowsxyVMwcym+
xdJemWv07KkUrmuQsjLu3dnfnRNXE+kr71KNzJgmiKWwtNaLNFwSO/3ZLb25Q9UO73rA4gAAfU/Z
VuQMMCOYkTeWqc55Ov52t2YE8psCm6Bpsv9QGjJfYP6j3bxeCJTkZFLq6ABPoNJJeA+Ink8IDwK+
VkeQ0mRKRivWqP6p2KNC2HIttNKwBcsxtPrxHfkaAHpgWcM4Rkc6W2JLNfnpc0XAS1RmKyItGBMj
xgekOtKDRHnVh9/Fl8fkCiL2xY9L+kL7d8VdlRmPZu2QcyePkSkrgL/0BjMVysatiyrl3kgbZsKU
BIlg3AKLp+z+H8mQt3+WZ2TQf+DZBg9Fw2/Qm0LWrIxVWVEwBijYOGWn7v+A2iRtt3PQSvB72xEp
GUJxySQRUlbLiBRNpXEWzVtnqfbamsv0nyhRJNWWHMhBsN9YGpee4i8YDUhJbRDFYfZP1Vbm/UGk
Wxpda9pPS5Mmcer4CsM64sDLHVlR8R+XiJMQ9zqbjbtJMEzlOOb0tvKYI9qI1fT2Xgnihvqd7NAz
SKUWjwGbmtaGwHCy8FEyaDx35tQW/l6xEClg5lLRAlkrgJ9AqRKMDI2tY0k8OK5+pPlsc0/ZwJW1
TgdL+xYo+URvPa+WzZ306Uh6Osu8Re2DxyW7t2VjqfySXrjNqUj+S8fbE5FrZpzvLttxJfamNmO5
pe/HBPjjXcJr9YqdUOKb4z4HJcIVJ9D8XjTkBAe8vn11R/Abpt8ZweSuWB56E6YlYeX3YBz/4GSG
88owienV/zO95viP39vnMA6YZGpFa09xsA3PTXEdLKlbW2vztKC3hl1PIhGGCXUl7rqPUARQYqRu
oedIYJnBVk4sHeHBC4jq7jb6mDirdQmgR6lH9N/odyqJdX8aJ6lqYxVTLR74D3wEdD1+SPOSd6t9
Hycu56otCuP3K/wHioX3VG97wBOIzOl08LUQ2MSjww612TF0OEZWdxJuVc7OhqyWnE7ukuMg6V2T
Y7DtlGflyJHnCbLEVP2gZZQYD4PbdfdlNdtDHef2MhgYiyghaDp1IDv9TMvO6pxbiRiX0UHwzvYb
eD3G2pAvDLAFI10AaQAWgFt1p3k7CujrafTU56tEEz9IuKCMV+hA3XAJUIGy5mnO5H2F+hqRIJ5D
lnu3TnyV45LBZ1pt7jZcmXcYnlkzuVedn6TWeREv97vTm7wVdbxtCXKaxm8eQndzmZDhjm289rU7
2yr56Q/lGzFXY8HNDQawpUhRCD34pRUavVb3JBHEwi7JIEC5lgFxEd05sb/QjThVcvKi/jiUspps
W9Ujlh4obSNUDNzrOXf4nbiZBuozYSn46ZZQwloXahDrb/JRqpFJOU4992RQ8p7DG5Ty4qMas9mH
+Z3c7cbywGMVjcZtWfP/o1dR3DuCnzdbSZD8sFcHaKlbFwb94WZGSBezTZrcuvnwEKHv8Kj8K3SA
PxC0Pzfdn87VXO9cgGax40OysWn5qT1po1KVTW1ybQ4bSYVckrtFq+1EUY4W0g4RC0f7EjYnzeiq
x2AMnAFLhB/CldUSEVJhL9T45iRlQN+sbw32ECfreSFvAb22sT/V+8uRBN56QDk17XTC4UQ1zfjW
X0AYTljIzDSUue05BzKEglUfkB1oy+d3Azsm3sLblZNHGwVk9MHLDjIwiARl6UpgtsPGbVNAHyTr
3vFhZx79rg0nnQ09wEPjwDSaL9Om16lVXqNaVI4A6rPB6s6fQvscFVz/Cc+ZuejbSiYFd1c9xFbC
TNaOB3B0LBWi/ELDnBtMoeehu9Uzwu7I+4Rsqaum3NNoHoA9InrhbWvUTK+4d3oSs99a41F1j0Us
KX5QqBBmyzNV9cOdHb5QTKKJSaIspkHELsgKXVSAEXhn/CTlNmwkNDkTlO8wbxKqFYyX//mam674
W4/4qU0/WBSarZYJwUoTnprhIjhITaLtE6gXQsj+AktKDmxEmtHDJI3aSrQ/LsuUXZ4LC+5iLf7T
llrOUs2dJcpgMUza6O6L/nZ6ESJLc4PeVXzTbuKBMSuAdd/X+tNgg1tViTSEtU+bNxqLsMzgxOwb
Q18TA2dWXjOWytQl8U3fqAeKYUkERo6W4017IM2RG9Ia2nz3765O9Bhup9uZpsPExwO2DtJSqTUl
S5nhKrKxmAsKQ4l05uzHGQP0adBKEnp/7MrbVnG1eC2Hk908Ij1JdMFfEyhG7HYQrwAnvGtAJX3u
WLhjbbE8o1dBMIfGQb2dWGpnH8iQuIBtyGDo3O2mtL1uNAhmtJSBiiLribLLF5EGDt3Ts2wm8q7Q
VcVC2waWpt54yZrwOmV0/G3TFajjjoSsWaPXIy3KJfyu8omyKR2DHaYexrhaZEEtX5V6gru4fKAC
Y0x+37k+HCZOrGJdgki0u5WFmqwLDnlIXfmuj1K6rWjPAr3DXCChFM1aYnIrmqi+fiPjXOPHH2tu
5zrEQ4hOBk24tVOPoKRArDnfYcO/UY5yioBG3KM8DoHwto7BXUVGLCs2y+Espq4z4IqpWAxhoc8k
93giPDMkNyc0u6MCnVSpOqy1GncvJCvJ8qka5YMfiUcR6QYnEEXqKFi8NMR3P/GvyHBy5PED5vSW
hlEoaiPrOWcIbywpn2ZA+x+sYDMafI4BVf9sM3OgWeXLV2K1N7MePK4NQtxZt03mJFyCB8TnuKXU
hjyHr83Wx0fB36UNDaH4Po7RdOAOOshAzg2RRIEdXjrRSr3DPbihh5JYVZGIRJ2T/Oj80Sd5wV6h
RkiIVbw5eVv6bTiqwW7FbEirTw7k00LaDFkeHVyauUbz3FpYYue5SAma+aLSDzC9Zl2ftP49PDVk
dlCFe7f2gTVXRUZTDS0DnTXslWAUaXcirjUYpVCww9h2sZBylglBo7GijFmGH6/s1VYgyiJusO+2
BelDyDnqJyT0U8rBWCUoCOA8sdbhtVQSst31Fa12A0bkydAM9Ww+PUQgT3pHHmOL3sW0R9Pj3hOV
wFbPb/lBV2cQpbLqyaWmZm1WzWHK19I+4YEEB5hslAewncc6N7ZtsxkcV+JK/g0A8AqETrKNeCHc
w9UVB/3ewgDJYqMH3EjFhrPmDquvcC9nj96Rd3peZpi0JjjjYpSvBXHoLMKqzZJSLE3Pf44CWO9O
lyy43y5LSOcDbLgCWB+TES8s3dzNTWHSucSdvQacuncn/Ie8O30NPPfjttB92i3yB8A3CzsHw7zO
J03lUohib72O4RCVq0MITcPhAwJ6MmtnUNI6klx0WH+T8+4FH9lwlkPVR+Zz2l//aszjVoOKmLCK
q+129v9XJ1Kl38SvxOLpevz1ubfeMYv9vTVL99AoRAVGSusLZAqnaPuektqQ1YkspbiA+E0J5h4P
50/g4x2XuMrfC9nio2oHP/HOh+xJkvEA0h8VH2y5Mh/spBHtlnWJ19qyUib2meNLtY8n3dKH05OQ
uY7nxfbFMdF3SBHyjP+JgNz2GgPdn9xZfgg0tbGRzzm3uLDAms89O/lVi1DENRCWgFwJyIx/T1Y/
CWi1whlkU+J8v10CBKgqEhmOSLp7IgVi5Y1/pKezfdz2Hsl4CFjz5gMIKDMWPSQg151FHWwcw3/D
iPmuP4XVFuZ9aYWFDgxg8fsAmXp2SD9Wq0LI2VHFDrGRAk4Gk0crwxaqHjZMIoVyFSHEWTWUCxP6
wSIzfXpIlni7qv0ygmCAFyH/v4RBX2ectq8AZvvnZw1uhWKetPmfq+7Tx0idXqEX80ROYwlq4bly
JSLRMMKkHXtsR7kF9O0QWwbFG+8bqAIo+9HZVRgFMqTeGUlUlvTsL5bHPPmaUCn4pPX0bowtJp81
xEsx/WaWX0uARe2iVOtK4XfGwV6rAai7GZ1je4cpaxvL6f7z6MSgogVHUlEXSrAmVAuj/CZqkLYc
pOD634g6BA5oxSa6oz2PJSzh1CBFPq0/49DvbisRV/DMAfxBw6aLS6OtL6MLCkfhsUiVaewIZhe5
IYbycQhjo1G8Bh5vQkOFJSyE0ZKjHn4kKc+D1J8UHKc7A3XOYNQ6o4nFVWh31SfeVo4hSgnEkQ09
9SQbjH5iAoCeDB+d3SidBR8BGpF5N8k8lNbVRNragDJ24Bu5woZ4TvgSuevJc2BwDAWvKLJv8VQj
EYfQYgD6I4QfuwXeja34YX0x0hTMEhqGjNaoAX/GilqthWCz+ODqcMLtwTpOe4FhLZ28ldK65p8a
Vmdt3T+FU0h7nbtAF1pgWLijFsB7aPxb+5HaegN7MHLwzqhNGwhKg+F5VZrQORbAkbaJOdMzMEPP
m3Oz5TpCC5Tg7/GW91vBaYjtN7vt6IAq0WCX5fN0AcAm0bI0NbDxFKCuoZKLGt3DV7D6N4XvYXbV
fP14vvR6myZhFYej1/HRKTG4qVpesVegsXQCu2HcTgxT1jSItujYvCwAEA++ox88CPZbWRY+M416
ZXvsjlpyVxw0T7ZIcgYlR8DW1iuJWR5UQ4mpUHKwxDd/eLLmOEUysv4p8RDduajipRz2TtBd8d7q
RjtqwNEZ1guQjuvracektBYETiMfnyAJ994v3uUL5Sb9D6nU5xdpEf1LY5P84ETex1iGm/lh/OXr
RNFwOhSFw0SuLiBhY1+j6JUU9re5clrYdYc1Y5jEQ0g2Hs80IjQdffUDXynR1e537ydPN+DJg0Dq
papIubP/WhljC+m7ab02vveQrKhInwn+Kt4IWTxuNPGHmzuNXnr6iJrXdyMzbE5qJ3L9oqhtvjfH
/LuoeKrAUL2X5JtdJ73ZSuGoWFwVdAQhbYoF+qpJwulZ+CiT7GZXzjT3drqugLb5Iqr7Fwxg8YN8
iShkDURTWF+7OtuHwTkZKF78JFIKxqBJUIPzCpSXwbB0N1y9iqBQCkEHJAfXBnfxaXFzJfhZSFTk
R0TBszBNQYg2g0bXIn/n4p9i4vwHv9FSh95+EKwg5kRm2cI3mUYYydUYXs0yI+GdXHaSwHjQnjwI
Dj9VPAn9KBsZT2IvibFTQfqc1KvpHEAmxfwKGX8OTIZIz+fEp+M8ohojS2LgZnEnpd8+i74SlMtV
hHRZcwcp21zcIxuy2txU8D0ueok2tT/LnRzNYgK1cpCEP6+wEx0ia5L5lf5Oa53Hc6A4ywm6eZK5
bZUaB0YopkTl6m6i0PZfDtVbOUKknVyudXAnuVyuCb5RyKGUvHcuIC90fPmB5QcNTQJPJ3ZGrbZy
ZgliMKFPtzPvc8jhucTkO/IiQeBTJPKUKIk5NBbUpXmnLphBqq8S4mG+McS/5enGxVnObKw9VoaU
Lfoho5GZgOjJCMMEZne7uHm1BS9JyjWVl3KlcR+qX457YhzNr1TxO7LJEZjwGq4pmByGBIItkLHQ
Wo60e8hatb9xzUfUfgHk6B4onE187gbq5RQsTV1m3Fgy/U2AsaqJYdR3fW0ddEIZwLvP6Cpr6Sjp
F9Z7lPR+PX96ekFsvBk/Os+eNyjxzayoYGrvoS2AOiasFAyW+yXG1YrgrRRsymPm3tmvi/jNVtlq
cQ92dFo9ZEyKWN71gezLwLs+fhcsHpKUBD27z0WgkGSAeGZewv6wr73usYnE4PxiDz8nM2QmQiXt
FiA7TxpAU89ffAI/g+rbSpZo0QNsXs50Y7IbhwKPpNu/sFr0kF3sc8TN/2uq3lrC0BbQeX8krgEp
pbDJaRJ7gzzNQ3pDsSeM1GWfaGOPiI4Qr2uTqN7k8XEAl3ZxFk1bn0bkBbrgwXXyDhZEpihCcZ0+
C3WSVzHreV6NeWywHakSX6gqumConB481A2rh8YjkS4kOaGsbJ54OfaZNnQ+eW2de954HlZ54fpu
DVYR7D21ZwjajT8QV6wPWUPkvJ5gyKUGmUNnBbAxGx3lkRiRf+4TP/xQKmnC+HDtlJ2Yh+ETY5vv
mcgcusd3Bm6bUypX0vIsDJjELp67PvrD0PXSBYh7noCpCLY9qQVt5Z08A0nGk30WBukNvXIMVOrr
19T9ct7hCs6giRalc9LjJyPpxXKA36Ubah3ERlSgPQFurwej9Zp5N0zrD7AVAvrnGO+xRYRIb8vQ
pKtTc3g+kJ97bnNXznv5VbUUnHEQRUxIRXY43zEG1guhZpYnS8hZbCWdZH/8BEaxy1zz76qXGYOl
q8dre4FEyuQlHiTFh4PhhKHfW7RNeQIaAQBew92Ed+YJGje7MYHITHactkBjfHftgj2zZHzvRWrQ
weWKNUCmGCiDT+8yPQYvw4eFJ2bZs1dXgIwUNT4HKn/NL+y8dYpeR44G3AyOsNN0Ghuq2PeczDew
3gWzN2DD02tKaRY1tcBRnGLkJ+CZAUqmlXSHxtnPDReUK8lTD1nER2fXxv5LQjfNYF+js+yWEMpF
fJsx8iFQ0nhCHpL8JCoH654L+c+iUejliuLccbAHQJStH8A/tSRXWHjq3AQjl+JxfTkfY+QRbrjl
GCl3spqZ7j/wjKKWNXMkCoh8+GKOcw4NtOXQRHZbEqnnF/SzvfpxQxqC78M1bacO7EdnnfcKDVOq
dLc/YV7ZXlYUjMRLAippCfINl1cUrSE6hkHsXOZRvQmE/mx5NA3yd+JrDa2Cm6gx077dfVgJjFni
Lx18dPihTfGtIw24XSGBgDFXDxz6/mJv7Yrrl+0+B2P7yXxXhyA4gZeEEOyI4BtSWTsAjgQFzJGb
hjFBzRt8rgafKxZmn3jhHqIC+8VKJyzo+Dot+3FMgi5ql7kbQsnEA4r8itg58kilcIqoB/SaJRdf
5+IYVlSFOR/M5EgXtE0+DGhPJt3lWzqR1KfBHChvxCHZJfmlECoO0DjvzQCA8aHTEqdguQAuXaZW
D+cg2KA5HEEMS1e6qD9JU92KA1vnmWsIzm+cKbHwxckgMsD3AsLKccPHK8aYB53KeOVmrk0Vx1js
UKwK0E/5nyF6/CRvNLFOgOGGC2kOXzGlCws+ECtQeyPmaBhCqhJYAJ2Rb0mJ3ox4NMgkSLOIrjT1
NgXRQROTR3jMpzxj8SPfj67DRDzCqOG8jGpIGi4o7TTyyH8WDogpr9LlXYNIEt57nz5LFsjk85U2
GZkCGFQoXOsxh31yNNj+mbTKTcOcJ5hiA115z29Pqzx1B66aHI7bKeMNvKaESiZs/B34AiMwflw0
mmxdldd/Ni9uXVELNXoSG/8zZexzPa86BkwlA7o4NXlYm0Sp0C+inc7fpKIchHDCPOb+BYKmfEEh
4fkpaOxePJgnsfjeHSVhjQ+Bze1vIN4h1W5rQMQEl0aucFp5L7P9/egui7jetAbPywmz7xavCVRC
LJTsgyTCeEnp7d9mR9LeD8s2QCgHeOASGM/GoY5xKGy4l4GfriuUSECc8TqSE9hTVb6vKK6Bw7SC
GnM5izu7TlWh3xmrvvaN4ycbZLtAwOLP7tO9BJTGOWcyPC9xh23/tJ1TC62MeGGEvsKb/9ClG4A3
rcc1iNJVU357iyOy1q3S1YFM1XdWCGt/UFXoIbvp06ke6VhYTOqJaZvDH+/8N6UJ1OY04usJIYrU
ximF07VBCQZJbdx5aeRxbhPbtbzfnULYwCn6FEnvfL2UxdpOUanMQNdHy0GASagGC9a+fyPOyt+N
Z/2lPKioxtyBqT+godGa6V4r8Cb78Hov1xphL+EFXBDEoqNKNdkMJVY3JIeRTKAmysbrB79nJozR
6GmRGkbJRXV5PW+AGNBB6aqiQorjHURBuPoyMtRM29806N91grssVFslI72CUblzyWAMCNXopmjz
qgZNpPoE1szG9oXBBOgNMswMUwheOiyCVjsy7GKfPSGJjOUUzIZ6caBwSRXh/AdfOWGH1wqwbGlf
/W+XuY21I97/Lagbl/BdMs6rEdKynFTNcAk0Syy5rtWc4qUA5+BSXtP5TqaY9kR+DZU3cRfEPJNW
5u1hBmhOoWwibhwnujAKgtWVj4uEkWmYcnWF4CE0w7GDM1tLVoPoKE6R5FeiLnDmU8yWOCK0z6yq
7hom31Ojq2kDzTUAkE+aeKGJzIUq0iG1qJ52Zhg1x2snAbauvjH2dGKXBj5GhnU1yjG/9YIo2wAq
bGvGM9iiaB4ExrbXJvCBEX4OIz+AHtQWCavfP5gjM008qPGOSf012Y2ZsR3Xvtr0DXMnS1v+EmIj
NyBMNXgl8jRkvGQoTwQLXUCIwgpmM6EgTvMMOW3nD7Yy4QK8CwLx3Ge0yE8ihWq0qh869IXBGT3g
IdV1R6JR0aedD+wvFmbRRBlwG2aXugSxDLNC9jd7KymCEvdXcVdEn2ujYnGqlf/VcDcpFZdyiLFe
QJ96G3JJ5M5Px5BLZRzMSi37NgIzQ8FP3pIx0ktpllMn7Cm6GlhRVrJz1n35uF+QA7lVE0UQBQBQ
ImAU/58NcInyV9kMT2n375iNLF3rz4eGLlPtOz0xO68WhSgGP1wcGT1Xv2ZiYRlpmffcFBNZ4FIZ
9yrEjrFKE5LcG9vx3MbQbZXxTI8LiLcDJ1u/9e1ixE3ocLhF10GG4wOs7/ADNlW+zPuVKQ2WYfDG
Klh6ldjo7M9K65zgqVPfBZo6tusx0lCJuwjOQ4sVFEZot9zWSf0A5newMCPJYUggegx9lbC9slZT
c0QcMhx1C+5+zWkB4w/feNigX0YgJKMXmhLEJNZ7LFQ8RWtImx/bj4m+3t9YUi+sOnfR78auGtxz
RWFvGg4L+sWV0XNabKGxW684QcXwHcTp+28BkfMlRanOcIsl3xvV3/bol8KQmTbjKI/GCaB+IuZZ
sp2qrI8n1h1PAoHiTiSWUnBX3jVllhm2fJoF4POcaj0iU6CGkR8W6Hmsp4WCZkWAHbQ+CZFTpsa2
zAgRhLQOxky00+QBvQ0Gjw8JzecXgZ51BzsGEoSKqIw1Hqw5bWwhH44xxPWLjvxOwmFFVyn17YY4
KOqlEbIPGcSlh0hrQM2FMwjknPDfHgDoNOkwOuWfR5YJXRclOh4SIEk0RkVY8WFurChsswWT7ZUS
NaQMq7zSQwJGhpYW6SM4xvLaMK/mxWE/7rn30WdBOiJ4N6PS5cXvdIM8tP9OfaadHPTJ+5w6YpRh
4BoOmvr7+jV7UFjP60BMdHzDIYzY/IvUPoXAdDg31lKWBQrg7pY19B9aLQRI28N3q1yW1hWnaUEN
kOf3dm7yiytQFwL2rGwHjVRelXzreAhFctZx6DcI15Rj8/BjBQNTQKDQqdNMm2LZOtR/jyHzAcPB
02yD1ctoOsuJrihJRJpOXLofFHmPVx86jSYYszZUC0LUqG3fzQE8CwJ7gp5LNLv8IBgXCD4Bdyjn
qx/ISqb42XmSy9vhaNJGUQvd7SndktoY1hUZfe/I/GZNsM3ErORBYYe4tNp3WRrmmZLiC9Pr72Nl
cZf1fORMUpl/hTlw6cD93lzs3Br5l1WtUXg6laGoOaYS8u3uB++FsKS/qlfMZrweyUxhEA+vvzak
kNJxmKyTYQD0zZzj3ZWFxNs/OIxkjZ7LRa+tVSNN9QctoYeHde5M7MgTvWncc4aEnxPqh1xRW5en
uTTyEJTF0AFIhdmNXy2bCUj9CwCwNP2aIQAdI6durAcA6lcdPKs5h8OO2AxpyVIBwB54qOKx3kCn
xut4Voxd3SIbSS83wXFkk79EPH0ak5VTpVOREdmFhLJHI/aBUmF7bOULDdNlRwEix9vEhioUpmEh
CQJBowt7zVGA+6zXOgbA2l90Rows5l9Ww81vXQVYe8WmMb0YsD+VEoBtMicgwXpK0TL3Mv9QIFH7
POi/u16sD4JJS9OZxPetNOJepuEC1CVo5hSvnwf2a0fvyLOuFjMpEVmJuCdiPb1UnHlasR0CRs0T
IRbWFcd9EH3MfnqQuhQGI/BMeq8CokYJ6GIgqHMY0lthaGMk2+PTXdVjiZpoH5IRqCpGx2QewhZ4
WdCI65LBtG8rHKC/UuWjCWXHkhVAog0tOlpvCh9H5/Oj++P3RHcUCOEu9YcyfwaG3uWnUKrfNPdQ
ZlOWRzo12mJCjzmMKST/d3yTBUPXMp24BspoGOk7uZyLXhOrkG0SyiXDIyHVCCvjzEEaXvsDjJbb
YGgWDm80Ia0cGxAug4dAfYfWNhdJ3I4MMbEyw78wFj80odSdo3O36mG951Y5Jd5iKUch+fN9gVtm
E7TZot2zV3mqY58cGDSTsrJX2Vo1UFxFvQzNR6qg72qPjclJNztUH8pnguAuc8YzxjJe1wUZhiou
oy0v4OGLXMH9H5pNQquFWNwcq+GrL52fGsxzkI6ssDZuIAif4GoZPHDnYl2FtRUEjEHw4d9cLv5s
6M7trHokZNYygwbFPrK4GKU/PBgLezINZVh7dg7saSH/wxJo72VUK4n7Rl9uYMuiZpR4wwlaqNmV
XOVv36XC1YOHOJ7QPPHE8yssyuM7ciMeVqTwL6isY6Yx9UczgUFzFkE0MJfl2LnolcQAFdjbnHoq
ykJxg2Aa3ZFDuLLCJDecdDS8VTbaDShuKR/Tmf4iFf+TbdjmKiEow3AMlKMlsKEEXOMHveBBmjlX
+7RBXl1PMR9hdZrrF9nThasehN+cdnU9b9VSGCoNj65rrCglg42Y11OeS2vDSToHCKH8gLbXCqeg
hrLFFknMH1CocErFldXCT60sdeZ+4TKTt3qvRi9L4lmcEcjDPaa03cocwqPR3nrGsSW/bL7PoSJ0
KCncjhD43KyMZ6QiCRj16n9KnLIRGEWJzJvz9NFgJktMZ8/gK+BwTbPJ7XdqSvfxcoVSDRj7TR4X
19mNm1L/di9eYoAJJoEZFktyg3zAaksrORULVdRSjFnYBCojLr75QQOh6MWTf6oMk4tXpfcXJCce
dJ9gKLHSvKjMm+ShZiYyrv/4zBLpakv82dtGqYtw5ppXsmbrylzbdr+L1XblpVMkgoPMqY3jbPJi
i8ZT82I4YvXZhN1FIyNyfAn0SqNtYvwVJBAoLki6L30g+ROZ6hchIUol0k/5H8xYWR0LgS73uNWD
RPn7UYK/A+kvfdzPs6HLvmUd9m9ZDB8nNQ43jGF3nAyL2LkrbZNJKejIh6cUOFf7/l6wFDvA4Jj/
LqhOsFOJBYVwCU0Vb5hcZgEIJ6Y7/KuGgiAC0a8vMlik5I9BJqFIv8YVAQdgUI7jOF0htH95s2ZK
AF3PlzSvf2TE1b2ns2kQk3yPfHoWWd/NJGJJ4Bb2PXjMk01jj1N0ki9B+6Tnl7/r4l6BNrvg0Ijb
Ti0KjRSQ66o1G/bqKqjrPaGD/KaG7pwaQ2LGOUjDm56f7xMSf3cKoUavrfzI96ZU3rRsu0H63+nq
wbND0eSIt3Y8mUMv8p5zlXfiiSEwjPG6G4vK5C7wbydPN9SZn5Ybbfa4OocdycF1ppcV19N6tgIP
kJQomrWfADVTVVLWEZk8KtBTpgoU0AYsIRllPJMbdNZwVoyvYMLgUmvqpNr0o8KpVfktvxsyOx85
mhRQtYPW016d8Tf68QCsf+8nISQiy+RmCXb0IN2MH+7tBOO8HY7LQFqioKDjs8E09pPjxnqgP1Tk
qOc4GN9m0iZQykgKmh2UjKu4N/otF9Rceh1RmMvkbsKU3CEbN1s+qtn6opo1vciZ3915+SFr64yC
eCXKzVNurXDmE6Az68FI8Tb4gaSy3wUxAjbbs0o4ZuaIEuyix91epFtmRXiPX/LNxUyFFc9mowX1
kda+GcX5bSuAp4fNEqLoeD9BIMG/7pZoLLhbvagcSYTlyyHuvU/9uV35TSuWg8t2AMKfWzZ8hVNJ
Lu9EaIYYgJ51/zKrUtAY3p/NQCm4XvhxuZnpkp38Aif/9+LxrH+bWM8QiI/ACs1O7GRwHYV286SK
OOIi1VLEBx0EyL5mq2jZazs0ccHL7YgLkFmAgY+eIOO9FJBHl4VCUAKnCFuhP9yUkn4p26HA+pH/
fHzK3KSOauYjXaQPYq9kozE4FB4pDeVFvIUN7JxbDU78UfOGym4X/A8cgOTtbb4t7zGWUCiVckls
KlUPba9s3erfTUkyah5yue7c4W6N2ZLvgb8O5eOqOScml3aSWZ5HLXKTJggJnJpd5qfFXf8wsPc5
ouy86flRJZVy/U6jLmlI1oGgjPXgORsw8BiyrBpgKpLDh7yQmNuiGai4PAB8JeVgTxJVRW1NyjCb
p3AARo4zm2UbneHM9X84H7ebRg4MTlipK5GrmMDUcC66rDs4kH7p5oqS5Kihtf0JGvXhjw2Xkzah
/Z9Y5TcoR409WM8rhtMItJGgug0LKChnyRJXqTKSm6dfj+Jn0/52m6FNrcYG4Tky95ZPTcTfN5US
n3Re2uM1ulTAj2MXBgF28j1rUE2V2sANrDWdag3P8RG5JCIGGuDAOkdYWC2aDg7VvIyXA6xwvhNM
fAZnF3756LPiwiu61jRp3CTCYViMWFw/sKZ3Xl1BMGwGqFbiiP2lDqm5SIJI9JNcOcxHxC7UDTWA
tsIrR0CuM/DKa79UB5HA0DEGjqAUHL4WeueKV4tgzbCeNoAklwGRv2s4By0gRP6QV4JBF8lwsUmG
RsCUzkUqImLF7U5sKW4r4Fm6ob2dgEhd61+YaH0aN0UixLcfVPAGXEShH64K0sYLYOHzydq35e3a
yZ/SiGfxe3gBrGjTfy/s9C1rLdetjKUsOm7PoEk4re2+z/jRiFOg6KxPhUfTwWm6UBx5agPfIT3s
Cf7fbLMWPC6HvNak4CYigUXeGv1/83AdPQtTwI67b8WqllNWH+6ZVrRHcO3XRzIEYVQ1kdQ+Tnp1
L5+/vkxCd/WYLsXPs9ZSmxg+5f+FbMg7dPGpt+r4Om1ggP8K82ejpOkF+F/vRjmM6C74TcsYCpoc
ZkMDPB8Mu86lv7zDK6zD6a9NHZmneRrBJ2un9H3isCP24XyTc4x5KIFhOrx0VTGB14AfzGTIDwez
vaPiydPpHP1TWJbdzrt39+CcOq3Np9to0hVJLmDe/Iym575x5iPnP4t+mA0DbQLO/Fkx2cvSeeRx
fGTrWkKBmM7QPyChU8gnZNmZmO5ulEndRhEEb/qE4UQ44NcCbTSqoXrPzXvUZEpuA1Le+Yj+6TBY
mKbsHna4o0N2LZHwK6BbIB5WA4JPYlgHr1pcHghdQMzQLcCldApbLab1pWz5anGvaxMDld6WrDkz
xpWQSAsXgLAsh9xQu2lRtx0du+kcrbUZFmjcSL8SyzsGIBf7dMdxP3HkIq6H718L2sT1/95wIkyD
Kly1cg8PUjv2esoxgfU7rUHuJS0hqpCLn5KrphNnvwq+2sbIDoFsD9HrSIcOVA5QeaQGtym+axCx
e8TQPvqUey0i8dyu7RkXYCxzWX8Az3TBtx2oUUg17O/yhncWbOyYUiNyCDSDqh1MfbAAjtPUWlRw
gpqON0c2sg0NVfTY9wqLYB14Tb7pMkF8bw3Yytfh7JUNOgNB3P/D3TOeYdFjpGCZAseSa6bWDdLt
Phg9msQzwBzys/a4gtaJ8mkTtQLC3b81qNExr69XZ2Ue8s9poFS5bNvfmjQsdNRpabEELfGNYIgo
hr/6QMRoQqUDWXAFRf+MsbWtWlL/w6+nWlakOECJUUqs3fHwaw1ZzbjHwBlkmVDXhG4jYbyxPZkc
qahMhwUMcqV61EygYZfzKwjnWvsOnXcjTLZqW2syzFoMW4CoRm1xPRcgirZ/Oq/9KVJJAOqB/GPX
YVDzyd+V9DxR9RSwDMnve6xfNaEdBn3DTUs0IiMYGK0I/AVW7yucV9Iw0jUK8BrRff8dwo4Gk7+f
RTIlWwmFf6d9DStDO3MuBMf8W0GLBfvNyDTZCgc4GNVGqVU/zosd+vArAToQOi3voaNKmow9Z7e7
RL/w1SMctRCtBwwacHtm1Jv7PX7W1dDd1ZDYCEV/8CsxyOgunRxm5Wg5cHuGxdwbkDQezNUt3SFV
pTMZwC3f6o5cz6tfeqt2gBgkmZduDpzt/sUqSK7vulMjmZCu9/2CB2Sf9aaOjYNJAgof/DW3gmfW
9A5gRAnau3w5xeS+xwJDKL9IzwS+ZCKr/ENFdyf5pqx+jt3sbzMx0iql+US+bcmVUM9JQHZ12jBM
WzutBmZV0dUOHWSd752VQv6W1yB7QUXRL/FqCzLXSOiblI17rMqAhmL12gtT8oRto/15hpWVaIvA
OWvum+MGiDwy6zFHU2IjQ5FDUb+A3uDkjXu/Q9FkUAP5Qu0kA4yDc7Ji+XpZ4j7kJno5UUws1x19
GqUKgsjfhSrcCpZox8iGsHjZsxC34U0cWq3ge1qLqkADBuc6Z5Td5fT3CcoEc5V/BoJ/uD8ZJvBg
2h9FW7v7U+7MjRFHhMSzuEugOX2+/a+32G/0vF6pCq21t2EKD3bjgl/54Am6Yk/ea+gVRRxSPx9o
tV0qstYSrq6gejZ5MTfN58neZ/LYOKpGCRlbriPJGLuP35nW/mS2eh+m9/wQgHeCIslQbrwS43iu
UWR5CyOlGPEudfbuuU0Pa0nRaIGv3KOpKQLXzllNZhO7suMsIXCUdwPU5RWIzkteGcyOCOu4RK2A
sMKvOBR1nDS6fpqKyF21hgz0Nsf+REPWCiEC7QVxIqhRbgR6tHQtxptmxV1dUs8iYG156l/xMDyx
qW2oilkvhdDl1sTk6grQfZhyWjB0z43G6wGsW7xOYcpsATUQCfomPZDV8K9SMPuyrfBB0m4VdH0U
UnPDWVi2qD3o5tb4SpRqnMHHKeQW8g+YttulAHeQCVkcfJZXINdMEHEh3Hoih7Cv381Qr0UWgL/P
rXjmJtsKHQVUY+MNPBk8TST14MpI56+C0guziGQv6QqmBNOAtA0EsMm0C7tybJ71T8/IIXQ16JPq
ZL3MO9Jpsy1jvOr9KYpMwpNUSRwvssoEiFplZ+mwmP02MYk13uswHiLJwFpQwEZJRFcrvU8x0+k6
T/GKRWCYXx4mijHtywGue6p5jER35p83GYeQGT+3oozurzkwifSrWpV2uWvEIRgyBm+kbvH1+jes
R0uu1NCQVCBdKfzLNxunpZZjHCXiUHPavVL2jDEyu2tBK47CXwTGJtNRdBjGzXMedlLI4BTQU6dr
VGdEAhNfLIacw3PuHPe8+K4Tt76tRwXT9gXAeISFRaC/LzIvGjPc+KJVHedjXjlR6Ei7Ouq+6pW1
BA5H98hxHnQtLpc1iEHDwOQmLrnmKqLhKTzPhvN8AeZCzaCLQvU0AWqjYBDSkMyjDZ89kjmhOWNk
VfUBCKQbrctvlZDh71OWd4UroUADIWjsB87HLFfCRo+AhxJpB1zhHEPTqw52L3/7WYUNWOdxYFOd
ewuMJO6wERXHGNJ1hTLk21e6w8vMIA2R2sBvrQ8GmYF97hpWWWCxh77zPrqmixGQHahlORovnm5w
wOaKr1S/pmqMVjcSTeQJXNhGrLk+xHq9ctkAbbgikoeEvZ+KNQAnwiY/D0uWJmOVsgM+J/eWHssy
LT4jZ5SjjmSk1KquOyNHsQjlIUKM+rIv3PMsKdePl26/JQIRu50UU/2jqMqt4jsjJr91lTi01iU+
+Vt8FKCrLy1BjTITWoUFmbpruL8aAWUpmNP5kDW9aZe3ilCppH9uSvst3RJmQvcBOEEYsB9UazOl
9AVpxcqLJoKgxtqETA+rBAjLzJkxM6VoRMPVRopi9fh/e6ak2r+h2wvFNdNfmyu+7TBwuddUde6b
6T/0RqSttOnoN04todRkS7SG23NnmAbznIBO82LDq0BZL+bGNZlG2kKLgohRHd2XBAyl7PBI0p7S
dtqgGnd8BcUcGIpyE+dzsjiLHkgbpt40WoAC7GG5AfWkM5edaZPOG2qh0WnV15X4j2EqG+HocTQv
GT2U2PU+uZsfGh2ruAfFyI7qZ5DXjrv59rSjd+8euLv3KLeJcCBcGfOBcHeeh1pwYCsNdRtnjNkx
rl8F3jDdYvmM0P3nbYlQK8IM0tCLTxdd0QjsVzH0NCF7JJnBbhrSEITeILxHJqykLYsNUNBZqh5i
cZVHNskDiHh0fGZvBflDqzZ0JQ5OTFUCph45RxPjKWunMXqtiOWaNpbxecifyh7GNnYAmo4jA7ns
9p8y/dFmtVynEh3nNSTImrxDBXFar5MvlpXLCmyzM0SNLL6fFJpfmn0Cs7AjchFxGDOmAH15tmrM
jqth5ZWFV1wuO1gRUeUvNvzDmrgj46ZS/CcCcSmq/eAaD/xETbH0iJNItBLCkUwql4BJqwdoT01o
rdjYPhJHl7IHi4N7V15ItTwn8XR8eAO30i8ME4GpMf5ykdoOwUtPYBiHbZVaKD2WsiAgJolTirBw
rYQVpk/XsEYXYtl7XnqE3U2mk7ZU7EvyVT667AZCvOHh3z3pW6sZbaK+d3x69xe2qYVhJdJVzCtp
m11JtcUV1PFBwYBUicS6Kx669UcAcNqULJ2RHJ93V8mSRPQb0b2DRzkogxfQrPR9l+G2pQe5l229
/IcMbwt1TlojcUr3Wpz+gkKB7pWgjlc4chMBEQDN5FehYG1B2Ekl7MNGvBPKahMctK1/bXxDqOD3
gEQJKzt+z9fs7TcUFhDydWTGunlZfA2LDtAhyQFFYChq77Ti3jj54NQUWFkAOoGyQMzuYXSvf3K2
GeR1pNBoW2Ofcw48hZ9d5NRM0b0dOSQ32lhovZBkWPfD8o4yrEhvLVaOT9jv5oOv5J57X6wpv+gY
FhvM+J3ob9Y0ZaB71Z6Y3Msb6lE2USQzQPzzMvr+7lvv84SOgccvFNCMjczXFx4C3iMjpe1ukI1M
S565ipvtfTJMf1taBHNiG1Y1Vr+eFsHpbsyh8WXPTx5+9ijbjoAMwbfCg6XVWQA7SMuqJd4FmjOV
psjiBMhm/ptjNLmeJuszpQt1uopoyc2EnVDc9GkehV2KGDPUWH8u1fxq4ZQ2FK4kHDAvZJ3lLq2S
5akhzacWKypgtVAYP04aq3zI+CnUAI20gE/ZU8yRED3hpVMQqe/ebpTqvmmzwdKZMlaVKIdP1ObS
4nwfBRpsleFe6oRBo4K3U+54Kw+i2B4b2/Xdv89OGSgHJ18nJDjsrEZZ1t/7cX3JUfoZ7Dx0UH67
2g0JZdaWqsn1Hgb2VqddOm75cJV3FM3OzylMqZeezRKNcvspke/QAM4do1NEWY/Yzcx0QoRpGYnW
7runpGoJX5oa6B65YOu354tCUOt5JLYNwXLKK0hhsI879Syydalq16es508RXpJNywg53kiFWyAY
tl7U6t0MxIxAPsiorEnYa3RLz0g7QNbq8uywIRVnfUdsXnrZih/p1ZrYJr+Rt/Ijicf5AC0yLu8P
Ywe4M5pZo361G8iHwDJyYbH1szzZqGNqC6V4+i7bDW+SUbKwHr0WEO4K8sBvzMs7K1eZk1UEqh5Z
rpaL7/hXzZEaw52VUkb4xZitbaUWxDLkkweneBlFqdBp9ZIGUOSvQEqdwypZnqWmde9DcXfZ6vKB
EJnmjx787Ccvyf3t2y02K7R0oKmqH5A9uK2QNbHRLc15QU0pVD8urUoTuapWMYG84s1ds7RJKzBI
gvCxDdJv83BZTQkIQmv2fCJ0DE7lDoQ5MHCIOVDBMwG147sDRjbV+MVuhxMhOWLACtYIoGoE4opd
BcGqWf/Nh5kt2GXL2pHcpm+mao4Jr57vPvdOvoWDrrDrxbXmalA3SbBjWWuZ9OA2LWDy4rSVcqbH
KR5+V3C1FvfPYrHbVtbPk8JPW6LtxHDKgbf0beVxYsdZotwMzOuPjcYVfz//erAa/aS8ftNJEb8U
WPul7OQ25qC2aLNHhipINwW3lwMVEOg1noitR1fl7hTwpy7BL5BbL3PwOqnpLKXBfKV4/bSfn/1O
8h8pCE6V2pLi1qxJ7KBYNaXxUYACQ7JRBotfg4R38E3ryWbo1vRglxRFTWbsymhVkSf+ACTtMijt
+nSxm7GRiebOGQxGQTfxwZWVySCbRphc7lrmp+W1mKEBTKhp65J9bJTn0YqW7v2laJTeZE1bxhDC
M4tzstHNMV1A9XQdhV0iXIMItQ6OOOEXnowKf+y1YKz2OCVyG3JKPWV1UX7LDAy5ctkgCe0umIUj
/2F1liSX7ZfGprJvp0uB4DbR69PwZY1kqnzy+yiBTwDABOVPj1C5izPUq7Z/GBa55kuCr66l1UGa
JW6BHvE3ywvNz7tk5mjOGyr//cQcmsPxJqEU7q/9unwxjU/XDntIxkV9FE/Rpmm4RQIOJwVLY52N
X+ixwRJ1ovRaLJluVe1PYNB2QGhLdOBSnlGat+liF0DQQKgODlIrfmq2EdMxPXUy7mkP6YmdQURA
Id8D5Ovi3kdQbDpAgckczX2+aXlUV49+D7JgUBwdpvvWq4mtVycNbxksUUqN3CQtPZ+ByTZmVH1n
zNGfZBK3vsFNOvPUrFBHgXgp2Ag1qwjBmzVttfJIF6tJzOwyTbUgSRctRveK32PCNXxtA9kFBex7
uWyexLJZzFKNEAIXWkXIIEPpwNBCk70owcvp1cC9VtVW3oGJ/9lwXxwe9pUy3j+FA15wWPQkNpJd
g2mC6ku2pwaYYBkOgoOxbJ97ye0an8qs/xT6Szn8gH+zc/X32JgrrBtJRIZpx5JBTbBy/l2jWkzs
CDHDfsf6ItqPXIFViIqfp2FoegvAv5h+kXAQlhv+cLz2KaRS7BtuMkl17F6UHEYjZduPwajPm/uC
0wjYSv1bOH2TXy43Yex6zQq+Kkx6m2KEAgUdrguTX3tb0a3f2wi4glXF1AQmRts2PfnkBm8q0v2h
TbQywDKr0bJsSkOKwuLqmYJ2cKxBW8zoTZ9Z+OdZfbYRzdKEYS0S4msO8Tcs4vosUYUDRRENwrAZ
k6mFUY3OVHUFVw2GDW6AXmG/LgOCuuvfQv9JDUn31wU05iTKjESD2/EtfQ8cTnUZ78eIVLQ8FGNS
TNL+1q+CelvBQRqNDLhfLga3m7OefvFzCC72Bizv3fiSrl1Kb5qRuSY7lbqucF4Vn9iE4DSmmGiQ
/v0VZrBURV+zZ7mgIsv28dOHxh8CErfy01ZXhshov1Vs4yyAV0bghprtCCSgt/p9QlSgLKmNP6hf
K3w3VkBfVq601uihShx5iUGVb6UWt3X/uxeiySlqCUYpqsqfXEdagzhDZlTZ7iRcAbaY9mXEItq3
L2L9grnCWC17zRXZefIS5uxPLYcugAsmktEycfQLyom0t5YJvBm5D8Qimf3eGNs+j7DpjACHXxas
kwL22eKIJpG1Ln32gsdsc/ATIeuU1JkfVpsPJSMb99CYzReJ4HYg+cvQHAHNa77tBY0Oo4C5/2bA
o61wtwRrj/Y74L1002CG80IoeMPDSgTWR8tQfxngncBhnfDOEaZy0yZnGJiAFhbSldcFBHJ300Ho
2gGHDQyXEgwom03dUdL2luXxXJCMQT9103O+GSgwt1jgNAg8fo08ckbxo25GT7ULSDaFlVTS93Ka
BVr1pnk8SkYuqhZa+VSq44QcqZ94ONKKNuA9R8S77uonza5OKtxQChfvEKlo2iMoGroYFQPB7Ckj
EGUdsfkTn/QyIK8IHEpDvOEeFTBhoVqRcQ/5pKZLY0ytt0Hb1AdSFzYZh6uQQST5MYhIiVyF7nHx
p0swwKpj58AGUHDWZEhW6BpYTEskuPuKaFtBPvc8DjAgSBb9IViq9UBNoHLCVMfgHKOUkncjCgEa
bUxJHEmbHseZ4cqTHnQN9O4ZBX6tgbC8wc80OIjMa9uNz6i/l3o6EciMGaL8iFBJB7JRtsBZE2GY
UPwY1OYzkPKXJ5ONIc2uBKS0981hKGjtVay0LFNgWp/Cte+Lb7v6g1Ip49UndRdpu8J+1QZYRsoJ
DvUrsyHamTXXi8vMkYQ2QXuEUzd2TgvEJ6vb52RSEv2qCZbQ3aki4MebnXi5Rp1lmkhChL0X7/zR
UBcPtYt6+Qmqrk8QhEWSCGsfo5Rbs2sX6VYudh7kiDem5ZVUhV62sCBBnsB9RN/JLSpg3eTlwzJ/
KVujKTMdY03ov9cVo+T1bzaF4IBNDe+a4t3aa28E/cWUIv7XewG+tz6bQLoXZ5LCH6w0EYomNt/I
MzK9FTg3JM0SEZ3B3kL/iEf0PDPmlaFWTz7VUr0S7123w4TuMMLTUj2Q//pjYySMt7MD/rgIoLbx
bcEiHI5DT/jRzx/2fgFu8CFGc7d83tlIOoIuGAjQggCYSbfO7/sjrdzlbFtsmdmMl8DEGtSOg6GQ
DypGss9ILL27A3U8E6gliJC/wvxYxo0omBJpR/BVlKXng1rS7WyY7puakAQNdgsqv70F+5VtAERn
UjJ+/X37+njKU09dRBySo3DJqOFl9Qw+l1R88W/Lt/i87qH1+em5/CjBJPd/0TjdrXsFGIxZgSXM
GPTD3GDDY+coJEu2d1HkhnSS+TWe7VYyGuNxKHugH8rarRPThOkU4IuswgdSoRtKSYcackZHhKhk
lknyKoutXhTJm9/l+W8soAUbDiVtVD5N4J+bN/9fjzrfyf51x4PM8SbfGOP1O4LNYnilYYjJ63Lg
QL/D6wy3elTwEjzQ/8RbEiojKbN/EpHYrKMNeUKhvc+7gd8r1MQ+zH7bBpWXs4Il+jmrlvTxaOsX
v+960MhaMO00nfuF9D4zoYB6chnexsq5OOmcKUXxX8dLhL46u6G4sLPJxlMLACnjjfK66igEJPrd
Uj890ZYUJhT55NTlRuhPlvfUwo4kEXDCbjy25Dl6lhId+CsgSVL53j76zKLdO4k7GIXDFACANSzd
MfX/tJl3NosWf63Z45Mqm4pjdm/XoMNs07uHuEqoNo00nHCaeeBgkVNR7d6/f5AZMvXb9xUWnUBw
UZaVDf5MKuNyqCfl7rnl/OhmurMgQLY5d6D8bZnR4bgNA/GePkLjjhDqMLfKM6BEFuJ3B7JGVegb
kGvziarMkINuq/b9WyzJhCekRyxwB9piQi+K85U85kc6B3bgemiwm4tN+y8hxpi9+OnlHxLn+kQ1
EJN+vPIynGcvxld4k4ihvXAIudrl7MKPXm/G4gSjTorrgWtgMKI1UJhMUI0ZYCx+vJsWyMgoN8pu
3UnPzWthXcUdfSsjar+1SpbfM4c1+66O+gmK5E06GsFB5mhqH0R/2QGoQ++nTZ3bsp4iBCFvpduP
f95CVfJer5vCUkYtFRpcbvXomUMLHMUnsS0+stnSmYeo7prLMXBq9kWEPYgf8JNCgzSYA66IccX5
aDk2+hTMhSXi7BYsCYjUctY3a7pH6RTuG8JwZ9FkNXULhbNp5oXCnPCOmDun0WQJH45JmBkfW5n9
wBCNwfThqaeEVy8sS0ZBkT3R5soSiHBPUhdjpOQfJaEgrk49oivDaTJq9cqzvcA1htPvmMaKgt7N
1rsK/PIUJ554+RnuY6AwxxvS1e6cVP+VP5tGJUtp+ilcEQ1kRwSnh9Jhk4JG0jZl5lhMR9tpqUFA
CszEuhHPOwc3zEEgn7EmLXOIrEnC6x7pUuSCMcAjcUCajohEWauwcqc3ueRHR6xlvYmH1Rx3kTJg
Y/PfcRfxMTDM116H5pQ5p3FLQ9/u7b5XYrdwwRbXArSQd3m9bF+gYtXjghT7zOxv91PaNk5gmkpY
zRKvWBspIMdcRChy7ARRNQqlxy+5zU1OlvHO6oflhH2W9ME4Nijks6iLlmXoWYuY45iH0V3c8eJN
UdcToqaDoas1MeO/pxXr/jgx4li4QhY9ZPV4o+Wv3aLvzNrH4pYAFrKG29qxZ7BqhY54AdSXyfBx
nXfzltFEBe3DpAysMtM8mnAlq5nZrRGtyZN/E/q0/43wZXLgHPMmyvj206+wRG1fRPe2LJtvQ8YR
W3Fl0GhZ5Q4cJb8hx07JdfyNlEc/a07711F4hV6B65audtstvKztezCVOOjPma8AEZN0FXWFIN0f
L90yCv3YjERQCdYoJQAlcx02krlBaxnX0J7f0vpGK/PeB9+VSjNXhHb87mdompxy/j9M2TGWuZDs
m0vWbR4D9s44F5B+5lOYACVP2VipVCcDfdKIKZdn/F/g8qUAAlw9n0gOZhwkgtAR1yQxx6A2ONob
TRLLvSYYTnYNw8mO9eucqzjgAcMiJMLfJt4EqgX61QnX/l5jZ1NWvSem9BxxjeIi4nxARy77VlIV
fDeB+n4tE1deoCbioa+flP8Z/WW0E1PEXOzZWixDs2Czz1VlfM7LMawWRE1WPGCuCzTMA6lpVSCy
ZKFEj3nqoBBeCRlDEZ6l/yGfNgNht9y1C8chs3nHKr9a7AGkHD4fxEIKC+FiKWer90b3IOWwPajr
zxTe52eJrjUln5f1PbhnCh0eGPj20jK27W9mVufN5kCZkkZGqqCCCzp1xykTR2+xK/Moq3EHegg6
iPebU6rjJoRJddg3kKpSLgnF1UGG5g+MnKPkhefSSGDHwT6zQdFzFzdxspe7OBLe83skQkZOQBOp
Tmzb3zuDXApMfv48SWSC9oLAImubWU+PhlbJXcvHy4sKWidntAbYTVpVIg7gJX91pXSKfiWhOmvv
TK45maxhduGQbdGsXJXkaiF0ZhX7v2BD5V/a8fbO+8+6cFdkp65cg5uFGE0a7pB0Rbg41fIbPZUc
2K7lNzK7zcA2684qvaPTJiccnNcvpbLI/y0843dfJi+ZgF+hWCp2uxWdB18DuU+rt+TbNh1pbq1J
hCPJ2tXcR/1kch7CGoWWYIX6oPzeFbRParWleQKeMYNNnS1E+WWEQstzLF0AuHyGL1S2IyYI6nyj
nr//45M/L/PzK9cAwcZA5aXOvdcmg2jIFz987J4mtD59uHecYzlhmf0j7HJKBkq6s10MGCE4M9DN
flnW3t56cXoTAtUvsvfS1i/hLpDSVr6UYprLhX20AB3ERppdXe9zyIYRh24B+cPGqPzUfGLC+Zwq
+UCqvjY2mUj3oEgiNHMNflvHNDsX5z6saRyP4KLgdHbKUAsXcbKpe5SWMyMJcdAWCU2StdS2eFyo
fY7DXL7stlzmLRLz0FclLJxRH6UIJI0d00bGPMe/pxUlOO+MPUuNSdikdNGLqddLCsmtF+aaLjcH
TQqv5OC0W+wKynhIOjh/RmYsNYIru9OGVqqWSdowJgGu3g6Vr5eZcJCQ61Pj7c6XZrPicku6AcTP
DmwoE5iOQ+wl9qcSz2xb4vHUH38BKMymVEE1dajBnKKxHTomEoh9ifsioMBbfMyh1NCS7c5lXT3h
ya9MjKz+n2zz1CuDM4NQ2mSIjtBd83mQscFkoll5scsmWAl0pFGk5wanc3/xXnqq6zttgp1K+Nlx
b+2DH3iu6K9CN19yrarQg/JZACAUFNBcqNaEVaiTGdsuGNn/dgArC0Ov5+MisDA3oFS1JjY8bcJ3
o+Dhl/JNoO/DfvPznSl8scBcZLHVJQZx7rkm1C+OfEFOmbKRPsWDA53EeqCY9UM5+JhRipMiilkZ
SjsPx+3/8zphArY1kV+Rp49AkPx9fXd+AmEd3FLzZcGVmP1/YpWwHeOhAbXRQaXdckROpptwAd65
o8L7wk9thsSEdoRTSVK9bYt1IC8qx9ebrLY5rOaUuFHFsf8hT8bl6gHzy+aLWajyuw1QEbHkRagw
LEih3hLqeVhBBrMxj6TlTGrBah0/U4PO0IDVcmkTICxWCSjcex5+mmAQ7URhLFI56hCd989FWazl
WSq7v+5e4MPFFms3tuB7t34QFZQ3BSApos3Rojda//QZXeAlYDiYhYKsGd9N9ZQvrVfnPGzlMgNf
YdPV0DJA0Ti6EAcftfIEZHPBGmOk9AwGIf+/0+MIhgUU+qTIg/R4eDUrmfb0KaxMmMHRvQOhuS4Z
gxjqJ0nS1FIlMFNC8EyP38+KRG7THM1AYdCqUXeqIuR/ZKORGTf0G5jlbdC06zzB0+LRsteyIfwU
+OSZ44mJX7o+0UD+A44p4uQPV+wcvML/INnFZNad0JnJrZDZUK7oO5aRb668+HWLYGHwFTQt5SrA
5y4j1tYWFtC851/pi1oPVCf9NHlxALSpI4LKzbobcbRsQUJCrN3GzD36RO5OhbbLPHZ7Os69T9uI
dYZZgJjeAQqQCL48POPN0dI7GTuCmGk1XYzvusTo/UfaT8teo4wof2EoJE6uKuOo8Deddw5Ds12F
k8GXR8nAgmZ56o2iUMOi3zytY7musPf4O2FMLMg1OILZTlqERVJRO1wP98tF/IlOhLa8TyF7El9c
51XaZD9hAr7sGcNolqBsYrloBEvpLArDwChjUWdpRLIOjBGnYHdclIUiKkSuirG6oKKJiwVQ5S2Z
rBdQvSCtyItmtrfZRzR3iKFjuPkKwqaaaw/kSTqIKFaWvLk6Zn17cII3I1A/1Yi7j1Cu6LpWvtV6
wwuRDG72IS+Fzc7/ZzFbv2VfOOcXYUR8OCkURgn9NwWyFaXoUU+2xTcWKyr7iyeVyfMqa+phXYZ/
NqcS1RAN1BaiMDeVX6F4FH1Yr0wuIkFd0btNJEoTQ0DZd2gatipAD0rbHqYWp8QPg0LzMsEQmzx7
/jWp1sPPXb3VV8rAU00rZrXXLvSixGG4rDJnf25mmnf4bHDbAB5s4xNqGzh9SCOm1U0rAiSKr8Lh
8yKqqetCYqng47Eoc5yWIOhec59xATijTktV6szVq17AWxG3DrsAIYT1EGTBwF/GL/Gdw5zsP6aS
qP2hsA2lD/PazNEvMcCxDWwNm6mB9LqNniqZQu7InNyI45QJJiOtiH4OW+Dmy91g1IZkQFrbtVbg
6U6QA6qft4rjEHxz+ELk/22yDbhxlWuYTYcMvty53QxFLD44aw9r8x1IiCiCRHE6P4TRKKooS3Nz
4nqpEILM1fI/At2F1chQLJN1HlQFaD5r+CMW/q5ZCyTDE8bdGhHECU6dVk2HLBG8WS2OYc3muDTw
/JcqOjEhZyDW64Lys+e9qLa8DasH8IsHUP3dUSfEE3VM7Xx3+RkoTcjg5O93EzRnLhcanI0vr2Qo
Y/W5eaCUUbihfVM/6BNmQ8RkYvO53CwyKkHjETqtWba0W+f491xuvO6S6nm1PI1Cps/B5HG0HeQW
ip62eqB+zFB0G6+RYbKo/dce826LcNxO25BqKpYE96Uy8KUNOTTcwo5dInF3jEC2D0t4C8ummOZp
vTAP/jeF7RZVk0b/wQpRMxWo89qEz1t3BxX3wW2SDrfy7bfgkGe8N7PNYiV2Rwe+m9pjP/CsTLr4
uDSHAXjKdCrUe0EOlZ369lgdRx7+0/SiGHdM+MkBbWeQ8FdyRNEh71gHc3FmYJAPoDlq2o5ICvdD
qx0hSRfwszJHfCAge9cRhoUj+DFOz+VUHNcAICF0QsMuBckEUr1Dm3sgaX0A28iQermh9R+oRLRb
YZGlaV7kkj7/+7F3YNlu7S6D4i4FSkSkHS2Rxd2ZOTOTmOLxeZPd7S5din4tv3PlDQzSpgEcP2F0
EfhAs/ptanUm0aVMRNiEbFyEak3WXi/VPCm4J+iqc3uaB/K86zis0JwN5aIn5j35nRZH8zhvMYb0
UqanETZdtBzkCUMCT2j+xuyonePoe8wmifSnMKGDM4F+NsmoZjEpPFCaGosohe9MnNFEYtZTRTDs
zpctdBBIXok2n4v5ngrXJidbd+alYI38eIihOMynhYrNFkjAqTrK22qcGqww9AGTB8gKf/wVmwxf
a1FFgkwZFaoHOZdyYYrg96DrP7jfKGG+uff1/fM69MiBhjupM5y0O/R4FQbUBp6MrBGXXowFV/YF
WiZX5zHfGWmH8rTvJuJt0E1LqzUEpmDYabEYn2rJJuGdzxnxyyAO9faO02lMl7wSQb2Zh2dwQkga
j0H4lerU69lcq0vzwHqt87hA4IRYe/J2ePuDkwNtXw28s4agw05lrSQ2xLFAfL9YA4AmkaQ9OpT+
Nn5/wVf7WL3cuYb6Vr+WSlgVNqXYYzBEkuUrypOUt3ky7f65cZ7vyuF7KkxX/O8s5eS6gnY69P35
HgWz+O8WyRnoeHrKXNSJ2z+9Rmz88tqFm8eSmyBCy3sx277Um6UAXU7aI28K3Jz1VIf++9FHCXfX
ism5qAv595fQeIbHSHUeEi8DU6ziHx7OewSMUgLsEA5oyu9awDYaUNBV4SGFWsuZ9HPeMhxEN7r7
2iWgDqw1eSGkCbR0BHRrhUqR5nHhijELH8OH+k76ukvP0YIMw0T/Ybb5rrCUmfq5LfZmtIAdqgIs
3DuRkcKetpiy8U9KFE4H0PXLRyMQmPOJi3PzcIo4Jx3UkyqYGfWS7SHiEo/KwMjreg4Xn5I78wqN
jQFVgNv7uMkq0lERrBhbM0GxxPVdQ0kOFJp+7XD0tiD3HrMxp2ElFp82UuQiW29pUNgQUS5nbRlE
CMxjr03CXryouEpkAUtLbUj+1Bg9Y1591w8bi2c4mm1aPAHs1rQ3qiTt17onv4zDXYfLljBs+8Gx
XoQVh+4fdO0yrn6XDn3zT5YJQdASV9B/98IrL0ERe2gdiByjIAhuwRyqYBX7xfCUZyYDfVmY9NaB
I2ZBB5/mOGLy/9gBtCwnEmU4r5QsOydvxF/FesFwIv3GItdKfLVL9eZI6GMS8im2pziawPv+V40J
v2HDLB+soOC4kJebuGV66Q0FtYWtp6R5IycxVj4NJABz+Bmd/U5PmKVcFY5naMmuk/gg+WnOWCw4
P9qMp9vhaOlbB0aBfM28qPKY/dntCy/0xyJsD+xVqCjI/rSSNgoqHZxsfdgAehDjOTBVTcyyIASk
tIzrqceSbg0GJgQpOYILMARxWoJ4c6AOjOfYtojuZgYbd6OnPICTk06RV7tzNAKmvqY7yks2QlJT
YseGFdazdaCLlZ+I9XJqJijRGAzf2SP49nOzyn6Z/IcTCjMXTgA5Y0ox/zY5/utQ1TZIPSNjjhaT
adlnNA6k64lO5+FuJ63ZuZrBJjOtNM9QmBXOy5fdhamhIKZ/QJRDECOwLVekeq3ekOWBK8Z136Zw
esVfRcwLO3Sy6iWN1tjdM5zvVFRXBphdxbiVVSQW5f2qM7eW08Kb+l29vpN+t9EAKkuhbyK3S6vg
K6y8JOq1pUJiSmeU9GmZCOFxw9rixrAorBGeL9juFAyLrtFSC5oaw3g0nxtaIOtzMue6fCcDmibU
V+f9tXJ1QGU4HTlsmYiP3iRH1T7gCNFAGCnE7cJDjN/RR8qOBhrJ0l+ACGUtSNo9xnl2Y0pP8XUo
w2pq6VS01+tH0Kd0fYmRqlyrpv0sRnpjp2BWeG1fumnHQXKmJz9oqWobTetJCFZI4r46qmQ4AfqB
WuAnflQuJ2Ue/hVe1C6thTMVQWnWWop94/yKQrV1Y3MfVoD6z4EmnOiBedvDu2X2UHTtYvWjtihw
UkVZdJB1tYmodJEUVmKNxi/51FAvKxL63kbwyDFZ1p/T3Bl8ZfughbYUKZIRmZ682ZPE5ZHhSCpJ
pj/iwp35PnEJb0EyGRdSDotzvoF0MnO5y7zKhZ+NQICT1QcYujvMd85niTepwZKJfoTkPVUbQtmK
xQU23bBW0HaZUDyN/J3qtKdGXZ+KCEDnxsI+v+ZZD9K7oqjxRyrCPo9yNWEr6BtThZgDbOGp33HL
T6CIVvw3AP3lXMRV/ZL9d0bs+SA7ATe/VcA2wY4tF2uluHUOLVrvBAZ1P4yN2e3Zx3+RTUPcXL8h
c+7T4dulBVx5H9z1twjKhkMJVZ1MqasRKtxXaQJ9xz8LVf+l+qeWtk7T8kALYfOCPyPMFNscSrJV
NB/TTYdCO9bs0Jr4nYIx6QmxdJzYNnfQItcWuLT+GliEKt9IoMbh0qQQ5d6Z8J5Ale44K5/B7Uk3
cc89QHmfIOzQ4/sl4QzPysHN3pSeoENhyQMasYbzdjfmaKjcinqgepJ37Ty1hYovDJu52ZDBKiIg
FwFtPXMEVovU3ceO1IEDykL9b4FeBS84edC6s6LH5VYvA4gpqt6yF8sM2oMS9CsyZ3KeQDOlnSeL
OGeWBJ9d0eep4RPsC+EjZMCYgaXCfijNqmcX38H4fU+Q/3JlI2Dru08xnHoVp1YZhhEvUqjN6Gjv
nCIshfgtqSsvsvKoklMtb0gcLQ5P8PSljvmMPYmTKqdb1XCzxUUNPcA9pbgKXMwkIGujmotbfRF1
o8qDT38cr1AMrMlKX+DeF+mt4lm8X0E/zn3ldFU695hEwCJvrjuIUgeXE7Nake6aB329wilT/8Mn
aqcrLQBKjnuAE2tDDhJJtomGl4JK9iVip4SpUIfPgTANlnK67AREDWgKi/JXMQSAUgAdMK1s0khK
k67KTA7KVCaK8wOczE7n0UK7MHndwCib1FuRcG1KdUm3TQb/AysSwNo/aGpgtYiAh145ect/5W1J
wB0D/TNFr9L+aUayBQx+ScdaX2DHxzK38w1W8i/KzOl0caiaoFjylKg6Uex9OOQiP28rLHbcHcYp
6WEcs3uowWIwpM9XxbhrUlDHRZtG373kKH63D8ZAHljafKmRZIij8J2UNLy1cWZsQ3zcnDjwxwyX
DpDQoAJyfmtWQd7wpjngROTLxd6OBrMyRsLXtnFo2GSHjp8uQJabqlrd83OFYL7xx4lGISd+EUtL
MLWaFnVKn9tOf67fhfzkvys59Oo3mkZjCUmNd8t/4S3AvmRLgnqHBrmX4KSBbbcBXNwVH6BNWbw+
oNmWbLav/tkG3WkBqXTgBfT13zHYcry51O0+Om53ZAca2wYRj/zMXTp0jG/nhM5mzAD7nqIMAo4L
qiEYUM1BItne65tGTY1ibFUU47bRvD3Fok3j6Cz4bjIRvSYe4gyo+8ez9DwnqAApY1BaNh2xgwqD
N8XUWl0eNyLP+JjTZLiD9geyF1EtVtJ72OPEvKyjvj6lQIQ6MF2QxEEnOIzzEaK5kVH1lJ0q7GX8
7ai7blAltICNWSJGt0mljnaHs6WdpMl3wT1TOMuej3gN2N+oj5wN7wEhSC5Z5WSlx7lxw+gCgvCK
OkCLk678ZKJ/uYlYtDmHvHz2B9ZNM7ABV2+O8+K1Ht+ByyNd3mQ8LqgNRnAFWl1LqqLg6onljVPj
KDwrI73p/02K1sLoZCdibKfoSxgMPin/x5U/pc4DyBeywXqqmTEpJP66+CdKfEfgO5XLCKKwvsTL
T2Gazw6UocPC+hvT9Je2fxoVJHMPIAruQ8MXcVHvCcRyI1FMW+gcQdsdfFnleUJNgWxKWtEMwfkL
tHcJb3XZ+HVnOwZ3RgZvuop0ZnuEU54Ln7G+FJzYtGRZ8Pec6FUYJ4tAYwzIneGGo7BFYdJeTtZo
T3bi+VV98d2J4kBQ0Adrt4x5CgbjkDRJnWDPOg51H71lCq476jY2etYJRJfJj9f6Se3aa6ga2ZFG
yuasAmBEoBXFK+Y/L5cTkLM6nkFArr7Anzy9DBBhqjf5pyslcvLZ+PiQAcYG8zYj1XDbh+LkJEiI
wGOZjzLAAK2uY7FjlUa4jWnjOos79+QFmhQ2/NyDQjKd+EBpIgZ7fXRRcxQ5zYkoVcL36BGKH+f/
1PqMV8iYjvOPIXLByOf9jJ0Te2NlZXntzoaJkDbv6eg5zACz1ksMRRKD+s4gw/vrWaZ51/fMWtHC
ky1u5r4QVmLDQ8E/WvbpoeVUVd02PSNkiDkFI6lQeRJtXXDUr8AYB6oruWGnC4x1bcR2OdXbzE72
BpuxBJNDJgw+XwTXNZJ9KjLAxfEtALwmKR5LCKKr4EfFhHp6oDqV1erM3MsW4Oypbbku9w8Lk90h
8PRZ8vHk1IxGH5onynoBj3fteiYY6u89Rd2B0K3ekumDGAQJzFS4Zz8nc1+DupTQivqv6RaRNBtP
igEaZbr//S8a22LKWQ6BGowxb8Qf3ZwOndydGDJHtYzVRZ2p12AcwrzdEA11/yqX84zMesCdMr8L
zFsEWZF7bE96SauPolnCu2ZnBRAM1fuaXrURPU5cOLfLn36pTCxGJ5FXLKZEvODMjRSFVGkwG1Cb
mFsVy1ikPpNqLsFv+7jrd4xJBiYM5DZ09Ba9uUSMrPP+cB63wfd/uTuKOIFBSStW0zC55b9EhLiK
dlaZwCdIIxSRu+GB+gNM4nNtco8j8A0CJbzotTlfNYj53gNUM0XBGLVGKSx4C1lcFnZbwWDLtSOA
ghKhHmvQ8D4YnXekxsjZR6sKzv1mTRldn6rOVJ2NEJDoM2KCaK8eIxkmk2lXKptWUxGLQP1MuhHD
NNRPA5Vvg7LnIz0CYeJcqeg8Y2kbtDzc8WJayhhnPlMo2o1u6a0hpwD//d0gdt1GpIfxj//i1Xrr
qAPm0ts9r3o3v316F5flY2YsJTV9TePaDsoAelzVsuN4Xyp9LA1gx499LdpWWOUXG6e0u7NuEZe8
zmQpInHAQocGMQgv0eiVJdxh8vXpKRV42SlLp+c45OCh2ZDYcMJqrkZBRerkkhjt6nnFULrXvoLR
d02uf3dCru/CKMkiFChtwoeVQ8+R4qMafmRPKduaj0khPSQKXCVMb+1v4sQSVNakzNLfSkeEyIdQ
FGpnK+RM6Sxj6Kd37DsoMTmyLyt2nmEFBPEJlxdpnce/AUNOsZuy0sp81IhJjuZL2/OrqYVm/f1+
u6cRLGw4WX/zHCYfZG+X0d+Svtcbv97000CzsijQF4oWGxPy/uPYmSSdFycTS66TgbLl099xpBfU
ylJyYQ/SBg/2w5oAZfSfqIwEsaHU1E5ieRXn6/QetU5WPDhnveCL+TBvk1PliUd+BPUA/mxH3LjS
SxyfW25z11My+q3746SGYUHVVlPkakRTgVe19SrsZvjagottYPkk165DTCnh1I1hbhTQPCQXgKsV
u6oEtSssepbmMcFzbWEQ5fEJ3N+l5EDRJn+Kwe7c72ECPMbIM7uvea/Pn6rnYrOTTswcgUVR8LMx
/EJCzavpapsrr0RaZbNyFiPpkb6RDQABv/Qk9gpDCU2jBxthccZtnzb66GeoXtdakZc/UsOb56ww
o80WivnTplqK7Qd8qn94OAgCOQ2MjnDsVkKsiMJOEs9QX8JwL4WtxlB0e4aqcHhk1HEubxPKdn4f
KchTEg03RVXsX4CRvwKlyyxp53du0WWWC6uJXj+CRzxGo8LBUCLAoFAaJzlDJeRE57D6IVBjv9Ju
wzpYYjOcC86NumILVuNzr5hcFLBI/uNcl/W4TN1/bgqKnSo72ZJo+7NhH9scI3Mi6BJURJ02eVh9
2ih7Fh2QsKcSkix+L9rqrdw6l5I722KvmYCofqCg0cS2/Wo51LUK/cqxsnl2G5Yd4Y7UPncKqgRD
H3JCQDuFXy/US5nJhXszUoY2UeFVsKx7gJfAPwNsxwiVuzjfaR1DUmbJEenK03YjRQQ4couSH13C
o9danFIh9kM8KPBaqWM/3BtzXoWbObAy7gBtEA841k+jK3ADyUbSDAJ6WVWQFzB2/uly6EW2xlyI
yuV7GqfmJ671/eRcgY39y99hYvRzQd5UworiPWobvqiI5+FRV8YN4kNIPsQ6MAqZY6I1G5HgCPfY
Ldu5con9kTwzpRK1Uy1mQ02K5pbawClTQhzhJ6gEsBWh2I/RpxuJszHDi2Ogd5LASB17Ab8b2+qn
1rsYNxqVSB83sNvFrl6SwbGPfj290h6cTTc87PkQzvcHcdwDJf8KaLLjkZEp59tOSODnx2mhHhEP
km1hil69rpoxoQFVh1bD9Nw3BoSzmSxFw6/rJrM2Hyg2S0m7hzgZpwQuZSbBJELCkVmLPgpXoPU2
G3RZZhnQ5qrQLwWgEI/+BI/GO4QeFv5NvD37L/pCYaoYs/bXPLUsmdfyV/cfxesKFoN9C/EeW6wC
c0Z06dwpKFg4fK/OGC1RXA54qfngePwNhHvQmzIxaFpPfEN22fe02AeZ73ghB/+0HNb/Nrvz8xVL
pDtdM+QUhPqT4sZBG90/rixoH5bKzOXyBPnf4vSu16n/N5RgeRfkVEXXgiDa8uj6xygLCa4VR+wv
vPafidvJ+T8N2rE3hQAwjFCQGx+CaI2RWZny355Od5Ozz+59qSHohT3wkuu7QwpYEdIEaTbPnxbo
DJwVbjG6peHKfT7mZmOjGT0EgbROrO1rv+fPYla3XwbAONn8p9B2Svok3E8x+QnJ7Idk8X7RH4DF
IBMEaMTJ0gWFXss/k+pKQxrt84IPYOixEovPu3h/EjbGD0EwJ62xXPEcIP5kBRnP3k0UOkyvPNEj
ZULqJ2NjId3vCIhJbC3u0CaDey7IsERQdE/0rC5LzJiKIz4YA2d8WnIWmKJrsysTACrTn60Xotpf
KtKaQTQ9hlE/Iqh3cgs13fY+/Hrtmta5wILV8AUD6hqiYBx5pcYAm/hbLW97NkxeKf8KGqhwIPes
K2sLhiQs8/z4cx0AWi09R870x46WmhRH5s19fLktM9oh3H/XAY6AYPihY3xFyR0QrN4DEL5OJPnw
T8TljnzkwODjyITWs57rvIgYz8JZuzuWq8BtEOkFuCCDF2dsoIWFB3dt4PrfVNbAqHpSrmXvRExO
8ws+MYrlCMhWCi5SgJyOHN3t8QB05VXKOWfL94XvvK8D/JV9SFAmM6T7lLF4mXhi0LHCxQQpWyki
g7g7HHHXfRdgmrvGsAy/+mv+p6REHQhL2Xgax8Bl3Jl4r604p5+Fn9+cxEdjJ4Ug4XNf9Y3xrQfX
3cGcKfJBmicd2u34kkIXtnTcYkxRTk6exGByQad5AFV/G/3kqjwQZOcsGLK9veNYac6j2kTrmkwk
uouccrbR/lfg3YFVp2DUq1RiQuEFF72KR6OpJRFZTFBpVczyv4FLXrl8rp3lAIQEdVZZCi4SU93I
S1lGyFbZBqknfg8DMTIsmV6MeqTd9yqVmGyU0rZCQ6qy2kU7ALPgbqM5f/w3TttV5jMoTNwDyNuD
cCMp0OWCdLhVX66YEhK51hJBiCGV8+GuAatpl/pJrgKEgAUNruXgn6XtV6cPdheyLq9HBhE1JxGc
TkD0W3HcUm2qvA/dU0Ud9f1JdXZE602nKYvU8WGU5IzfAtzWLLygxVtWQ6iAgG29z3iXwi1ThcjD
S3AGq03LYSUUlZ828N71mxU1DgCLPdjVHGmX+rVdNrvyL0t9rWNif7E21WakAnpyfih3FLVFzqEP
8c/cb9zjHxxd8LEg2ExuXxTX/F1lHvhpCvADkxeUQFhnw+HdVmT+S7xyXuNCxLwhXhAsQFOd8QE2
RY7GvBOyeZKm7ljo0mp6Jqyv8rlQJ3KAohPXXGTasUMp6I9XSMqCDe/ZyvNl4o2QlXJbj2xa9M4D
V35+l3qSv74JIPEkEaK66ojSI5hYEB0WD1EfBQM4ptXStAGBVLe2ez5TqRXKPnY9qAunJG4HmjKN
mRXNW/q1kZiV4nEKqVpBz747u3EUBj4NSt3FUbwJmQ9LSDuIT/y6v2BUpSNXP2am83vb3kKdo2Z5
12nTFmnQ4kklDzCdQnrjyCNNp4RNmREMwhX7lABuY/w2TAwoQdJFzn0X7d0irqWiDZ7Yc57CQxuK
yyt/613ZMEcRuQxuLRlvLfzDUqTe6ywjCqcq1Jq3LjFlVI9iyUWnVY79P0wG9U/jk6NqOGcpdNP6
TOxmSVggQHNGH2Y61+1c6DK9w+9K3o0ihHDS2QHuaiPyZx+U0BM1sTz9SfR5sdZDMsVhdIQxcgrx
MMJ7T+oLLR8CuG6N7LPhB9E8Sp4NVsjvnj76se22L/Hkd1OXeodDwyNIJGb65erZPWbkTTvChHc+
VDsGv3AmsOtPRbiJLQ2qUzGD8QxoXVr3BAAvytP3Vaa6fNuRd/31TYoEOaT6f/WemodU1zCquhYV
wjwAtlwAevtXFtjga1xKP+ooTU7pRyuzntgOPI/Pu1d1hwYU1Ig5v3GWoY+bBYA/j0yEKev46wT3
X21r/txuv379+CmM/xVzmYnj6voYCqIxnx3hxkFRpMZZQR6+kmoeSM+8SfLnfEQQDzGgrPIVJiN5
hPC/fcUf4GIGNZKOqqucc7gG+dpvb0YtqLlNuqD+A5NUg/WlB2FMF1K9Cd9iXK8eKlT5fKBt6dtD
LtyXXFSk0YUUXKPFZoVpUwJ5vTCQKXwoxYMLyBXeYZ2asT0Oyby+G+0REHy/YSs8m5SqAYeyEidX
mNP6bcEORj9a5W2ifD9pKxEHaGeh4mSBnbx0Wd1tALJRhDSdVC/31dxFgBrXKJ2Xy4tnJzIgbDH4
acFUrsDDMPvjxzAYQo2uQA7SGExtldShMRTdxvvwWtP8eW1cd9vvM/FeoQm3U5wQSVDlkPPkrGBM
jAPH3Hz6UpwERAO012R2pRbsSBWFPL9+fR6wK6wSqDMYyaL2r9CNj7+U8/RETJJS4PEYInRIOa5D
XEhOfxI/5l+1Kbfx6SRikmO9YRPQ39NnrJ+DjPav+XihNVP5a+lZ20W6Xe7Be+mfDKbPho8E70A3
2aLCfaqq/5vTk26raJ5LO+IrV3e7aGvdETYhm0z/EKDQyQCeuiJqKbunDJIYfrLRvTV1xm+B96ne
F471ZOth/xSz4nA7bt+vvOCKoWU0Bj8plHDMzBbMyNl1LPQif9gTmLBKFKIoszWL5vjm8sDorMCR
cynWxPNMlrXxJzhVVk3rJiuXJNn2T9eKyaiZR5qvMYqFzOQ6BK36kdzxZWRLRXFVTcXeAVfR5qBp
GC/umIbzvdsWZPOWSh376cyiVy4rcZ8AuG5R+7M31R9pc8qH4Cd+1mQLC3lcWbwfapxIKO/FXDB+
EfqzARetI2hoXihDzvgbKAWoziSL0PeOGs7hqcANj6zKrx1/VtVkLWfGaHczGMlRKPBJXEWJSeDD
+ABqBMpCF+wau8E9YfbA9PKIBUY5EeAUsV37eTCoxck56rskA1TShBNzI3GEcwNtr9A00FS8Wici
lFTfOrLsh7YoT/wwKZ6ZXQNFvr0nyJYmEem3DzsRxbogSxrEI+nC7qClVFWTGGLEWf3Km+Hqv0P0
68phcmdDTZ3LwyWcLT8bM6gTDPLEhAqczMNs45BKk6WiEvth6nf4Jy5ruja77NsKxTzpb0HUyDiB
SgHyjiCFrc0o2zq/YUtu7xKfL/UM1hwpMYzKw3S2gfk09lyEBCzkJEVSkw+/ZaxevGH4EAx5eSzd
gkenhi7039F6ocv2HUriq2qLPQkXztOZ33Jobf+NCJcPOVYuqm14WrOk4m0L5tz0ax2SQmsVWSj9
jmeNqZGZWRnFhXAQGMV/IezYGNyyu8bXt8g/9GlA7SBmri4u+6NcSyA1luDXL4Znwg0rbz0soal6
LLozPOxxxX8OK7QIVLQOdDz3hHFOt+l0NhBSJ1o3QetcPUzV2voW3o2ceRlWTPD7UwlYuRsrEPBf
KhJ2BwcbQSvWJrQSTlvUC1vsDK1T1sm5EdmM9J7TXHi/YggfXDsmobHWLawCFnQ/WFxp5HXNaG4a
uNfcfMUsWQpIGZMx7ggD/lJQPkCaemZgg+wrJNZeJrA+x/7A04zJ0YG8+inlAxyEsAKMsr7wvzoK
cbslSsC+rZKOuTvZ9i6iKNCJXNaHJ4FQjkBfjdmO9Do+awT7kPFml4p2obVOhoPnp9vFVcbXavpu
5UyB7Xqy8kongSYFXGF3FoQ8g24kHwHakpAB6kTkHP3mK/fTCOZmYbZH1BwNZ/L/1uEgUzomvpjv
RFQ0xt98hbH4kDbzIra/mcxuNoeH8v0cxrD6YXAbigWgYMRv4TcCdrXTWuwVKek4IBglT6NpX/UM
GTNudOdMYAJ2wDa2O3DGMFt/CGbVVBonu9KR5qpwev3HRoZyMPDHOv9KnJDjuH4mhGppjhesumbZ
lVLZOJGC4D/rHzxyQq0dca2hQOO9Uo9THZChY0Pro1bwmaYPc0+sqOeqWzUzDqoL+/Rgyy7H4M3p
79MMg/N8OqksfCxYSTZcaOZijs0f9M666MHvc/zRHTP1hr+F3ntYHH/TGxuwVeP4Pp1gzGFpvHwJ
QkgouXt2mtmLaW+gC6w31ZvQSsHqTc+RKnGCp04iZ3gD3BkiADPUcVaELSVQ3iYN1J0uaLnjQ2gu
KoPkPVt64tS9qc48XdQksDIWsj0rSqw0lfUM/Q4bL/8JxUbYWuhbk+Iliuti7vj8L4T0rmXNHdLg
Eaet3l39EOE8v9mMy8f1D8tId3zT5B2hQA8vd2mWmSWnME3cqr0HOw8gdaS4I9tWEgSDo/mH8CIn
346sgdwdgC5tq7Sibe964XnVLsOJ4wu/hrEI2qSp/6XyzD70fQ1jyUd0FvvSw0EwpcqZEIf0HR01
ToLfp5lkiqx/iMXV/dL3r76PtZjAGL6k9U1gJxEMptJRuxyz2DbEHlESFxn/EmAVHCewWRzEVIt7
Q/yk60ae+D3V4rz1BcGnZl0+B+IB/5CG/j1WLU8o8r1MCJwpA0ZD7tatKShKOQqNYQUrFC/Aw8Ts
xFnihzQp9LHb5moVeq4VA0fBAgnNcuJTEh2nQcNfEjfsZCwycY13eEN29boTGgTBgF97Ka8Y2jI4
a+zS2U2YCpeMCpZ7LvsVEqZD1rHEjU5kShd17lljLCeCDJ57JixbLjZYB4rY9+SpUywIFFCUA8UM
d7wXegw+8ZP/FzMGlxMlCv8sLabhOMG6Y9V/aekZUzHlAMRCOH7/qWF5H8uD2aPKfXPmSX/6nh5U
K8/FemDy8jJZ6EPCTfovILWplAjf+yAZE+i/HaFxge/rpiA/e1Q/LNR2ioervOVvo3BEwSwXami5
5cqjUUfaiHLSDhPNwgMyp9w8UCkY65yRVsiMUxqqLEk0/36awYXprrm/sNKshZ9JZtNXRpCS2gD/
WSew/9/IaIYoKP0ewUbp1z5sCDGJHZNZvRb5+2u6fp/079oNW2eAK2jivG7ASb7GffBgi2ZfUsxN
e6FkIQXZsYqBvKIuZ5rpKEhWR09bHoKjWlJOFycySKTr7B8Vcs+3PEJlolyMDlZH0kYHt1ZOjUoH
2bJ0d9od8jA3J7SiIBRQPZjEWWTWyy84KeLlQYfUiwUtYI8DpOeqIBRRdezrvt46EIyg1WnBkwbP
yHv86vyTAaWB80AgBcqg8crm9x+jvqZ4GGry9SZocAPMVXpKerpzInyWd1QlKcF5wQpNSpWHAiSO
8Q9CCBoEBrpR5c4Tok0kbNnrZpjNmz7FGrLkLczfdH/+GKjV5byVuvVdAYYRVZl6/wrb1A5qhVUP
RHBDhnfFoUqeV7Ru+MF3KT5mKK4qoSsb21Z+XgnPxah1lhN22G4EL/Ka6BM4apDGlkPAT+Q2WV7v
3CEpbDljC7hfjtFBR4hFaOXVW1/0CrGqUdO1RDfO2hXvsdxNOrQ96wXCrPrGco3U/xnhgdHgBneI
q4rePZkrlQQnt3DutK3g9G9gBya+G/sdwwfkS0pPU9arw5VEmVSqhi3Owmneja3FT1Jm1J67Abul
B/EOOSlXG5JaMNlzufJxfCK9RBzlFu/2bEGK8qUFpJT2zs2l60zg5d5S5hkNvIUcly4iyetcP3fN
mOavmRTA6TkOYipM8ABJ1EV8WCH4TZPNTzU4pj8wGmVEk8G0MGzeHFswZ/a6XCgRsw46SgDbsYhd
22mxDF8AcRkxZAu7HoPUmKI7JYWhNs6lXgFj75cUiXNSDiQ5gnPNd1RsK2Wm4mIGFaiY8XUKb2z2
I2MyZnGa6jMl6EZEnrJ2V2WEL9x/rwzJ6Pvaeu7o81nagsYuyDlYi8Soxsh54rfBBwOXkzChIz49
5NPzNTlk2Dxbc8L3VBwQ1y6kd07yiYnPANTqx5qhokkvWoIQHmW1sRuUG6wkfu2M0WgZwYzRN4DP
t+lLz61OEK2OdKvl6Xis8sXBUhAhVHYoGcMw5Vu3Wbn7Ljosx220fWU97Kj6V6mXKlKDweiUNCag
2afe2AYUuUV4WE1M1fa+BJqlKbK37XV90XTS96ct7VcI7K3GMwVBwykEXSpwFI1hiAgU98zYDJy9
1Dq5iRMPG3J11jUqjqvzpcliT2hKy8voeuyEie2NkCD1dAyfpmWWBlOaWXG8ePq24CjjjOS3JRIq
z0Kd6PyoUrK5xNZLTIksQwMAs/Qsq2g7iBQg5muaPCDHmumHlRIX3UUPg3zwHaKLa/PZODKYUoyb
80Mi+4Z6YKoJMQnXLsew97Dv2rw9y7wD6591YhG5M08tMMP6RDBNYDjVAzn9+pV0gVdxZCFRQIpM
ZnrrDBNDugvPcFC6MVimC3kyN7GRZhU1YSBdItlECfvho3/lf7fQpMbDYSeDk+tvNssqYlEPeX2n
BjU8dIjFOmxpAXwGWC/yzfIr/L/C2Kcr7/pmPbcFex3N+PvWpK/BsUjtozq1cNVstRlm3X2cJsJg
JdT5PypYk62ZMIGbuAfrXu6jS/t0slIMHQdHiWQIbYCVROy7HWlR8JruW0+g1tVxsxzrj5ACUs6L
sd3A1Y6d4yGsxRTPftU2UJOjbW/k0IkdGFuNhQT47DBsf4DFfCHt863PIyaSpojuZcPvCSgsn6F6
lOdCnP7HRMVvbibKNBjsedB6nk0T8aht79RRMV6rHS8LiH4/y6Jyaa2ywqZlidF73PtWbsn2RYyy
THyAzi/5CFmjNiV7HYABf9rcOzf58rSozHEoZv6cMcAKk5uIJP4DkggbFWZrkbHmDI83J/rIuVyA
Vnu9pQ6Is4ny1vf8w2C1T9AykhprUtTfjY8RVpt2eH72Q0f89T/boj/X4ZPw5eN63LCcRI7Ai3+4
BhYLEpm9UqW3c/R6AJ+VpyChFR/ISu+NpYvu+x1b8i2PZmAP4pWAAyr27UbY/NK1kMhlJckLVG09
CH1ZEslOPVpX1UAzqGN3DJ7nb0BFDaNUCfW1qp6G9soloTnNr05OzvGjDauNVggoCq1g+8wvzZu2
NSb0jLiTW+3JiH2FoTPAu32IsqKGG/JASokOVKhct9Aue9rFvGcidD4e/ruXYBDbft+J7H4Sklxz
krDtqwiv1KyBL493sZBxmE6hntwVDk3dx+fA0lsy8TSFfeeSDREJNYDeac34XVw6xyMyYh/lhLJD
NvVON8UlwjcIM0d93NJNBfSMEGJex6lj3rv3kNDbi3U3TYvLsHoBUhHuo/DHAI6KY3mGjGk/7dTA
K/wDde/zvrow5RuoLm57qW5m+fIeau0dcg3ycJiB52MtEqmZFej2oapIMjxt1+SjG428OC4L6tE2
K4FWZVoVS/imzIAAgWt/Eqf/QtgFbDsHfDCptOaNWvE3q00vkb8ONTYQyARjwPB693wB8Z+0TPxc
ULgkDM0UTJyum/0LgwSvuRVQYfgEm2qZQJQ/rqsAM3OC2LF2C/v+q8YiMr0ZrKJ/0d9sDGPZY+E1
pbbuK73muL0Mj3v8x3RfvsjFHr5AAwOURJ2u/wFPXLKpRc1RPEgolgYGJlyhl7vtXEXhwty7Zys8
aibUTSetrtszp3eTmUEZ26z7jKQeKJy7oq+6PSydZKMqynef/ixRyiKLvkYC+GTEDXc7tXEmjOsi
0+VJ0K/vS9AxMi3kIqAOevwtDduABjVw4PY9R3wjWxVb+nneO/N/Yvhx3+duqIDAf/IEAjY46M0t
mxlIXelTzm+GzemVPWPKpjugBjQrhvpNaTfoSov9+AG9vcZRX9Fpy3KGNwhy5ZR09ts02JKBrblV
PKfO+2b/S7zIAChr2kF9Sgd7KcrIG9NXmpWa4eSFnmu7mcYbcUH5NEFSPSF6pHIBbkobx5bW/zOM
pOB8NazdATkSBQqc6cHz35sXk3s4SHyuUVv0EteuQusiTzXARaPcQw/9Qoj9DOWv6lQrR0G4/z+N
LhKxAowjkR4uxyONJR0vU646hfglZAOs0EdAxodrgtOh8VyuHKkKn7O8BiksmNYl4xb1TTcPgCNT
M3mi0UOjbfV5D9bPvj22UDw6/eDSxqkFpvf287IS8xyKrRzHPBIFzjU4oOP39a8+biTj+bxn0Q/z
uMA5DcmZMN9v5mibU6lcy82UXBhqbrMDkekpqM1ov+BCH68hl+bR3UGnfCI3Lek2JWZixQ7d/nWg
wARDJlrbHTSDeKu3P36posyZFyAzLRH+UKHGmPvWCRZnpKRq8KQQUOOsARd9I+mQPcGMn4GTeqvY
SluJpp5IyEUkGS76mHjGLuKzzQzSODspjdCsR1fuNk8PryM2+6hvn0vsbP4j82IVaNs2dVCgxazw
+ffp5fz8rkC2gcvknI30nc/big4Q/LjUu0T1GktVV+e6EgTIpOF3rs1dLxhZQ0YT4leni24sXWz5
B2pYq+7gopWleVIrSb7QnMeihKTJHObEdqVU0rGwr8fSmx/0qypGjYu9DqlOsr6481GKpWq+Pjz4
UtHP94WT3p/+nloHpeSrRRyCifM3aVo0AwHcKe5pqDL6XDUbOBuafl+B6nHKypE1lf0J37vx4+Tc
YwTLZPdYWplB3vPu0wDflNh39sGuKEKfwMK8lyuThFyH/cbomGAprFtBDgKSFeVDx0PGopO97v5A
KSIE1m30Wldo0vL3DK2ZGnAggUw6GJybml+kj+w12bCAzz4QXYl1YdqlKJjHtszKiizStcimf6+d
IwirACPe9ruyK3XKuKokBM35rSM9MqFtBh8Et4iggwzYZtjeUDidAMEE7HaApF2yv7sCC50yIRtd
9HYRtUYs5matNyaKagSGibE6j7UlWJ5ckOQ8LYz+oqyivZLUgRPch2A7HVVNzLV6tnYvYXFXnX93
i9jGzIYfrAKqF4jD2Iu0LRG93QPEVYITGN4nOkyOc3qrpo9klXtsE/CAjJt52gP3kjKqsz0qxeVG
afykb4AtsuQXes2SnOTeiVgtWwV6QenKd6ikk5lctduQrcx6txmJX9Nu98kEtuWNh8iZGCqVCBDl
cOf+8Inm87GKPtMpahtAlDFGxz0aYeiAliw0uDOG5EefOQR2++bD20pnRbraLp1wJ/1zyw2uRVCG
TeraODr78sH7knbes2xuGP6PQJhSNOWosnkS7ZV0Fvv7dWHLgkhMLONDU42tDsH4CkYidpuew3Fe
f26xQhr1Rfupzp4Jb4geiTmtRYf5vvhnabP+9UXIJwZizYg/2rUu+VEJqqC/G+3lmqngGtMtS79+
eLMqGRLKOdDxfNApnwSEYCtN5Zuf21ywmJqAFaQJ+1c41E0BvBdzm9yING18H1JRD17RGot0gt37
togeYz0FHhusu9Q74SpvFmHGLLKju8r/tthHQCyugefTjfBPorNmoTihKZ0AX4ow4qisqWWBJlW6
oCTwBhhI2WZdoFjAp6ou9mr7Kh1KmzsQSGmlNpnwCQxyXm6TOaJX4cI7jp3eqatPZXuh6Qw81p5K
hhlKIW4ny6keH9eAe3NHh5q4jWSkS3v57grtm6bdGGrHRY+9LJjGV9ylARPPHVczydrp5rcqnj5r
Y8WMvTRCiefG6/VHlCRVF0u36kHecoJBdXSA8jg4fSGLKOJaoacpj+7Sfo1eBuIesZGKoMTbwzfi
tTYzY0P2kLWEPl7BfKAUzQ7HTBlWcEWnbqq/ni0g/nPmJNkU8ORtLl2m2isoUQOKeViwrf5TV6LZ
obSFoHpj6GvCLHNIM6hXCFjLbRApdaJczIrFWqvQaaqR8AvchAed+lBP6TYHylH7PnJXzp4IBeMe
XKxj1EuCrsl5xybm7SkFDV1rXCTGnVWZyfbxltd96ExsI7hK77oljMBOkVtUZFfs1K7d7qqoAguj
s8FqJEN97/AvQVE52H3o9dxeknpmL1BathmaHS/ebe4e8eV2NkP438b3iY9mrCusXYZAXvk3GlLz
M6bgpfcEfQhHRfvna6FeVdS/RHst2QxtivXKhSrYf+qmjo7bAf1wbw6VqtqXiq51hhTsXWRa8XbH
WQ0Mqz1VFHZCy5Uvb2rQmmmkDCRo1myBGlkGLQnUoJce0NEIBgD2ekObE5v5lyjy6xtDdFuR7sAZ
gFgiT/7staS1t5iA9nkxDY3DMrSoZAUSzQUEPuBK0iYhw0yUkiafVst1RDl72pGmgQYaRxehP7r2
5GrL4Nu6iaznYlo/POyVKBYhkhWs9Q9kMTCJi6ZILjSkwlsLA0mF8ObQVHyOKazRdFD5ddGOp1nl
N/cG8LUShUaYwtgmf7JF5r8XzvLFiq+HPPUmtV6mXcv67ddxyP07/DjVu8mzkCv8TU+vePyNxDFe
+5tn1zq7WAQhd4FCxLmXX2zGJPauggbGbmUDDdNoa/J5SzVh8umxXBGHy8SvFB7GwWGM30aBWtWz
btA7S+8mjFxZPGfL2oPqVBnrM7rgRl7CNsrtxE3PHtqNEQAk84wIPCvxD8f7r6BcFyU8dfI3Uu9S
V84BIlbG27QrT52q1lt7HHFTkdArwAsOx0C2H48gORs04p5IBn/akjhuEas18jDHDwsIrmaUCDdP
vY8RVStlyeyPo8MTLk2Pm1x6ADaU2MA7z2OIEXKxxdGtUsiqpRp64TxmWwduXCqDbkTSOPkIamqA
EiPGGf9vjaU8acZS3XZQYGlZNIWtgOFZ8RnBvZfID0yLdmCFS/O8d8dP0P+YcY855hcKIrmUyAlh
WbdGtR2ake16lQgbHdun+MXU/LCE9YQbHE1l2Bnny9Y1yuXYuN84A4L/7tKcUYFRuY5mRZUqctgu
9Y+0Bai5Cf2iHHvQhrAH4oC4OdiUxZLG8jQ2VRhQ2yPPfAzp9uoy2N71HM4e2ruYX/dNMFPthsFQ
NYjRBaQZWwSDDWc5FogeuosQgdNMyuHAZz0AbIgZWgU8HnEvFqybZmlcFRtlMwZKQqikwdcX1i85
7f8ABxswxeqQvXq6/XUupLgWaaLl59aXjkxGmyUfuMqz3eNjcFgN4nnWsHrbquwAPjfBlOZE3Bbk
HoTqS18xV8Z1IyYfFFUCqEfZNf/XYAPg1QUxZ9rrI9PWKOrRPYiy+EE6XAhYnGxOnAmdiUOf8QBz
zcMshfsOINAwohdu77klcYTBbRtUlV6Fl60C8IqUEFG1i6RJOqvcayEmKm11F6hK2o06wSCaRlUc
HGwFZNJ7CtpDdy1Cl2morVgXvxbfbGQ2z07Rglm4kJ8VXeJwnm+5qREy+QdpmBDY18DFMJyhSpTE
aQHXxwE3x1Ehqbim1uwmjbfFJEf7el6usz9Jhq1x7eJtMtgsCVD5Npm3JNw5sRiwgMspPgT4Gesr
wNULkDmKivY5TxhtU7vLPn/CCaUpTPvPFIjjeEQYZ0b8yGzrFBcMOi2ZPMqUSTJKfk/rld/hA5PY
zU1N0kKgVtYIwOow9i6vydijgyp5YD2LFSE0gig4ZAHFbN8Ocrax7zfphXz+pniQ48QarpACn0U0
8Bk/JA+VqzrLDSeqf/EJRb10K6y1JN7VXKV113ZRdyTFivDivHey31KO+U8R6ZbFlbulMLg6t6OL
jR/gcQp8L3+qdA2UXzv5CawWbt1/HTq7XrLlnN5wtChKZSzHsb/ak78xosCDymkGk52/JuKvkaNi
+1zVXkJB4OG6ML+zJlex2lZijklWM/P9xzUNILPenC8Q/l8IVFMHlwBznDFPg4cHzCBLxkNbH0Ol
NhNEVfnHPG7pdJvjOxCTdDdoUh++d90YKkCCXM5TYzr8ogilpNnClcIkCXArs0KSkzetOu/gcPyo
wVpXlCw17cfpu398VYgr46y25thnXkmtXF00o7vPFBbpDmRc1Nxjhwc5j6fdXulhxjHzLV+GtQvf
nYwtBFMUj2WFplHe4QBtpiGtrQtrMueddRiEJiglY7guru4Q8TjQ1/8z1vvulcaDB/f3Vf8QLNGf
LA34E7H4Siu83G5AMdxTpfYzqebH9s9dPYWZqdi+Dv+zKPga7rTaLanr4eB/HdQhfNyW8ecarGVv
Sb2ew+6plKlm4eE/VECs1vV2imQ/585rn7kPYnNX0NhcIGAohxM7kDHX8F0Fh9G29LPmkeEZY5h0
z3kNhVYa8aky+VXwTi4/55GQzyCM7xXr6FQ+Ag83f3YS7HeWlI0+qqwECtG4h28fw0S33QTkAfNK
+UhPXCEd1JELnvztNbt5AlyBlMryiQGZGTc6LuVnJKMwwhyHc8FAe9vPLtlICz9X0CwUPHLYCJmf
yxEOQTRfpknGx65g5KnF9XmLmQa32q79Kx9OTH3g78bn7dk0SJTt5tk8PjkUHU+oU7L5mWjgmvLF
0gskaonyrmZjis7PqOBJhrW6ZEGFdwf20SGpaOAk6xiQfSncCUieUr4rUifkPaE333/gg7UrSts4
iKETgNk3vLt8OASdgODlrlmQdhsu+b/top+/IwXrsncKAY0y7iq1NW32QH6Z8oEyG1u3HHZN3L9y
XFyvBEUfsWiJe4l1v37P2caT2ASgpf4qSPx0AYBVXR++sKqyk8huUvaWV63G73E2e+938Lki4N5s
CSovnSk6Dxx0jD6u631gl8nHNwOmzoV+06naPaSt4+B8Y2uvIhd/kazdaQn7qcoEhjt867TO4vft
H2wEugxKjEGEGn4rbYptryKqg2GYOWO0oyZeIaIDPrSSU3vDE2MSytEBq31eDvAgDKwNj7F/r/h5
kIjUYvNacQUM0Jv74y4k+2b8/xNqCbWI5bASnSDhXGNZMMdsqMhNbORB4T48on46JF8V8ONLXqqC
vQpxfTnQrw2sPOpWa/0GFzpKP9XUNkQ5ArZJ9rRF32TRchXMFjhtr84LEEVEutXZlrwFiiVfjS8U
R6UocdbksezsH6Xvg176opAe4AC3xCKKCBO4Hnai6QOB6eOGzdP9A5wHmWbxvYgUaa21D9l4c+6q
K76NU75/XSION26V9FPapjPaR+znPlESHoB1FMgRH3zmqVJBGjYG2R2yQbfMi9k7HgsEMGTZEHeR
7YX16pdyV8hG+mecvQeYg67tjYvzE+YWKB9dpM2t7ggg/7m6mcLx7y/0S8Zn+ScpZmbVH5359h4X
1AkRzmTP9Ua2ARkVCwNPCpFlsD2gQ7tmdZ5PZ07SH1OnQu63ANIIbQxDExpTi4WQUCEz9Kqg/xlY
Xt9GQS06ztfLTun1gGxDWwyZuJpNWYZVud+XuCEin8efh1AFSRfyyNiu9RoE0LpCApEMjG1SWCEC
M4WXXtOasmanyrCTcwfwFCxFIrpPlA7ipiuILSaxuGjdfRYoJ/dCsXcKXWCcrtw5g44FIq1U7GO7
aKPEj62Iq9j5rA7Pn9or3RpL1iAjyzPemZNbwCaqWXyKp7tHGP0soEYXncdNi2cqNufMkn7GZLhJ
KCpX+e/Q/Tu5d2Zfuu09vCuYHJR3VswYnF8i38NjLQGxpLwxm+pQZuMlIaKLijp0RETy2MmjoU2W
8r2Xi+4gX+mbYLnwPEBeJ2vqPN0KIYDsOOFStkcjrDYeabiagYyrO6mkdf2OT0d3qHJDABnCh98h
bGaAMbFFlo4X8ve5LeYc3VLTLMBLGc0Q0SHJQ6V0KI0jbDP6WFm63G8uc/+GpovMziQ3sEC2c67x
+D/PjzBo4e4C1tXwna2K2Xg/E7mw4gyfkaJ3gGWtLDnZvnKOCfjsKnPt+aaEMzIKE9tp6gn8RmiG
ouPtBzmdqw/R1fXnDkXO7mMfAK8QvetvoshZ2JEfbeArf9/gfzjGBTlQkE0ZpqjCK/bcryxJadvT
Fo4NBy1++ykuJzYTrPDnaxRvql4K4UPuJorcFKdX/za8sGK2BcfaIuDSqtmN+tuUM/E7Ce0O97Vq
ZNY03wCkLismGlMv3B1Bt1sc4xL3yi4GDcfzIVJN3MYJ1Q2pZ8dW/umpCzZPTYCuSlKKGd5oLFm3
6S6UWzhBXvoYx4jAvr4Y3s94gKi5qKZhmkfZhnCtViXC3K0ekWJpaLCsOSxu3tXuMQL9Kb3fid7p
1oW6EipoASjKF/O+fScZvuNCfHWzpJKlKg53jXeMNxT2M9zsxZf8aendhKcFhWe6XaDA4wChCb11
BRw387elcrc7dWNCX2Njdit16qPT6JhUIB+iTskcj94bcjHQcsdZueqnBWdXH2VztK0j+5nDOvo4
mkGcfDe02h37NNkTampt6MkTweHFhbZWbLHwrVqGYF8iHCnFmrfVNTuvIEhS+mcETt96eZtwWJ21
bhT43XLuGjp+N/T3YAk9blp+howjdlhMMaY84PF1oEHy0+uQaGtakL31uARgG0AdjRRQ/SKgyvJE
ceEZ0fakPaDN8p6NmNYd1qO36vLpgF31+CLSaLYGpO86LGwzaOYcbLORdmBK7W3YiPIiKNUChusQ
KAtH2Syaa9tGLA+UkLBwYUZrVgbYa+Pjqot2A7rz3GGdD+M1LMFzLJ8PyrGBeV+HQ3qJP74POvRf
dbWPC9TViYGcst0t99dBSl1YakIMXJjhjQzWnP+OS3HOJ87BgBFSXEQktibazwMU7Pp2Aa5bQ4O6
N4ZyPG0eRww9eiXuu/tFU64p46mUeoL7YjHtxtYUe8uipDHyurXbJgaLg1VJy4SOvuUstMIcEY5U
frSFRuHjWIc2UIFI+ogSpNvcqZjz34j8DkgOo7Nxp8zc7eUmNoRfxabiOjSq+PbRyQDSz6Lm/lR1
VveewMXzNJhSw/y7f7hx1+qP+AOykPcZMey5RIAP/H0JikCImXCYaFA4oF1TiSoEluXcpws7TiSg
uPPY0DV+sxVGfsm9UfuKKFXSVy4t5iO8ToeAVHhArmUjJoORzst+CKgL/M94AKlrHez4MATndVb1
gaXSyGrtDrWaHnuvoJE3v4JiuzIwTIFhxu51ShYhpsLMRvefOGTBx4KDDIlZFZjy79psh+5BWZH4
S7L5cahHy7rYBCNt4WvK4CiWmSy1GPXkOwd1akXL8bGyzqyLx+KQbkUlP8gA05K9Ts34K7LifMUo
q5oJgHRc7v412vcCCAnwvObDe1nWtVP4mXq+PBrv4Zj6D8DdKf6fVCJbKeJRWQXqT0QDKVoCWmLS
LmvgT7R6M3teTMYZP1y+ga4LjKxYodxg5B8THFr0h0VSW3E6uMiYtNyHdGsnOZ2JKvs9v2C+6rNz
dq1vzmASugYBQXE0N1Pviow9MQNux2KZCRoebV/FYMz2W75+LlGmIz4QVkuEqXHa/MffI6dr8j5A
y4skuEJdUaHoMa4aTfrbIeZA28lwCB4qo8TGVteCbApqQmuG/kG/Faz048+C6uAsiyhRQxgV9sqr
ls4+s1biIlYjDCltcETh59BOT/xjPR/Rko99tt82C6gc+edxNCwAiY27x7pVGk2JJdPzpsOkGFGJ
HWrjLp7hRbp1q5hGwBM0m917yB0YLuuKsBYqAe8lBGZiyIlST8v1YvhwV6+a//WPbApOcnjEYRhk
YNIgszcY6LRks4n+TCQJhg4aUY6nwXYTDe9QFolBsfzo7qiMv9PqwWzo3g1ZgGj5lWv4azYySQ9Q
0+GUPUv6m3NwW9c5lAmxZYEvNIgNnOrhd2p27lrCj/+DWv4/s72TiwtjQ0HeNEQzpPZfirfrxrnc
uMeVTHIrdLynvAcZ536vXH/10HFHSL2OMPBl1DkdW7yYFQbhXhcPQmDo4bkGR1bmphFvRbEisRGb
llz1XnPKBvcOsidr+tcUZ4mndWed0GjPwRVVpU0qUHC2CsIj5DajDRbd/WSFTVAfjwomTWe1B+6f
Dw9W1RJehUy1Dyj1fL7IhdqXZf9mU+kZ7NLFV3WcxGvOr3HK66d4ePy0IDDYW1EyOhJtuHjVCGhT
X6DCz70hJlKcIp9EvzgYVhpQ9hpR16WDtKMGETnZkZ7vpHBcxZUxDEkBot7FHsPpMTmAlnevNnoT
rwHO7UVuCGSb/wF3xAgGE/8v4ZEtwDdT8YpwJ3FWUMtWLikm9qcDe3t68bw3ANeMxiYU/4kdctqH
jDCxgJQ9SgFcEwkySqWjkl+BcRxYg95PeKZU1iuEGReYpE5gDqH3GUxByiuIRMlp6BPLRjD/7XRu
UEeRSTNc60tz9+q15GgOhR3eg7/0/4m6IfKmK18AhpnijB8fPTtBFh9P8E1IIGuEbrzQBp8fkOdE
dW1I/zOqMuOprLpU7XKiKq/5441e637Jg9VDecUN1sn7ukBTJtaGj1WRmDljjrss0HZ9jvkFR10u
iRO2uV/ZOV5xkgjg+JKjftLFza7ip/4sQ0Fbj/1TkPQyNg36P1xV+gUnNxiuSzfeBckhixQM8swx
toYnwFJzkVTVM0gaa4aJoNRCzIRSJSZbxvoEeAk8iLo2DjCLwxuA4XYX6XakZ6+d/i9ueOWBFWyq
2FGRAsBYNHlCbxR5VElbydYg+iUNgHroWkXM/20wvd4fX80NhEBwHjagTs4KvEtqERyvHsiA5ddm
BRKEXX943H8z0jYavhVzjL0O9QR7NeVBxuePAPgumKmxKEEIdFpehVtTVq6uMlI/bPn3YFYG1gn4
j4o/V2oLriyQaZLA/331tuQJOLMJ+1IcnxU/dvTHBR5p+Q9X/wSR/o2NrCMI4jJF9qNIR9mJCZ3R
AlPwAuphmQS+n3xyc8NUpbpJLVWyQfdPJnvjndpgwXyW5KPKyCA9/FgjutUELv7IIuimd3QJ7WrQ
ilV+sA972N4NN0yVeBtpFLMXuO8Pn+K+21ectBP979O+LUB3eIm2nHidYHCzSB+3fCf2WbCatrPW
5yukDg5Z+Wdf9+jQvG0/HTVHVOemzsnibqt5Fy2oi+sxDDIgmsRNEixxuE+BcT8cgvL8DHyNRlMG
AhgfgG/P2i68nir3G4zK0Txe8KLqas9tFitzsBRQ9c32VTcUvtgBCWcZYwTA+Wf9mY7m/9Iv86aj
LuwK3wcxx8LCB48Sxf0k+ngGz90GXR5lO9KmLogeNVj7HWcfnmpaCXZZRWCrNWqGCRKpx1u8tY0H
4UtiZ2AqL7sqA5GihPC3hDejP3ZUuyJ4vf+padLZqM88XlHbyTVsXlQ0hTpXuDaahUllVHd4ksdZ
7xkaM2u2SuCZCZiX67eXeMBaW/FV7R0223rCTCFGOdZr3nDIDAMMrPAPaTF3vTGUVqD9JKhHdF1t
/LgpJN25IjCuKyZPKSpww9+EFVqc3evCLJddPD1cD3OuPs3WrC9NnWBRk+35La4120vk8VHJsoZO
cIuOwS6M8vTdMGp1fa3OM2kuJdiHTsOC4gxPjVqykuuHpLdIXdBP7liFGqev0zeH0SFsVBdT8bZu
FJsL7+RYWw/egshREovtBLnzZShNtn/yznczgIzBVptE9GvrdHiVQuJL1YYagtTT6d+jCbkhM6gH
yk7v3xz3U3CI7Gdiw5q4isQRZNAtjLbxaJTbd8bPi4mhltA1ANCTdWTUdyk727F5wMpCRoW1XgDQ
oDO5hkD0Nm1h3JTmZNxjz4cp5a6E+O/0Qn9hMmdh6xLMQbZEwi6LUTtdEKV3qbUx5hiZGyQbqHpv
vBRvpmVab6aEgIyvb2R71xBCHRh5QCb8qLup2zJTa5xtHZXpXGYrL1mXcjKJOtQK6nBzD2whB9Mt
j8htgCZUNZLQaUL66dRYI6sJFXfe69CEYxJsC5XLrijaKd/YpF7pm+wXFH00YLsos0iAz9ztM7Ku
J7S8TUq9JMUEY+f1sx7ZhtHo0aYa0P4qAnPY+SJRR/brjFp2zOQhl03SMyCRLumKbgMyrHOzmrjK
3A8q59hN/q9ZE3P6hQOiolnkiqA9ZZ01I3jVS+iXrgaMBOa5PHfY9kjlDm8LuXlvbCBHWoFsYKwG
XfJ3iH/12bKO9PucHKYNJc9aK0DlwY6qTOtvm/rqFUO3zo5n8QXs9cG4ZtAiwAefZopX6SLefkST
SfV6iLb5lud157EjR15bvlF4PbXd7gpn5DOlMlTGbfStrmpxPGQVmwByhzinOyM2UefOyNpVtPch
tx5Kdd19CedqFyIPvIGBB6Qo1NrxgmL53msFZidxXjEe2Kd4qeaQGg9TvOxXJyv/P/VDI1kNbREt
cFtvaSONW1srQ7YfAXo2BEiwN+hUnkIhuWXrnb2bY1SMIp/ZHo9Tclj/Bzp9Yl0TPELMT7PzY1JK
33joTeyDj/pZuyVgKwiZR+1kasE9PwZq7T0umMOC12rnt49nq5kCZCjRlg9GQkrrXE5sGa0g8SNh
d/9fxT7jWko3FXQSVG/kWk+3Jd0Vjiq1pQS6Xza5P1mEi6fXWB/L+ncpwo6pAAPZQu4QdyUFcGbW
0eAWVsJ69G2t477QeVHjYmq4sDt+P5a8J9Iyk68P3gaaY5DcmkuwM5XpILj7zy8NbVZ6EZlxaUEn
BlPd8pCN36rD5bRXDyx3MjPyhJXKxf8/7sCUCdZ8Nfwcx0Gmtne2CE+X9ifnaQtRHoiXanu/BtjO
iGCcfIcA/6cl3oOCO+0/smFIKzDo9X8K6OsLFSdlpjTGckUe9JrxxCKVzdxB8cGeesAelGZKzkTf
xc4Lzf8zpciOAjtNvYS564wt3n6W+D5t/76Nxg9PvZ9uZLHZ2yDPp2tPqTAerTsRSqBJB7QCsj+R
+63gwkPY0gExR+8aBCEJ6D9ojJnBtBZ66b5kfubPP3wBzGJ9QTS0DLoB57S0ucQ7fN6eUaR/5uNb
S3O4tOVj/h51DHfowXLEHs0F8Kl1ErGAwDJ0S6ekfbM9Sqck4Je+40/dkoz7+HKyy0CmK16sspGI
4ICStn4VnreqQh7hLNTI5SBCsJpgtHFhffy6Bq+tmVPzpGWqYQNcRlzmQMBbCUm7Jsiz1xSzGaMj
d7I8mKtUJDFaywtytWhU/HAE2f0vYS0yM6XBv72Y8KKq3qdjKFh11eTlXybQngAvOh+2Yvq9HTvT
uTYNvte8of6USaAWJIYSfm5hdmnGsJpcICpX8rzAhjlKT0YJQgxzIJx55aGMKpepMCqG1Itom5t8
OTTW2wWnwa7CRGDSyrimSGZs0NebeLI/R+mLEjbKD1FfimYpdJZT6zMNN6Si3dq3TL1ccC7t+VPm
kNStmxUca9W6fi6PRZc7rgXWJPfEjgbvybHaQ9l8IiplbtiBclQy/FAiuyoOkcbnjjzEingmmftb
Qc7lcvuKmtigawd3QD2g4mnga2E2/E/zYyoh2Wcow9CcfCq1Qsui4UDpYmIJf3w5+aaT5jNg8i5R
ZJMvKDUoWWDZAfz42oEFMPLmctMRWAfwz1GDNjpZjY/Beu1cwMuDK6qJqWrEvVRZlPRExhi7pxpR
LJXqTsR8awbNrvyZIPxuwXmjWKABN8OC0FurXkCrJPrwjLo82gW3xBmWYCCfLpoa/DmPspcD0UGd
YaJlxAjPInEZjKrWOAuK04zHDU09bdmdUHB5BE4XR7qsti/8D7TAgHFbH8kctQuOAlhS8Il/ZZFN
l3an7mTlKTuF70aOJjMGF3hAWtZxu9d196LUV/g39Gq6ee08gBLu1WYp3T7DQfxASV01aJ3ysX4b
/moCy3t9sbf0QHfaWyULCVht8WpJkerPwiRLKbXeJrZBR6zhLXS8wRtUKOQwMkXXi6gaZRwsvmz3
cyRcE87QTmz99X28Q0au57clc34TstXsDwZ38eESbk5PhnHKJbvSGVRk+Ee5AEXd688Yy99rp6+T
xt6uAieZ0GpljGJsLYnQzAS3X7CXA6a1vsleHmI9mwTu82QtUFTD62cUBLjN+qGX4mJDva1gOU6D
ZFPW5GRn0dg477D6bjy/pkaFYdJFdNlCsJR/vYaEwho4c57gOzf7LUenODK0ehDr7GhDPIdvwJ3b
Zw53UDi5tYEAIxRuLhrGvjeHIKZJhbZ2PhIzkjI1zXElMJdvknUG0yyDZc/+08MbQlxJJFsJ+rho
jtFaRpLXIelTJCNmG+Kb9mHDGh7CGoN52jTsu0NkeAeKeTEB8fxRLNqCDECqCbNKytTnaXpQiqZ9
j0GmaVr07r+ghEwlGksrsM0Zc91E4eJNmz7ICzMnPZ+dA3zVMAWxFm8ykRmZHMOOHvcZr0J3M2Uz
vw4gSBLBIKyYjEKB/8CRMoh+nOjLn3c5Z6gXSh11GfsRpbkoy6J++FdvcDztkDJvqxCMoWygiml0
qNO52afCx1wpNbuWOfqNE+S7VQQPSk/4fAZFAWXHjCxs2SUYjipdZ01LxBtSVQyvGkLps0KShmhc
THHUc1XM2d5OvutnuQ5UEuXZHxGCXyI2E+x7F1GrSojlNGk6hVRxnItK5Rz5IaqhKDtO9Pd+vprI
I/ZZi162diVf5mBQFhEVhQT2FGXUHk+FrVmWR6lJT+PBFXo9cbY6R3XCaIbeBivKvIBq0NHvyerE
LDa1VOKX89HOXLDN/0y8GLo2SZ69WENmm84ok3vP45iipKvewMq8Nk5O+iSBzhehL6pa0b/R5J4F
x8zObwhm6/3f08c4ne697JF23srQnqmqSRYokspbdvMZAIERILeEZMrdWs5RX9aiLcI9yl3ijRwZ
RHuqQmRWLHMwst95MJ3c+DUFz8fMBpWid+7A6NwsaCkhMbjNHuFFDb481qOhUEyr88Y8++nWBkDy
+n2npCrpcyIe354Zoh9pBrJGM3wPuw9/qk3XtfVDXzSfQV85WSRDZgbWWVamiCAtN+0/m3AZwHq5
DUhtpl8BaXYKfgTmAcBistueMwfwRP2tqwN2zfrDQ7hzM0RXBnEKhb+/MdO5yPZJSvek9U8YTd13
e4rLC/LY8gZGvsQZ+/3jtSMfoEdLKMYXq29zmnL9ReyMeyxfKM9gfXfr8ScLYybZnUfQbZ3fqOpX
LJbg0IFn3CxScfvLhC262Kom7jyQX5vJbnO3T7ZM9hn64YR2H6mTcfFQasUDtEDYd9zOWx2kJerp
tBQdY639B7cqfeKBZYdho5E7SoU52W0OSdWCE52HBBjM8IfftLtWJ1MShv20+emRoQ0nWtOCGjAy
X40QGLqXcwKqPdZ1zFu3xb4pVbSK61RAQVjwtswtnj5POFXB84tB2jpmVJBeBlw13NSnKycMFDi1
lnHe2q9flIwrmHYhsmeuu2yZO7IomznRFxltz4Kv/HPx4IkMZhq5o45nPHIsTFajP59L2IO86KV3
2XwujespfJVxpQCXvM9nGEuzv1P9jW+LG0v2wFOGvKCOaEKCwTVOrDYlOFjxUbB6DQnO4dsBeque
UFZKB5o1EoyAJ1HwHsWGLFKRUM79hz8dzeuzUC3JLzw2CknURQK4d3VveKGLTmIIp1oLes5i1Ig7
svLg8CpocTemFFQDYERGYJyeSqNZcVaQmKz/IXu7B5R0uHttZqq9ctfQKx1S3xADOwHd/v6ve52M
c/WbqvOau7QpzDU1SqPvsXzVrVIXvt9i7wNjGSzvd19WWL3oSGI1rzZizJYz+hz2QPk0es4W47py
nXtc0x/sCm1i9bxUz157A3WIkhuBTqDZtT+NEnI7F9zSpu2PFlh0KssmdzhxYV96eq8X4wAzTiMa
JMug19XcN1YBFHfPYbj+cg8OpIfnEYN4X0gBdKkwHRM0VR1xIb5fWk5DQEnU1FbQ6sZynq3UPdWA
FDfzMwaXocyzsoiBqkgAOUMQlXx2AWVjby7H7lJ6SsIsyDldQdZnFiwO54uP5W+Vop3TL8Q3dFkD
uVpp2US/25Jy9/r/jMnt4n+GC6tN7ksLObbmeeUlGIdlStmEALd6bk6In/Fz2xJ2KreNU04xlZOv
wckI93toH7N+R8BLH/qn66G60xJ776vCjub1CoE+LlczlG46zwGL2w2DSgsaKVaUB9MHyrqv3RWs
F/ZEWVItmHs/2TQ0Vv+24wLWy0BYqdaEUoub3sxC1FufkBoPF37CflWB+EFofxXZlh9k4ktu5+gB
SkHnvgNhDIuymFgv0hvoVYq06+HOdbJ32+kXfe8imHC4K/G8a/rvF/d70j2w2uaPfwxWpF7Ksff6
Y6vGMRxiPqAdRQJ8vO4p5Ff/zTF6Sfli6XgcAxWaUmFCvL66w+1K+7dbejZ5fsIOVNnHZd+F4pMo
OHz3p03qy2y6zT2MbDeULT7OdL+RG436mlrxlc//JO2WdpEwRFv3w1cnrQAQaJM6Zm7XmXZaz9fw
QpjpsKwUb+85FiLxj47ZcyPk9+r5VujIGU6hLB5CXhaHBC2h1983ZS08aq+OwDtHlaHXHvif6a9u
N55MHclOiuUqruF3KyYEavpIkInFze4yXTFnIwStW/EQAt0RFa6K2BHQ83gstrF572XK/uNDdNrA
QVNMlVvpTEaEMWHATT2b7ngdEXS8/+cRKYO3j3G1ZEviBWLUkeZYCn2azTLVlvyGYjdTKShkEPSF
oqNavC7TmvaocxAX5/xOKZ6Udl8vcHyBJkFiOwxw9sA5wu29dXhjU8KmPPrUx7QXYHV8d0wT7MVi
ZrN3EsyqwiDlKvFEER5yIEFETOzWfaJGJoGniQTgqUyk/VQ7HE+hhAs0iz2fxWwYm6xd2o3eDztq
s2aTqNxXcxIr2M3z+HrcmTlmRaR8QX4RkgeOFGgAgxeVsMUJTDABGVWrcpIafdAdMEp9bK/oVrM7
ir14lg6w7kuE7jZWc8sTTL0Uu1dCkasShvD2SfliXVP60HHGWX2SfIy46M8xQA5pkWmm9PmdcAmJ
5yZPbXhFNIbmFnvj+QVfo/Lw9ogFg8wHP5/LVYllTdIP9hDk1zZApzQpCPrXp+Wcxwt5jCycLDPu
b/NH9+I8wfd0zrBC3+ig687yBy+7OVEDveefBOtGd8y99EEdiQhyP2E3Gv4sxv1cVafpCwpxcp24
tp6A+BtjUTN6KUeeJEhgT1E9cmaEmjky1dJvCL2+ssWsfeKDhYqENCXrVvb3JPLvvH7woXSmHT5J
DAnX3VQYcHMk8NVHPm+2djsgWKXa10EmifkVfzY6dJX9fQ4DeB+p0raqxbU0tqLsjmW8B2IxUwPN
ZhsuSFOe2GhNRo/o4cq1R6iAorawvU0pCdsw+yvmGkwIYDM6lSKE8iPyeax3rqewLzG1OFNLpqK0
t5nnycF0R878Zkf+TNyiP1JIFc9hwklFtLcp3AbBxIVOEfEOKgGTyShF89OBYIc0DhEI3iTgXuEO
qL4tEXx8/qkK/iWU51G0BivP+/wF2NMfNrbJI+jWZtI0KTBqwGBaf2Bbg6UcjPy6f2CT/XrAb/ll
dN67LIH0TInuUH8iKHENb6s8lg4icDGM4mhqMbSx3I9cdWOpiG0nRz7//YkRzQq5+TIncXMdym4Q
7mtA4wW6ChcwrSBaQ72JkEBowfbxCIcW6A5+7K1YkV9mbUySnPFA8vw8AQj97V9D3Dj07vZ3cA4D
1jTCi8WtWw0SM4lOOUH5EljbVQ9vOdIBZsm7/xHLBKG2NskMQ5DbCbJVZEFL4KACTYsWi7H5poF/
8jOSC82jXeunMwMSAKeljAMfS7J0PdSBycCePKKoSm3SZygwr47D1V/+Q7wPg1EcaXCSr1nt0hn1
LncA1vlv+Zjj8VYw8gCBULuF7x8ApT3UxlYvNBg8bVwcM7hIPJQbFWmWWs5JvQeG59Jde5FzfYsS
NEWNOX9jT+z7ELNxfIjuTQajgL+LKOflYQcN7sfFEzevk4msgrr//Bb/4pdImNppSnrb0eMZ4uQV
yJaMMzOj76gboPCeoAAuJ4lsf1CL/rSbf77sdsLvzZj+WMzwYEz0HiV2daVdI1KB87/SWk9xa1v7
bQpQ15PeFd0j01j9cduCMlu9SFgI8rITi0BXX0cqVvJZO0EHn0e2r5Ek0hOEM+W3xDtNQYDWh/gO
K2hVOHBViNq67nIWbH4dI61tcY6yCaijDgM1jSUd3yiN7ebxNYoS3EVHxOcHeJqcJqa8at/MvCFu
C1pVz63o/5eFD/siJmK6uhNWKV0xA8aX5tbrCTf9481O2KvTsmtwxIn7MVgZun/GSGPl3OmEBmSO
Z9wRFNKS9CSsmxDXjPCw9hOPZq2h2anKhWhEDqFl/4XEpdek7fR8SssG6x8+ZhS9mkHFzuKW1bnW
MFW/Rm4qk7LN9YJg/Bf0Dkd5phaOO6pOFxFfGocYsOW1Qxsf5mOWHMu5H2eoCghxEbZX4pnZiWGj
ctT/D85WzoqX1NV9xjNCpiH/e0R22x1C0qZkKuzrIGkawYbOQRrZK6bTKlUw5ghYmyeGInRpQlxP
sZpuCakBr7reN5afdol1ijwiaPrMTn33t6QCGYpuNl1AfMCYUuZ14ADulqtGnHSiTp1q6AdeFjFr
s4FrGadKZu0Yb6yx5SoUeTmSKlQNDgT4w3+ahA8InkGZr21H5iwhjiQeoscF3bNzVeBUYpG9GpPs
Whx8AoNu0TXCewYGU8cNHLQkzofU9U+JLtMFWpRpb3h4iKbVLdf65+OWKlTQfJSqj1J7mP5IeOUX
SF8ShvieMQLv1pwJSyepluMKNDxAisO15kXnDROyWXMCFuXtuiQQXLpEmw3RtGZirtPOs+k0lQs7
HBLuXTKIUp/uGtoF/4eM6gmujpdGVpOpvJOJ/3bWLyT2AwhjKwpLB00BfYdESc10NXaTgubLX68w
SZyiIm9IZ9ArKXVL2LR4YalluHfObUU7ykwWg1SAerra6DfgimNvZ2sbRn3KIZdSVf3hOtbWQUms
14pXMVPrAEu04z9ZQyYczI5AaVNa0ER+T8+eGSXnqyJTMRhNzmvyRjzWp/XzCzNw5pRz4/i8RPDP
FsRSDlF78XHqCj39IO1rjVXVsCJ35MZ2WHg2rFBim5jKOVJVb41+sxQz5qO+xMC+qus5ZXc+abB5
D0vmVOMHXPDzpqRtGdXSXlm4DK0x4hspDaj6WvYfLEDTAt2k/D+y9jdy4Ob28911qgBkkqkpE3fI
Dg7F47+3ZnDoIRq9YaN4zaqa3diy8fxEDAlvQPQ5SnhaDaUjoZT1+fFhqVGNb+k1sX0mAdnbJBYK
hgUi3Ucwjwzgp2cHk47jMeaGHRmtOGqWnsHWmOukXRczad0nfJeKQCyi9QemzQCiiAE7+heUhXGN
6gJEz+LR1z++pnSrML5/YENuOZ4N4/oRy8lr1Mser0mGvrftbR0PGU5jtKoB3A9dTtlSe7DUmaFP
gmdHrreZ8WUZezHxRdEGNjUiV9HM9tpFFRWSaxpoUrB1LqY+pTLr+dn+60TOnFMFouRTGU8+B478
lSOT0+OK7tO7jJfidJZ44RYWRBGyYVl505Opbs42Bz0logyLQRZ4TXW/E53U3CklRH4+biUHeJGq
0/NLAO4Klciy+o5EsFFt0p+XoYDUGwawKd0JViQh009hyMDZwD5ELYEZMHyG5S+zJwh/2FYcIbrH
8nxqkg5t+vfz8ktsS7rO2bkkaPe5doxtGJpbis0tovJfdAO7RuQl/ls9e0qdtn2uoUQDN0RSqSj3
UXkQHfz5w4x6yNtlwjiFy6wRh9pZVIfabHy/Yishm3MCITK8TyzYapsPY9BBdvDvIKhsOjB44+2a
T+0GC8RIwQRU89v3tTvPSicunlDlBfY+SUipdA3bdIkGdcIrjRB8ZrqRnNRXnyDchf4CQaEQ9agQ
21aXdOh6cdtnbGncHbU7ciPbIf3WUeAyOPQ9QSM+j8vUoVdyuXC+04upfUsdADRB7TQx1V1Z2Fo3
X+8FN80m6uoX2DzEoayGwntIdHfAqtBZOW0kpU18AVZ64Rz7M6tX06sUIOjv/6xQbb6ZSUjaMM3A
N4nYo1vKOi4AiSnRny46rHj9atycEEi+0LYF+8vEP5gNBlrJb2onQU9fDhQ7Q5NImP0zzVM8oSpq
2yhdxVvNPisStLk0U/2Jt6KChb33uOEPbezkYZwFgVuJM6dF6tvw7egxeS8pFvvWxX7VUZncPYIX
BjyP0ogdnGU9wmzHbNBmJ1y+BAyQmAbOWUdiyFSCVv2uMxkbvWT9XD6gF1jgua+Y3xn6/WfjwPGg
W8Ep/gsm//az1GZXSp0jZkp6lrWZAWs6ABYxCrquNBHx6JnaY9vVi0/78NcaY8fxT9co+qG4r/3n
fUaSdxogAxDd7nBBeg6hHe7cVvlWV/FfvDsLEJTh2t+AO4ByZ/oBGV5jT0uaQN7nkzmgh5ZwpqXg
I2dDsmnLs1dN1eakUNFU45wJn4WJvZ2DtVqANUlpocvbIrsjRzjq7s2fKE/wwe5eOKM/5J5Qn6yP
pkOkrv5Zr+LyP+oXSAI8voAHkfS1VzWR2f+fssZj5wzY9CZOAgbHjByLYoz9Iq52/i6bOLeSJtzW
ilwlPpoN/JY1r3nZMvbgrn5mYNQhyD85NybpJLSVbBin7U/P+5WOGMOZD0eRe5sCBmChNEEktsUY
Vqtk7vi6lknGzqM9t1DrLZDQpjgfukP6yngEvkkE1ZzKKZFFy4ChNIQ+eXejwNmgFh3LVnTY0gTx
r4I82+sX49mqiyo/xFQmLr0S2hMEeh5wAUTWaS907fFZ3fRwh8TTmerBDS3pOPpT7VtCeWGhytlw
oTQdjQC8HfUs8Bvtgj/PSNhYTIqb8IXL1IoEAGAzMxzJZtIKk8/WHTdFD1ZdZz0To9tc+9rz38w4
cWtLo4mHs9KXZyrbERIZlek80QWIEfnxmwpCrr8kPZsCS1yTAl58BMzluC/MfyQ/5+hAua40cT3O
/MQXdkIAIO+3n1wrU77kktcHblpHRDaD8noC37YFcxykmUSb82r+FU9RRepLvuSEkgbaSsslD3hR
T0hER/WasUCBQsR8/0xWDhlTljafF0vVhBD2omTOAhtpLv71+YWxjSHrmNU5p5UmU4h8L8feG2M5
8hgD/oU6lpMgGhMjX2RUfphY50M9D8ob/Zg0iiHm7QtDTzZydTBM+XxrXu5r1lb4kSSaW5K482gJ
efrNXhncxuLRrybUECMORC6z3+4dLJKeCwQeWtwVLunMo1oaBSfvZ8SByimZVvqkqAt4iF3rjkIs
729FQnXEo+0jodOQfHkHTQjhtUmudqQCybNNsbmLrcUdbVNWqI6jzHhMEouyB2GoJU5TvEStonK8
b0xi7+m4OErR4ZCZ6gixFoaBYtdLqa/XF4dlLw4s93e4UEu6Ea8yXa372I8XBDLp2OQTfZARbCI7
e74CxED9N2nNdApBJ/4paEY3+NYjwUNW1rlczz4FTU1sVYan5FmDxcn4ilYDNn7+B+HzCGRF5dlB
+wcPT6tRZ/RM6FqwW5bedz3yh2RC/W+PIDtEuGcC8ZGUOmz21JGzthCFWsjCkEqwsoCGu+bb+NnL
esVXSk976bBfjrH/kr3uf0vawVdDbJ3Jyh/5zihMF/n8ovTIouic0pxZSSaIOltoVm7dfKxLwkQD
DeACzV44gxE6U8CEtoWn0N3lFfVhxXb/LNzdEOO3PyOQqqipw/0WtSgy3jF97CVdeakhgtcm0HJF
J33r7QH+sXDgW4I2rONrUHNEqEDgJw8xWkuOX5XTtughafJgsrOoDQuvXfqql25s3j+Q5mUDOPAN
hEITsEoYPty17uWPfje/lNcX7wHMXqLhROF0PylSMlAtp02dvt7ijJY2SJKj5SQ/I08LslHnmvJ/
l+hLKXF04ukaCjiL4/kF/lMh0Law4aZOsqjhOreYbHPhyNxE8LMRZOospyfRTEOHMefIdJ1Q4Ddd
8pL+QSaTjTc4db3XiYUbAXSk41by/XdtRj1ubA5hdPSZa2knzpMt0ByJYj09W0BNjyiYlIinFJlb
HqKzVRKQg/vJu9AMxZiH3IGvatB1+wZhe6YAMsWqKT0/VuERuBahB8qoHnh8FcQ8dvBET3eL0hKM
+X+JDfUyTdx4O/EQyzIwWLI1f92sfZhYJoC8TpYFgcDcmfe8dK2OpsOPCi0bTtJ1HQ2iw5NiXQmf
4okDfkdhMahItmrH5GJaHS+EdkRV/QhvBvZ4Y/QM3UThseRTMUrkbeA5OY6GDs+a4oyb1yAjVQrh
rxT3u/CtP9UUNnO+hHffPEG1I21wkU5sYmFzv0T1tvDd8ErT+aWlv0kH0j222tOBKXQ/45o4j84M
qih4eERZs/IUvgskOjBCGb5u/KOz6PEMIu/0q54R4BZlHyp4Yi9+5qa0FAzr0jbDpSBowV73e1io
jcFvITkqnR0qBOVYzfkHqZWSQR6FG4U3ZngefUKP+lLbwpmnrz4nE0FQrG10tzvu4IRrZoMZhogc
KbNeFJxYKUsM+ZSbQ0VWWF4h2rEULrsierxMZMoUpOLq2PRZav3Q6Dr2c21biOpRDMB0J1Sk4qMA
UVhL2b65EAMlmvUbQXW0jYRK0cHVyFhrpMEkMnznsP0UZRbkBkcrrpC7a9bO66MSdN681Zwzrh9w
PSWlEx6eHMMiPwzGvGJMRu43lTFqLHJC8aI7aTXt90rR0TpjYcaAFcCuSafixsfgsP9kzgGaYLet
exFmsw5SbhprnHOLhsax1HL6d+L0d4rOUfurzWmii9IChWYw+yDQgMv35ugWXBQNwQat5WUh8wao
M9/5dMwbzfV7gll70LmgKMS93vAnRybN7fUweLmDaqfNsTFHlOZY3KgSxfzDD1p2p36ugym+2UgX
kJzcz24XYHoF47RadBtdfVVcU0NqY4lT5tdBgFeeVb2RPSMDE7EplZdcsnu4IPKkJY8lLJFEd+QQ
LzBZSESRNHqVcrDc1JrN9e2D7CM05efvb2xnf/5v/ysB3jbRa4CRGnLA0lQ6jj1iXJ2HEdRrgfHF
KZ8vtyzfT8u40z4MZvhfUudQyaQNNTt8G3ZoAaKCyxgp7/4a1mTMHmWxUardPIWF22hyPci4tDRM
u4W0fGvruF3sexjmEKqni34qce8ai68TcuO2FAwxH1iknyRoptS50lEa41i4xWDRXBuZweqjJYwL
5axmVJyaup9pwHLesMv0/FL5PQGsr3lgcJW/xD0NdvMfFe7OAx3oRs7lwzg8TozKlYSxaw2WHX0U
1kL14sb2nOB7XoO85C5DWmRKPJhRdkPLg/7uBo7zvwIlCuEL/vBTAKXxdfLYDNDAfg+dFQRJE5kz
WodsNyRQ4tAlf4RyrSfuIx8JGDsvTvCeaAcFROvBQ3mj01EmRV0D3CoslylvaYyRFvN8SXkT41/F
xmPwngkG+DhfeCGtkqr4aB1izp3Vcg6cfVtMiEBEELjyRsNocvBGUM2wBI5jfKx0HLeSIyU06+J6
QVSRMxP6TFsZI7r0gpZ7pU1rVdnox/qwEtZG5reO6zy5e+KIOMoD3kOuE9J2oKFU1TixRYI6mphe
8V9W1BPyKSAK2UmtfDoVgysZaJ0iBKpwu9DD2q94jMYvZm/lMlTeyVpPuMfJuilwzGcMeUFNixuh
lr0DyUqT0xBPrPAQgq5yfU/DeE2To3R/gQje4vSTon+q4BAxlDScuaB4a520TRS55BwFzenqbjBT
MGDE5USU5v0+k7D57Bj1GQ+x99kc/hlUm/FXNeh3asCkWvdY2SQDaP+zx8o3kSg64gDajREt6U28
xBSa2CQFpkHqn9B36C9TEv3xXQbKiN4hYx53v18Ey3pnjAi0ZAaS/S1RzCMNJbkgbWY5wLCZ5EHi
lh/qfNIhnHvdK/7sXfkPs6I55nO3XLHqp7ommwVSzOoZB0DJV5j1BNyVh/qKzRrbyFvnl2z9p6/H
mHpct64FLE5haoiGAywxPQBKdoYmBAvbXzUE29IfEIrix2HKUWsWfF0+/Q9eOrAVgfskfLlhi2jF
Enamj9oF0Rz1QFO3asgTvODpRQ1Rsk/rmS0fYzFew7SEg84SHPSlhqWh88+oY3QxxLavOZyeoTQT
IIdP9Tkpn0VFG5c2rHG0F2uhl9185ho/XTrnC5Zktz3rpaYnnGXh0OSm981HIAgNYlFajqYV2DKe
XX9Y0je6lGgWBGP/SJTCaQZnOd3BRT3LYw9ZdmtMvCLN3uaN3K0rZbUWklcvuA+7efrBJLY/1TyU
eUTEQSeXvbQGwZZgYG+ebsuBts4LmfSUVsWTNDRVWrJt7S2p6ZXqKADNToHOz2fivfkShne0FVlk
CmBE7NUd0fUpDmc88XQoDit8DW86zivnPOGZ68vx613Fd1dBVVknQuKOa+WW+SutC63hwBZ42Tdo
v92BupsYCeLivXBtkoyj+HI9155rSJmEml/pThmkjZB6ADqs/d0gIEDnyKWRKek7nrNEw9vonsS3
LL5JxWX7zcCx4Ros09PF5V9OaMT/p6KZyur5R6ckHveSejizo4Reg18fbolaRTgFChf7cubeOJOU
TxLs6mjLJk3M6VUD92zP03/Bw4iLsQEydjn6bbYeX8UUUNhJAYhoZMFQzc4TvR9Znb8BrXB1xFeN
k61OjqzOut6o7LC7RldT8cyDW58VKdrj6TD/XufrUbLYbRWemBdxcsQqu0eo7vzLFiTRLpR/RiX7
HEXx9wNfEqPcZWPnU83S0rmvUJINsUk6xr5FTM1MHTqwAq8/UY3C5OrPK4UtmKswQmlPcdp4xPhI
eC7ULbGXoexWyjYw7xWecFvOmQcIhEPxuSg/FnX19p9YSnxE90+DgDgJRla8eMtJzgqOwAYiPdHd
YZQ6gUOUvHeztBGqoEy18VqMC7KY8Cdfq7yIzH+STmYtEzgvg+XPSbVR/3MG4S4nsuOCMOSVjXIi
e8d95B5jhF35X8st109uUKNPYs6gUROqLf8IfLEGLwwLfszXvamjd5u449WA6GGBkThzixBl8Mbr
6H5VbJEmCLQkoFNIIyOZ0TScCSrQpc0vfZycgG/Y3eKxZfFXf6/aP7EDjV1do+W/IqrznmdZe4Lg
+AlaC7ymXysSuYLQ9wwcAyGMTwJlwhJDfQEota39szYaTYCCeiXc+EjV0zmE2rLz9O7QPoW1V+lz
6BkfQDl5DewDyhaYXMXvPj1Ibstmk0j9NHUor9QJsAbqoBVk8aMux9wdG5A0eR78Q6qCh75Ri2No
XP19u2cmBIzSpYLmbAeH/pZX+AhqVSanBrKgcV8C1nVxcd/0zz0BPNMJTlVBu4nojZ1uaxfRi6vw
FKdlN5XVyYNqI/u7Dv3rlDaCpcpHsCgwzHFhnUer8JE3qUKtLm9/8ikD2qi2lDQXVFkL1T6Vjf/b
r/F2Rt65xAyxG8gf0xNwFq7UL8M2gdI1uwtp1dh1c/Gph9YDnyUeW5ZEdBOp+qsHb7qnyOH8tYFo
R8FsEHfxS17V1mbqJ84hjOQHbaYeIHGKoSArRtdcFp9mLed6tHBHzxrTqqrltXN3C+e8HwiW6Krp
lLHMy8Hd/QhJXH/UZwpAUpo7BSrHzZOgk8LQMedmWWFpOa5/7vO+Lgd+BWhCUt7nZBVgTmSmco3Z
AZhNMaqkyRxfNtoVJ+tBjK8mOsXEg7vmSo8jML/5q+wN0ubJ0GPWxuyk3YPXTSVQ5GNHgg8vDEJm
VkTPL/55QSZHt5ROHgwN41+92MlgYh65BYV3Ycs3liMNCCM2ByMhXZXlQ5olgoKPXt7N2A6RRcnT
11ylbJsiH3BBt/HyeE1NrAUupKE3+VxemEGOT3tGlkAo2DuXDoidYZmKR7n5ld8+75E3a7rD8VKa
rbCk11YurQ393YlFnl7cjcGa05tkPilUIl7hmsv9tleXtONCgqgdUoiOhLKl7N8C5dhuSwTUhkZF
wSJZbwC574LZX3LXC5PNp3drkWvHr4Rvv63SWGqrqQRndLpsfZeJiALbIOnK1HdnRmNJCPSP2IEk
vsSGMK+99BI+kLYn+7jcbE1BAy0hN93qXQ25aN6iBKZroKinQfnvIruolXqHySee1d+k9x2dsJ/P
KwupX6zoieldVnkzhzGfy6dzQT1fHfPMXfWR/HagnbKMQ4Vt88PlPYK1Kj+YejCn90z3fz/vSfv0
WXahla8ff8XN+RguRFk0m0cd2yCNlpphaW9Z1SMg/4ANU/Cf1Cc69ZKtH5T55g0E/z9A46ooQ1S/
ifGETCzSHwqr1RH8iOuli+nxtXHRTTRfUw5Vg1yxivt5eYDDaNQnvScxq0UhlxrmV3VLuUPfscOe
F5FeyYUOcvxqYiPFHaBSum4DVroNIyk2gS+IHQFSteqsLLi+J2YLl2aRlry2eYpdDBaOEJBXiIJg
Qt8X08+xWVeN71Rdcpm16ufvavf01EAXZsGvcxZcITf0thoZN31eDz3jthgFEMNB1zx0+yVuJtW+
cp38q2NOZ4nmO0b8vmcqQUySOvnsD5uTHy2OzRCUZcdWNTaioIBU9Bj25k8JKpxH16BQpJqmq7Du
4OwG+7DbTaZO5SkZpQnU7FXw2SnZDt14ax6yQFDzcoBaD+PUdof7R9tIXlpxqc5R6vC7U6xQPcCF
U3ilE6p7+1Wt1FqsWRQa22x3pFsni+0/s/gXNuyA97KoMDEcTKJlSyVj48rb6ghSXICINqeYhx/L
+s47nKEeiGEgVYbgWY6npRgb0S1q8ucxaxqDDGD5BKM8wqCASQ1ofyJUQWxAyFA0DX9wnXwOcr0f
zNFjK2WIMZ2eYs5F2B0oQiUQnOrNRLIIVv3Bf4Oifb09VwF3KlF+MG4w97Y8bnZop9KjrclYyUWL
02iD3BHjoyL6uz2qAfh6S2IQpCS5u97mGBz5b5aqlDmI/Yci/X6KUgx1Mkr2cpTO8t3ozt1I+38R
aPIlro0Q+do7qe3OG89XtsPHxp7Rj+ynM7VHKtcJ0cNGmumN3mrRzvatosHU2+EtCtrvaR/gFpZW
r1hMBVwkc1YrKSdjRzxSic3n0G3UY1C4v0er/9QWit9u3MtPBYFQkTM0HDrn6lZAymQ9RwkgfL+C
31MxE1V7c7thtpJOiskpUcOM0GpHL42YePeoSvQH/3w9OnyKqP/WSd3nD0KnS2+pLMxNZF9JwCKT
WLod8gcFUqP+dIN9T4hix+6cjtCuSSPqpjqVsxdH0oy5bOb73OYx24k60+ndaM95S9CedOqgBX0s
ctbbJKuMAacFEusTi1XDL+7OjDIoLNPO48TcqZENvMtpVP7/ho8R/Lz5ui77lFKMRvz/Akrodw0m
/xtIJ2plsIThn946HmwNM0XSXh8J9dZAj1DCtw7TYpYFrnFjBl7xunbhsOOQ9zuBgsdLhASn78ll
ySbZ/M0eN0w30jXG8UdfHH6S4LzMXB5+OHL9lvQsiXTHQa2i5aU3WorhxOQWO2hYOMNH5BrzvUXZ
juoZVT96lgpnrdI0mYb2VYIDINyER2sWECn8uigwmtkYuefEfwbSgGICRuqXVOHSik/c/YcWJ8Co
fmNNAcId+B5efDVOKwonx5ft4Fstvpd+rJvDuDXYAK29WPKQ7IFOmbCsndE3aK5rp5QA2lE3ml9N
e8xq1e9OslvqME2PkBmZC7JS7vzCjA2C1cady/dpv91xu6wljvsw9oqxFcVzo1qLqqd+EulLcl+3
E3NzqjPqIOzMo1TD0bHTJ/8JxfXZDMLB3E8KOWL+0t+NXa0DR8UMobBW17MkaJrTyRdovpnBTXai
H7y5T8NLvqsTvf9EzNVjK8vCgQIINHsaHnJ2ijqlXS5SCba346m2RJRNLdpLTYaHGOxMbObEQjei
hVA/v15fYiKS19MT8fiJn1VHDxRSZQLYxQ61E2+oo/nP9M9LnuNx+0ebVehwuhmuwESnDAR+oQT9
8zzbHsUIO3PxNaBdZXsNy4CqUd+MZTn0PdE+ofdmmT82MXZbZTyX5dBLUXAuq5MzADLzg66XF3du
qVBm9GSfBCeaLSd+lQZacKnWHmMS8UK5LnReJd9yoZcfOVjvolBamkCBZfmBs41MIw0T/GVD86T9
BeL5YJeb/hvsP+PvypS622PJ7t2D24CvishV3ZlDrw7WGBcnvBDNg6M5ymp/4v81ocucjm2O1epk
XP6VEyyS2X0gydxQRGPLx69itvlJaa9tKO9avdXAkUciOlfnQ9HBzitDKS3fNcmY8W7F4qHJg4fs
2A2jBEwS82Gkt1VUCs0m0+ZS5hxhxK8XsDQkqh6VPBUDAcYi3+MuoYz90yPOAhGe88SWqmmTqYF+
fWjHcRt/lHdFldqZwN5vv20VoYKIjyObl9qv+K8Nf9QG+H8qZN2UjpPKmLzv1/Q1VhDULBhteqSH
TPDDwHAsjDjw0bxYEIoNkYguCtoL8hJipAMQr2OxXJZDzzdk2ID5e+YV2ie4vJnN3J+1CenhmecL
XhQ3voUxczWnMNcW22xGHQmZUfjuLV4DPHKQDj7O4bTg8/DJOOOovmtt9Z+omx3AfQS9l3H6IfxB
1YBeSPDSGnQb9BoT++u0t0du7Y7eoHCY54gS76Ct3Wm0qkqi4wlEhgszDbqv8XzkEAlmEgycciyF
ZNxmXaPE1XkNi8KswJFcPRBqqASsNOmGRuApbxQdZydkHc+mfdP4Pd2f1lxSradCy5HpfwVUFrqg
Mcjj6CXGVHf85M8D/n8dHgVdg+GF1kt8Jk4dq0HvJEbqlk7092BiT7WIvgS+XxT4GBS+YwSlTLVu
YMktl+qlqFROqkfo/QgodUX9z6rIUDSMd2QroRNCmIn0P9y55Ne+R+KidEDtMB9NIdlt74IVNMQI
nR4zHT0waKpauxXgYiz7OdVvFzlHfC/p7t94FYE3xnvz8aray6lcwV7Bo8wB77zg+/LXFjirjyUG
g+4WgfHi4p/2z4O7Pjy1yIAlbBOoOJdf8WCWu/c6Z24UviUHg4Peh5iJvDp+NEEHJqcE0w6NUK6f
N6GCz3E0eU94vA0zDp+ui8kS7+1js4f4z76LRSGnO/kaVjewj4W/U33cPYpi7xJdxipUPCQFrRWK
E2mODve2eKkJgxFO+L8aRv3ER+3RKPMW5Ixrw2drGocg9XzC89vBdarlWsxtoE+2Fs2lv/ZlOinQ
a8Oc/59Dv21fxvkdfRDjQUh/OHIkxhMSWmg4pHAthelE6pdxi/xPkfnpyqQ1yudDUykaPuEB/vm6
xdcnKeWh14FP6ExCuPoAK8QnLhT0dK28J9vBQeHVEybrzrJcoTWkhPJyocE/lggu0UWGOC9zieku
zr2U887nAhcROaqyad8Hd2PCF8z88qsy1+vuncTIGsp4TQ6/7W2O9Doc98EKxrjjacUKyj8RMtky
pLbBzCZR1UH/9N09xvrI0a1G4YaK0q3EIOh6M8+vtdAHpDZlG6QmF244bVjeMvabrDiboJM0TyPX
kOro4YlJz4foJABn+j3chrvYlS8Pitj+arqWlTnJCWmOIxY4dob2XZLqBhOAgTDpE/mJUOO36v5e
X2/dMt2aKY8dJ7rYDQwWM8eSu5hY9y5Vh//yE2EBten8oTn8DMxIOeoKf1ql4IiSznvO/wwT2IZk
Hz8iw3uNKhz9ojB3pQrQdYw1W53OTAlwz+K72lXUgQxydgQVaj4yNNZO31GJQiVuAngM9rTferTX
3FCSOrgw2CMmMuYNipGFkJnk+q7Vol76giEyxi2fjEaxXpDljiuzX1vfnn2ipEdrRKivUt63xqud
h16hxJSTtT46bdmg3txdRL/IVSBHCfHKk8gfWkTPBA3bHp59HNf8aZrybre9jPtcwLwEinKUGw7n
EGsuINLxXCyEJGV5Whrl0MQkwbdR2jhtAgwJY0E662FlyY/lnwHL573tqLmXs25kQJCj3Xp4OYPT
cm51b6u4ZsdG0tjLergQTXU4sMYpmhg8s4G9h8jK42N0VX7thCHMdE2zA19/gqaU7nHVeWvQNFK7
6i9peBd+ZwF4ePUqYMtNLBeUjKnMYYI+xRh1fYjgSjSlbJL5HxtcIBmiPE5o1BL6yb5hO8aRiJhV
F4oQtFCceO5M9GrqRamMm46Zclfq4BJlpngNXIEjqb9KJYuQrYdpy32h2nJ7VRKp7E8dRvB4JIIW
eas3m7FUyebPv9/0NVbTmY7A0fBu0SSS2XSoNPhMR/r8mkSrIaTEumSy83xdsSbwRuQbJjHpYMS6
2zNdS3RL67r0lQvGpWulVDY6A7dJbdAgiR9CtM4ZFrQWINgf+MY3uFA8/f2SYqdKV2KLigUi2Igq
0f1t71rrn6jCIWaxSYXghGm5lw65Sgeh+TRvcGqoZjr5awfwdEzbqCnK8ZRzP3smHzwMZYALziuB
MigPU+QzK8hOhWKwhM1lfCCtRruBLNvWnxwLmXnUfzTpAtvhxOTApcuSOfrrICyXXPWs5jCIVOhk
5ND+V7Vu9hEp7iMLIelp+mrbTU4bwZfW/S28Rg2QsrQF6iB6kPHwYgyZQFu/6VdIPoDnjJZQl5VK
T6a4mAONEeCqfuuXLx7ECuD4W2nJ9hFmKvNMURnM96jpgSD4ah6PvK5fRoih4Wd9VxcY2aK9rrRY
x9ahrCx3/PGPP9/D274cJZbHH6J1iftgJhWgtWmCJu4bT41KgoTwOdG0iebF5Wu9qgSB6yYpE4/o
4G3DMdEzkS1E5M8mc9gX0en05nsvulqwuZtCD4W52wHVhOcy/N2C0Cos/XErZwPq0Na1hKC2Xj/q
IjAOzbXiNuYaJZFANAyJav4gT4lL5WU3sIHgx+r2o3FfWpkWLN1g0mjn7E02HNEPlHKVILuaBldx
Xv8s3gEEDhIiTjQ7TdM4eIe1dwAEul5rJ9oA1ZRKkrskzPAa4aNAjZdYtzMf9nZpfPr3k1ZIt0kS
4xo+WeiGhIg8Ik2cs+VYqeSFc7gmAz6UgV5V0feM7wWOK0zy+duDEMvahHtNX5LVvuxa5oTbjjXy
9ipCDijApvtVWMVNzDHSk5xUDWHaf2mvCVad4DzOZ9bbSzm0ym369nwtUeYYg5YRSOLdxaDwSU5O
vOuwcTVeSModOFGEkfmYxl6v5m7pwMimLkml8wpUsdR4hkfmHUzDda1F5OyEtTdghQrAmYt8E2WD
AxF4fC3lcRUlzH75dsMjWKwIdwyV1p4NqzISNQzLim2wWN15gSComnEjet0J6aBRZYiyUMSudvHn
uyNr05NQa1x8zmtnJBN3Q4dz2z0zC1LJb9r8CWvY0xrh1ib1AM0ylL7yqo6TMyRumLYeh9IcD3dS
3vjux7BOHe/1ObBYnVldV7Y2SLx66Df08BkkE7rUfbzyydchPAtYAUB2rUjCNgcaIuR3qDREeT+W
yjzPkIEU7ApXj143LbeykuvefBJuDuzH+Buccp8SKF6SxbmCzoc0ECApMaoizDbBMrs5+S2FJu3X
UD4fVEMmxRoB58aHH28sVIK387srnJxs8wSnQVrWdF6GpqsPII1d/8kBRvPnyIDydy4N0uR8aOwg
QKCllvNKOv7We3ewN+lWzL/5j+CtyVpQOvo7+NvGTs/cuLiPr1fE85SZm69/Y+6C5PLQwarieupI
aafs5QCcQUO+WepNRg0nbehZ3p0reQO5dBwOEM84wJogt1nYFxbgTzf28r/h9AzM6DQV1dEZvQta
QcM5e8TyL8VqfYEXH8QXeG6CYoGs0+Pv4c6xCmP9jPwtvRGd3sh1In+1J01tKtZhjVjtK4YqGVfo
zti0UV+Dv41thaWLLxM9P89HE495G1Lds0y7SoklItksL9HK2H5NfbNLOQytqXc3GKXW/XhCv4TO
5NxmJBaCp00BZXPe4PuKQhiQnTNnvRERP8zKZprPuVuUhYRW28T8huzUwD86Teng9y1iFoUHUjCC
lpl22f+8e5Hui8u3xAIj98dKutiSUGkBTWYrH8oH/ZMZaOOnfrXGvCtpz+7WeuUUNibP+Ryc4qUj
YP4LhtTqAeSYdio+2S3VREG5ZHUzY2qBDMXQZ2/e3Dq+c0O/G+dLEeVv3gGh6kxFKvyi4TdQ4J14
jJdJj+jXjwFdTqbRrFb+JNNp/y10ZVYypyBzb9lFKqrWgC+UGfmGYoV5ZZonQKuLCidgHl3s5Deh
JEzXmCtNJWvwoazeRWNQFZeYNf1G/aMiPqL0mKzMo0jRpr65/cj06UY966LdqyISR2ONAuHbWpq4
U7eJDpccC0rXHaWIhb6wcYHI0ihMQ8y2EWmMAodtPa2PsP1xlUr7M++eKY3TuVdSPVbOKQ4Exgr9
dFw1bgswD0OKy5ts45XC4OUfa2nbMhPyA5N6mVAIv9qF0O/Mm+SAgdFVpTu7CqK4CAlblBiTfxoi
Il9H8H/8OHqK1zCW/TY6gWyPYgd+Mg6u4xHknY9ZUwflusYK5xQOVvsViY6toyYjk53YUY8worgi
uQ4WMXqGY/+g3E1lEQ4/T9cMdwun8iSYlv5oJ98kw2Zmo/yjS0fdqJuW4WgGl5PN3Z1aIKmCUEFW
smidkR5CiUu0sYt79bcT2rrX2mxyW90QVzx9SPBMwD8kpnYLeWshlm3CYKLj5Hgt7+YefdsCM2Jg
iTvrJrJ/kbt/RREMzUeToScwf11fPVywH+q2wYLdNG1XPjxMeWRx9U0lYRhqCAseQb3jvfTOU5wm
I5GQZOOlEb+8fXPAUs/9jhvqmjQxKvr5jGnkwkpFCElwZdL1HxIR4gZ9zyYn8uUV2TTjjHJ/XWcB
6SWGOO2zZWEVPFOvdghEU8sOw5phdf4LXOL2H0qzdgWQlqkoZW/8k2ggFfR4J3jFPfQoiTO8UA6J
OjEagN5ZTq7GlU8UP+mBzkRWfFK2YjOzbf/SAvcGAPlMoCNEGQDKHYUWygizjjkauCC1mauqKin7
j6AJGGFwz4nUF7G2ndOK1tc+qvbl2Y3+iwBjYMWTSlYf7Ypqf3Tli51U4V9MvSc3hqcWEV5/7/3N
XAVGJmGPvB2+SuI6bxrwmYVDrTfLEnXqdTRf/sFn7LDW/qUULJaQzJRUeEVOQHf3eWB8tJDgN4vt
3Z4qjiMz8NwzyJh17nQkwr+K1fDmB67EuTwHulPvlrHpPsnzFxXf1pgq+VAF4ECEyhwEpiPuMXZN
Fu68sMc1E19qnR4Uve/LPOApmG8BYH4oTpHNTgMsZ0pgcJtprepRVzs92rBtXSlpv0O+tAn7S87G
wqu6ODJaYNaeQjEFELUT4eBlnhjLhOh93FRXelNr/A9nASO1lphBIzHGQ67t7CidDAheLbCMpsz9
A8TKCqgGBwMRFXc2FrCpgguoy+Ho9n6yFmmL/QOX9gl0/dXEcEpvsPKGuDe9o1ftwRhCuaXbJ20H
BGeTvb224ZELcFKksRN4FzITwcFowYWd6vCjIEDxoFauF1xYYpPl47L43Vmcadx/cbu0r24ZPtwo
jw3nlShOg5Dy3FM4dT0gmtLine36rKH/3fhN8KGQNhRLARzZmB4y7j+/zqsjbgVI/SPktWu43mLR
gJ2nsgQtEGEDveQmL5GW9pzoqvSkfmrKrgwZNUUVFHyNtDS/TxK53cW2ut+WxHqKVYIPYUgBSkin
3N/xBjvpMKBeOjYtAUOBrBnpQ86HFzbyu5Dl1uP+wNDN7PWO7nJh1kWGaCVjQko7FQOHztzCjBx0
2jgQV7z99NRmVVYW67Kmcu6AMHaRj6McR3tKyxGkLZKH7yPBNsE1VUe2g2UdYjia/H1kevXEREml
jt/tbDxKJbX7B40c7drcyIL52OGEOMs/x8BPECbx4Y9S++MmDO64tmIf+WqXbVuB46qJqoUl6xnV
vxHnQarw4qFbNdGcoPyPcSs3ITEwxdCeEBk4BTNo5DAaRsKgn6HVwvR2c5oWWUprzBs6mpbmTOH5
TsFPydq0ipyhNyKNZn4HPdHUvdPHLHDCek2ja56RFb4fz5ljvzVnmz0LxuXALYmx+TtldD4HKUR1
oYUJXbb0c7AwH9yQgaEoRk9L2en6hFUTefyT+TK9rWxMlEaYSQ4WiTab38lgq7wjwHaxXntCw1II
yJised2BazPy/6scpxO8DbSHQgDyHbSrMk25f9ZYgTHNADEcPdRJgBaUFN55ZCo5dkcAbu2AYG+S
nEO3SOchyggMOJQAd1upZJqzNWn0BKN/Kb7piCOZDlqNyf6Vz4y1RVNyRHR7/nZEF9RtjMM7L5iL
38PFTXMS+fINkHdWHMR3R7U/m01mvSbMT3y2QEJF2Uf9PTWxl/EvyDkCXYyjrGHuTDXnOMsZZ3kq
kR71eMytpaRuePzXhp5CzJZAhqk2hMH0xVhysh6bifBKkZHmcs5TQDJ6Y6qqYY8/n+Upb1UykABi
idnmY/bkcuFet6WjGUdkwM/FrQ0x4gLJI6QpNQ+UDWjQFigbQBOdycwV6f9jJMy8EWfxN6CuPbQ6
8Fba0uMVGajN3rIk5YGeunTObjm6p3gBGvW2Gxb4ijJzrkZtEuOXLwBCYKBho7ab40xIeu7blYA4
Qj+tv7rsIo5TrKoO/PewznFnX+07R/oQiHEovgzmRvceCiACD2WwWstCR3Hux3h3wSJ1roTNkKW/
mleOhe8p71FUxhjICRhQrHQdy+j0D1Pt+L0pKqoc72aCBX0kEm5yUIryCS9kQMMAJjVedd9+mA1S
J8KyCIuhMJBfQp+T9C59AvWN5LyXlXvCjo/RYbXRHsDTVBUfaCRTRRDlJfhAK4NLhFGhYuTOMLO1
jGTCjJeKKBlm08qFFbO1M3grjID7FCcnRX/fDefjVAIla1aQif5yHcuauXwi4S/cErjbjcs2Vr01
Ri8US/gezH/QTKB+T06CJDg2idiy026YD/TOIBKyErJUyEhhzpOMiNL+GMlCca7LSzJsi0eBQ82H
FZyCTzSFt13MjA15DnNQX/ZrJHT13ussgBQC9s0NLgFw8F3mexS8cOG34hQirs1RC+pzN0IraHXq
qjsbBo00sgkmgmdfIR4Ibv+o0KZD7Br6cxusn7clhAe6gBklRQdJaY8G5oOcRL0MR0k6nf+dnwAY
SFP5Kl9HIXhoMq5+R/6jrJMjChbNx7rhCPlqQkzvoqU9hlDKns9ab+mGFyySPGBeV/evwlhQ96Gy
/wzgTQ8Ey5UhGN1AtSa4ehjH7pM1KQ2EWRb4A7kZsyIZnrkYM6D+AvTyLR0a//WiClni1YCiTz2P
a941cIE9BgTTGUUkdUwmZ96sprztj60pyrd8+zWSFPnR7eCSzo4SJvyuSycPaI1TZaFv/4v6bf3q
dnKX6RHY8OXLrI+ZkjnA+040Obd3qY/FBucnlTVR41TdvBGHvebI0I3m92nIefJG66tDYuw0zMB0
iOlFo6YpVWS6ZMdy3txDDEA/M/+0T1fZ4//Ly/08wOFSLqGF1ruik5EVKN2VNdHp7vbaqwGLApHr
1iNdbDijyoajtbujvm0WO8SeFEaAhFix9XF4NAMwZIyhh51AaXcNg3JErNevcMl8WmCKhQ101sEq
/yzofrZrADhDkYBvra4XG3YuvC4LAhmu+NoBrfcSEmL83mxHUC0BDVjN/F/jYlR5SZzQab+Z64ng
C9ANwO3W+nmeEboAeo1CgKOJvBLPsH2IE0mPUxckIQEkJfMKCsZgWNkWmZwCZ/sPWHJ6HnPgAKgF
X0I7QCNZrp6PDcXkytsrVAJ5VFym6kR+2IW8ot9D0E/yhsFWqhCBEwmp76r0xY1UTI6nPFu4BEZD
OmxAoaKiaXvEi8Gtww2ne/rp77wvFYfO3dSmLrJdJ6fNj7003ZxxFBHVOsJhikYjvXYWE1rueECy
qkYct2cJSJtrrbSZf29VR19pwJGJxFBkLAxxdp1teFBGjGNTUQuWewgQzxSjnq2kbwIHtuUd1bs0
HfK0dyM4ZeAuQifyxo4Ap3VRTUipHsozsoDwFS45jaHdSmgclTQHBMYI4oxJF61NpUNaA9gb8cUT
vYE7IQuZqXVdAcdeeQ6OKTaYhp2BKqaYQCoj8D0W9iO5RUmfOcsgwfk9AaJqhih++7ISgSPfzo5A
DXCbqauX6R1i3m279baMCeyz9gtTv7Ri8om/U2aJo7EW40FaBM3YedBfMCDJFw+MF00D9bddQQbq
h+Rhwtsnj8kosvbEHGjtCPFAxegKb6ML0CFVblDcDgkxGJhbq6aIfGniRhKfRrSMwB1KWgqgMqko
AB1PQD5P24yKfaQBMU6SFHscW19Wh0u3C6ossim9tYe0sTHowo3iVW1t9C3AOwRir3RfMNB43php
QV8Jb0mYmv5FG4y7IPO0Hn+GgWnnKhJQPkEZcEgGRazr6UrsV1WMahmdUh0o3WBoDzQRTEMY6VXf
Wj40UGKW7BBsN4Q/9o462seJ6G4eCCyX7QrUctFwzjlFRxZYDixilHunS5ZGF8qlHV8i2vNJaGzk
cq3HZRhKJIX+OoXRMyIpWAb3bwUQUUWz988uvO4Bs8uP8AePTODHfBPQ7u15eH+jWGzFQGnfDvcb
bYbm7u0Ysukbg5/FZ/bAN33lDjFvrGjQhFFUzdYnvBu4CIro0/hQgE+pznHlUV4QJb0N0PwTGE30
Kj0IpS+e04NyI+s8hSSnFHsAzopoP5YRADRWFr/VD7tGDgI+fqPSe0g1esR/b7pGnqS7lvo0noy4
vCYVR0ndU8EPEc3TmrslVm48yLDDuvn2ypBMT68KkGVzzSfoSSSTRncDBI0eym3juJz932+KbHpc
T0YBpRaQXQriGoQynNXI88zaUaxMVjmZ4OL53amV7Dl4tEIUaRdjQv7yqy3ncZ3usJjmTQOpTvr2
EHsSB7bmr1Fx4i5s96sLrp92rRhcqCq735LeRdVqgtM7q+srGOLznurdvK9M3jylMPq3dgFzppBe
g58n4xNgd07sVFMNG/3seSHkA3Y6RPXH5IqH4KOc/fjSv4j394llSATvObw3qErioRwO0/Ex+ccr
4dUQuDaFpyxY55CFTNKxABEumgSG2U/b21S9qqVeGJqb0ZnSXZuxyGAPtFCAAXW3UdQgG+xJE/dN
I877LzPpufKgwrIGyNYg93a12mY5ualmsJSVE+Ipkc3p8dLgjoVP47lgnC4i/LWawCPCy6TSnYmQ
ber/hq44iWzwmbUzjKtKVolGJ0/itXDSM4HcA1A30BTWJ2N7iMR7ub8MSRXuCFCtb4LtK71WbgVS
FK3MqLtQ3qYGKcXbj0PbBxAyXL4KaQKE/TwREWtze32xphYtAviO3eBpWlWrhiLIGVVcCg+YHjZd
jHcihTW/nqQx4Ixbb5Q22l38YJkqsuWMK6jcl+vQjaynrms2qBGA73Kwqv0B9zbc5jzAoiiB5WT5
bonqnBIZDiLWbF/pfkwayUdJaKWh/9KYi5QOh/N/4rJ+gz8npZ5NIQV7vv+UL1r0h9tzugjy/RLg
vaXnhJdSQg32VV8+exvjWCelRFmSQaJOG+U6bdmWqqvzIsS2+1z13JnIn1VDnGaL5v0P9k6Ms6Cy
JtHrPDhwIr6Hu4edD0JLfcpW7KJNhc6NOdb3VS0Ym2HIziwFiumuukWM6KIOXAVUFmdXqilm7YXh
NZDN116oS3ONGZEFfaYp9931jlJP7u8H5ZYvj+KD/OSfx5rJohX2DOHk1RI3hiD2d8WJVrPQW0Bv
UB8H41l+sPgN/Fg3L3Wkneh14yqw1uyrI1KrCgW2wA5NH+YMgzWrIMNKF0dY421Y21ix+RO9N3Hu
rBxytIXyYu4mUdppVsnLj3HTKchnLnvvSXGHtkDI31Xg/hwV/0JXRNb9EfxQiJB/yl1bnwAPQFey
IdrUIwbDrXAPXjZ92cee93qeYXtjmishAmMum8vNMYs6YUnwOzkIocFx73/nhOA6uSBmsIf3ypct
VtKXqWjdHGwIzL+6Grr603hqj2votignFFydKoMf5GM8+tpehlB/Ky7+EFpt0hVIxfxGZP3Erlbv
BihRhH1VveL1uB6Yb3pAIO1ARtbeV14VGUPAo9487uHsTY/8zOwIfvAPOJ4aHkVkmS/sRaLgQil8
Kef3Uu4SfHkiFN8OB4cbSb5OhvPOnGccA+OsT4HiZCGVvNwKKzms2BGwGXXpPyTM2nuh6sTv/dxV
xS+TdRVYz+Va75txDp2fF/bvzT9KwRdGZZ7UmJED2menBUdBR5FtbRGm31Od1cmWFHPbnWj+qvZW
hJGJgMVYM6MEV/LPSgMFHGMhx0ya3V329a2rNoYPB2J3SBV/a/lLHtKUrZZPpKITB6X43H4zChCs
a0mKu+S3Fp6SCeB1wzaY0w7W0Vj+tZiLoIAYMZT7BzS39uULaNlJaYNMLinM7SKVrE1YdscRjjhc
nnStdlMZUYkTtCKUpQusYeXvz/LsPimYROYsneQxMvgw7qa9dHGoriJ0AYjhfCCw/o1+cb9c7SWf
NPoUzBObZH4tGBIlcEVgMzL7bx8XPzuJUQrM5AwvzNS0Egjx6Hd6s8zq+VHeGksPkkciQyzIGUTm
cYs5/hMYTX+3y4QYBksTL6mwdVwCFart9Zw2Ug5tMAPmhlfYYryqrSA8hM7YHfECvHggga34n8qf
iw6FZ2TV0Do+Z1ZCariMZDfarq/qUZQtBwbY/2VFJkL21ds/lV7kgkJGZt4Hg4EVX+ym1bQ40E83
8XRs0FLkpxocNb3BTgIrp7CjmGZQlkNODONLzBYgns4ku7PG44p9km4PwpjYq+BRZVrhf2CKTVF7
DgHKaIytCrghhEUZVpPaBqd/HsQtu5Oy9INUFZypQmxF2rMHAatregobRUz9/+x3lGARvli0XKTD
lOnS4eAkzeKBaf4FmC4Yh3MYzgfj8kGEivrFN1osaPbfwxIv+Fw344q66ju+pIBV5sdfXJRtHV9Y
KeIX0XZnAMlJLQ3GX8/yL+UTJQUIwe2xZl/SHebav1fnVoqhgg/nGmC1gq/wzrn7J/LFp7D9rVv5
HT3hHVjgLYEXVxPCoGaj7zduqFACMWANOsG/z+SbPNGmcT4oulD1HvkChNqzU9a0wjyaZ9NEYcqU
AMLnzgtkTlDJgTaHEwp9MtxgQrELzXVhWCfwCl3tHKH6m6mK4VT42b/ziwYK+IyUbroKREWjStE1
mTgea+6dVbJTJ03L1nWMRxr9GbzXXwDdyWnzYV5jxonnBO0vpZPrQIprXRDMwIYTp3lY1j/oGHzZ
DrJBkvHZ9Lry3DBnsoFWteM4TPApbO9DYfY1N3MBB82GDLgIy2VgQ57fn/daOq7npD+4B4AB4uIr
MnaNUNT9dE0S9PnFc0ZlHZy07DAbXWUGeZZUQ4OBzCE2VhXw53ma+zcy+ugjxdppguWM+V/+KT2w
BHtxsmNi0OLyldWp4oNiAgiJDTqfjj8SjRhI6oEdV1z8Ipp4MYe3yJarRcVMmH27CJ9BmgISDW+7
0szIG14+vxSkLQ/mKGmClofvDLdM7+mXJThbLmrurf16SixJLERjNsmXiP1tLlGtJV+oLOqTXyoO
iA8ytXTXEyDRuXE0IqNqYPB/QJm1QIz5EYOg84/wxDDChifyTYTmg1Vv8gthZBmOmx1mjX8nwGmc
FJEp9qULx+9iADiKrKRcRjtk5YMLpfg5tQr5b4fGGgcPBJ44QutJC0ULCTREQE5bM4ctOzB0+g70
O0M2ErmnPKCTIymq78+B06Tp2Ai/w3Ylr85Io8TRqcXMPvL7NtSPq6a1Vo0xLfgnV6cnfUflQ4Fi
+0Z1tFabGoEq5rZbUnaALuayk+5fQS5WeUgwei7Itsp0t9npHXX3E1S6sfDE7ef5Dh65wrt16f6e
nZkh6Tdo2Q6IdjvBa/RKlnSm6RDDFhuXIQlzI5l0ocL4fb7FP3gsOokGQkMuEhTWFrqaWfTkVxCn
YzEOcKyDYYTGfizE26oQRz4nSIuKQpNT+64YCeZL9szJHNf4+sB3AB7ZrpNqgxDfkyvJVXq+7Fao
+rjAuQVv4CjZeVN6MuhVhczWPUP3CuN/ST0scXSzctCIQn5Y8ZvaN0qZXMwzl97w+Pu2RLp59ExM
uLPklXhxDVO5pbWpS7BeTsc/sOIwhiOzUZyCwE9dTgL+ONZ951+jkXp038BBw9p4MPsQucjdLXzd
B4bspx3Eh+Se/cMVzyvbdNvHoBVDhWTC9l0Wb75Tgg+dUB5kFpMO/VVK1A81StyBi9Gh295SMAdT
Od1uEazTh3bXsAzooAeh1U3xuSBvDSoxY5DK/CcNVpxnXnwt7Y7jbhzm8CSx9TyAq1zQUzY5AH/4
x12fWO7UNf7rb5+7JtlK03u1BEGEPv/ICOLbNP/ZzdswIJ/obZIoIBtFIb/zK0HMRLGEa7Nc+G6w
V6OMuX7wp2an8WywlXn0jR4dACNwSGJgfR9nb+Egm+AOtlXVJ9csFozwqicMlVY36Ixax/QdCJ0H
v/bu9vkqsf7VYhFJWF8qtGPkdlF0znh08WJMee9FsSLs9uXiEJja+jLcL8uZ4v24bJKN3Xsj61Ww
4NxUoI8hXPlANE8275BDs+OqpOFUNKeH5NEtrx+jsrVpgz19mMpOGcoO7ozfQTkKe5SFMYf/XZN8
lDBTd+W5zoMYdoH7WETAj8Vw/TVev9ikjYl+8dr5OOeqG/reYw5J1JtVz4RjriuRpfXlz39YRpgb
iaTl8v6zGuU3MjyQ8sJ5Lj94WjUEPJF4NixyL2H8uSe7vsUsOo33Yr0JDHPlAvuZOZa2thUBZZgQ
2IhnM4L4pwsXm1PJuGt6X/qHsd47eiiTT0nCcTg+B305VTp3sA6qOYbHn0EfyJMbg6xv563hysuX
uz46JzRobhdw50N5Gtpfbr6nR1h2slO4hdXB028PTndbzQuBWQVWwydjFlZhJ224xboTtvGv84Ul
l5as8N96/0NVprmw4LzQBy5mwKUnDr8V+ajsxUzRRzNhuved+wX0bVW/N2mXPnABUnRGV4NZ/Tjy
Jms5TVl0HHsTKOuxH5oBeNQrgCaoowEDByR5ofmQxXlVWtWw2Gwrh81nb0kg2zDXtJk+fHWd43WG
m69Sdmbd3tPLcKn/GhGz9yo7BocHC1hXNVQZRzj5BCgEk4yuochrfHobe+DmlZ19dC9Evq2r7x+q
gE/dZOkY9iE/hBIbNb7w1ElceE/JzNbfkwDKNvuvD+0LLYUbI0AbzHYZUzvl6evOii9uaR4mUPS1
mb+kQo9yGxGqU+lVs/96hQyUhbQeNke2LRzDiu3jku3BRAgxfCkbGNYdCZYjztyKhfofV+izyU7y
X7wfohAE7ZKY/Wbzneo2fF7uBa23q/fkAgZ56PSyghFsn5tXJiSHDrpBSPdSxqA3Ph46JvOUE+P1
IYvwtZIbxX92t2Bu7vvGOKKDc5sG0OFhKXS6Sx57OEdiy8soEkWa9dbDLYP1+Bv7ZEIriHosBJdZ
XAgtdWrmtLaaZm4dhKmameOqMUEaePlhK6bmLRiIUCasnMXmhX6/kF8kefgzB+7TU/AxFa7q6OKk
k2HpaYQd2YRGAZ0omb0NfJSOrEq1kFZ2gDRUm19sMZCJi9wCS/VWkdeEp9zbNQolVCZvmFseuCGj
qxnnoWzttLI8MQ7kAVr8m0qbULIW6yWjaDF3I6QKImYhktLCXCvcWSMfRI51eInFK5AU+8Se6dqb
0oKWjwKzvITX4DtpOq2n9q8luPv0g7xFIMGyOn6mvkMZF6lXy7UXmxFwrzQ9quUGqdC7hso6axhj
57/W+IH5nDHJZ540ZUovzaTFSpiyYuYgrxO+YuHYQxlAZFEKw0tp0/Kh7ersm36C0cVi1JVmN0uc
s4/UkYZx5qAYQjo09f5ZfS1fZt4fUxQAZzgoEGc1MZLmeX07fV3Ufx9vLur7pWXLpAkHRst8llxM
i/rNypteKChBZfWkPVXIkxndt5TSGOExfPQgB9aChnAAT/E/TGFFiiLSHX/xxnagOtORF+eESd16
CtqHPT3iWA1xLC8iZ0EkJN2NhCTX+BTUcWz27hOq6z0DzutEIV+OuXJ1T/mvNCXvJqJwN/CrcJTW
lsWtKBsbep8NBi3zJzCPF3FSHMd8StXZXWnj80H8XmBbvKteGMs/BHGdcTtIXbD7Yesr6HBmDc2R
CzE2zd3vc6HdWWY+NCuT7PkzVYp95ZP3J40t/arS1iJ3IMz4r/xYY9AOwJVri2fHoDGrlOXcaXbf
OG0lN3QREqp/s49txQymfc10tVQ6MpR7bqaDTzPx1HQM0nUcZQNgFdX8FmJSc6jMrC6/72qMMH4j
FQ4FVHhz6IaKstdU+Hb+F0xUw0E0pu9fXT/6+ZiB3kGjpLDb09d3HHPXKjJDIIwie2Npa0LLrAv0
AMYH2VLlO1D0eJd/muiax+WG4euZtsCpyunEwk+kx3TV+g0ATpMYOFoGvg6Hf90XprgIKvGPoOX8
F06a0bBpReZF8XD2dY2icxwfFY77E4UA1Ik6uvhObLsSg4qGTY0gNenC71jRXteojkjffUQtK7vP
0iVTLoOOhxoR4LXmplWteA1u984UqMRmAbUTyiWE6x++MaEIEXx3rorzVxQf8sFHvXbYIv+b0nOd
hn5WF+VMgDxnNlh7YBnzRt/s/+KtA6lKFZB/MNgj7vIwI7KofoCkngQ0UxbB267f+CElXHhHJ1PY
LSJUITkOkzaZJXHFr3vSXGjEd7ign4H5oK+OwnNlqhNASoUFKKpdob98MUtbvLxwekIV6qV+sirN
9sw+s6SkOYw8aDMx1Q1jeKxER2YO4me4F12MFmuyrDZ7hFtcVp7erIAV7zmo3h1eVg+w6nuCw9Hw
wYv8AyB4biZruHP/EOcV4ji2M7aB6ISKSZO6ndd2JG1U945bHjdE8Qb0ELogzk5qIuO5A9+xcmgZ
HAJ/pYBatdLCHNW9oMdwZhhweIg3nDtG7ADz1oBH2PTWjDeqt1ruMigs8iAs4c+XnkbTtrHV8Acn
HMM9WRnEdOrUsMMMHmK++qXpugYJprb8hzzT+3DVIRzb7micsqGgQYQf56GDpWDBC4mdj9pg+qVR
iFyW/rMQphm6D2WCySfQhRcKc0o7txm4okGVJWVE/zDqbR3+KsdRm4EQ1p0B4F1aJv3ekCB/8Vd/
OXg8Uk7k09FTSwc7Pm3fONSqah4CnFhm7Nnd3XOhQ+3UD8UxqS+jtSVPWD12EK1IwYj7fNvY8VHz
zS0uSrk7NDo9WnM2+TuKlABkCjIiVpTsCuUEbvujSjwv8SGwBqNeernpPGxcdOXeFRR7ud88pwnS
idkryltZGdX+biFIz/WLEL2L4j2pdxe9qqxHYW1iTKW0AvlE8YxxoGtuIJ8AQ6NC69slD9EQjvov
ormVkLgNGjocDfZotG4Cy9BC3QDwMzOvIuKCnTQ6YVYvmuhy0X8biVLu1oiMGNLQCf77w6ONr2e/
xttwmrskQTPez3k1xv64Pb/rPhuu+YiSh5zvXkB6iRd5B6nXiMzGl+ZYjbDMqpT9k0kBv0Cj4xbR
pfPEzVV4MASsIMgnrn8ovUh7hn7A5ifPcjnmvo4iydcn6ZG1zlAqlqH5SHcIV36l2MkIUoBnOuLc
EPxULL5TNF/u1x5aTidmWytURhM3XLvwhGCbvRKCRCDEiTD2pcm39yo/sQ3vSiJgUacbvf2Y6vlA
U3yRADoWUYhsTLIgOE9HuLACAp7oFGw85hrlqVbQIC0f+3ZfFniBIcvJ0BO9gyans0/RJ6aLC8xW
UnHvc0+kfgOwX1kEtR0esaeOT/ST9IYP5W8cNc2awyomTa1Ji1Fetr2fURmEsyUuUZ+cSFAgRft0
M+qKjRKJr5yy7KSvSsY75MTmGmac05AWtDsJIdBL4S4VCppQmlLKSWLq17M9oQytmf6X8pyZuUG5
ZX2o6jsAqDY43IVQ81O6nxKVFUqL5r5SQfLAngsBbE7+qHaXPngpzq+wcfNjRPQdJH4PnLfHBCii
bK1lrb/sey9vbMNtzvwNhoouRTNcAjGF69GB1pUnFy8deHvkPGLo6zSyAc7eO2nFDxSPVtv8i4E1
3ReY62DTgHB1QEEm0u5SjZDE1qMt/3lIx9lK30O1tKGmFmTXiz2OJew6kau7UYilfJ9x/kZEOOyl
B6dQmad201dZIk3zN+MKPOKTwj/OMHyJNNMx9RqhOveD8C//tLTzOGy4KOrhkSaudaUjs02vEOGh
nFS3qISB4dGoPZj4ZpL68R/4QtGx0oDfAlNZr1jBycEr4nxHWQs7tZ9FYAKhxHvgdou1F+BQ2I60
LTaWzT9lpg1U3MUIIjA5s2qgK81hQgpsqC4gSEUp80ePZrTVNpD1AB33YGGApoQDSyG2GHDdtBPH
SWUD+ptLbVzyd/4xlCqFM1nBu+w32ufu6oQKHp0h0/U3GEcjKeT+7ofPNWWRI3mbHYUsQP++zW1q
1VyixWiURXAej8qR2UWaYp2vWcSb83wlryZ6JkFnegCMTtdHQHkgiFHGUoKaz0eYvkEX+MuFk5Tc
bNwaz9dDCioC3Jqn/Ev1rdi7L5I1e5xPQp1fCSgpCmdm/kTpf5L+S6PCQifJ8CcNIo5CAr4Jkj4e
+FnM+UZsU2KqtJvWabzBui8BzUf+otxKSb3ZuuEX8CUWanFOJYicm8T4xaKSYdv34HQ45h9mPKtt
TDGIrJM1vpkT4Oi0vSVzuVRcf85dDjkA6Vn79A00JikBIy8VDldrRLEzc1S2cq00wVMKhXNmLmLM
0IjUjfyzLpC7QdaTQUbl6XNdE5TNO4XrkoUCe6dKKWwbdYugWiqkn2Q9yIGpmNk0brdK7VUBwiuF
O3Mok+YgOgV3l8nInzgfFDDoPv/b0Wpc03LFqVerv4c0sAwSA3YRmgAqYSvdZp7I8gbCff7lilIf
qW7+Z5vXRViO2e+LDxZ1qk8fETn3yt5JOA8UEv+zLs3Z92Pm0xsKZlQcVq8/PSy5IdqMSpLWKRwO
7dumzAd67L+XZC9vUcOEgIDXoU7WrLEi5kKIoykS9OMpnjn8az3OsejWscTWDuCTUUQy8WFuDgnX
DUViycF0hED6VaV2Off9iCr21ldo5t9hhyfPBhzNO42u0B5zrkoFk1jxY8e0oW1VSqYGX17jrdYh
s5NM1XRDNpezLvo4NXi1Z6zfm1OJrwuMVUvfvdt060ISH38JuUMIaW73LwnY8nvptrKO8qGK2Jny
kqq5ezU0vwI+MXDcdegincjdTDO34eMgU8r3zFWObrhQ3IA78C9ESKD7zuvoCyqCxpLsPRO5BNbK
2CgeRKWkIorVdFoprzWq4m1wDERmKlw3w4o4VqEWBi4+7HCARtfurCB2o5OYwu8Wz3uDj99jDbnH
5bEWALSmN6WapyTQFzuGucVY+MQf3alceeRVOaVnp9WKHoykcZrcuaQlwBmgdpGPX/jHDGhI+YQK
xdhnuJmGvxIagJ9fgXcE+7IBxdKgUSVoncg9FUlKRPHkX4qFjy35iq44UkiqqXsmvB/qjqSlQpEu
NHVlTJiqlFohTVmkiJkqeRbDsIOJtZ1/wOsL4LInKwjXV4n3IVkVY02qqLcRryBvXaFaYV/6YKz7
Oo6QlZX68n6Oa6OC4vGlsDGDqnpI6Jj7xRCYkNEAd89n2ULvaitSprjgyVNTqo/bRj6tjN0kQLOH
SkRbAAbjSu8SekA7/7ff/02oSeeus9MmSxD+5C/07YNzEnU+LkN332YEHhOhusnXWrXwMESJVMsr
kkc2HdJDLiTWMsYkQI6r0f1IoTqS58R3opr2b0tmkNWovmmGiY3eJynkeOxon8Hpmvy0ykrVJPPi
HGUfaOK37iVQ4NuahRkpePhEgcsXt4IZL+Z2aeZtsczAbWKbNjqtvtWUExtrIf46cydbm3MWxeyC
TpbUdyoOPSNsghgILW665s/JGS1h1JjKmPm85yDxQG5CuJl8jlrbooe8cNDG9QdGAQ5vJ08VazAg
mcm90BkE2BpbQXUA36PC/bBUrpsaTrulT3G+vXI3Srxge0iUC/6F3DJ6JHa5SRXjOXRzQ9vmQQ2W
ePV+fc/ubuaNsIAznGUgDzK4XlCX0SzZQNc0kgs+iQAIAO6OmZFJeIJjChrDimx+MYdDtYE2B2j/
oueYKmTb/YQBhDDACQFECtfiVVqZMUIWBH7BTC+2trVueGNlDn1wFhkmTJ6dc8824xTRvbMCdvlx
Z/AenKb+8H5bwTUwSc8b0EGtNN1YK6q9z9N5zj3W/EMDMX5TqZSWVQTCJ8/FAdHC1C7bRXh5fzx1
vaplcb5E6+503licjjFVIt/BTwJTj1c9IT9Q8+MHkOoBKkWsznIowL/mhkIqXW58MZt6SheAm/+Z
m9RIL7wSVoxSOFOu15yH7sN57nuaTeJGgwmCcg46W4AoHsbcRwILKH0A23k0bSIwDrOCuVyUZ0sg
QQ6evtIexMxpPKHPCJfos4G+xs4XIpRT/15R+WLB2O1CKkDa25kRtiBbmf5q8fQgqZ+kpcV1RC8y
vsXkhicdjw7vfHR+xcx7yYkp9QpizVtqHjkOxH6jjOF84dFkqO0qZHeTexxjUcc47eSuAt+Ixc1j
Tlr/lzeAM3paYcNzNOaY/+Q9DyMtgDa11uGonKnnONcc42AlcpWgxiw23/pPHILcQKp9QLLArb/v
xvecIon6zd6oehBq2aR+pkMPqEwercK5HQCjOiZQMNH3+/Ua9+33sqyK/8JOVhGDM3mLTFjlorO2
UqvncAUHIzsFQqkcLMc1ihSnbORggKn4LqdzCXdWQHFc31do9a6OUEnNWZUkW7MqfAnPWKmO78gv
FVnv0PCASgYVZqwpIvORAkSOxeZavM8CWsTWh2L4cxhavNJ7e5/RNV2ctLUoTBTy6SW5J+VIcVPO
ceCv8uhunU5RHGsOxWmOpR5HQVPINsTBBsfPqos9D0QA5jwbvoJSp19GIRuUQboo3HynFl3Ohyue
9+NMNHLaV7RyXAbZsM6/gADS+FoVfdRTMVEDQF69lz8NYtkLxG9/mvHpVTQxxs1AkohwM7+Vkbgy
AMqC3ugT0pTr9LlqQuWxQHJcaJskaxflz810QHcbISQCQAm94eyfw3hXsJkY2u9+pcaS04SrwLW1
jC3ZDoXfuXaoCdBw6x6dIG5t3TDBxtiOH74GYvS/8WSaef5N7Ty+g9pDM7Jkz/woRk0tl2lnOMbu
mngPEmEVnhbdOzNlHSM3UZOFfxxgCqXtLqo007AkkFYtiohYgHYG/uurR91EuXqJeTTj85YP5SNS
/SrmInUFDzTiOMAzll8G9bQqDAFSeckMqSafAHkhyHhHpizZTCfqoAYQPDteZulIQUjNJxYv/bxs
SpCu0k6WbCsGsBGeeY8bfc1TqGbFkbU0SquU+L2h7eCMOyjijEeZn9wJImbJn2a+oHY+zDe+h7ja
JelY3K70kF7kMzgUBRHgWF55IDeRpJ3Uv7f0RZuUmfXdHlnMnwxs6syMedCQ6IUzC8sPel7+3Ys6
W//CETz5zPjV7kiIUfmd4Qz+liWKm7prLqyMgOZR0zF9pOJWwTlzXUIy+TngF9GKMyiS38SGRoH+
1j+mZccqm3JqLFvJaukLNVGWQvxL+LV63R2l9bdLLXldIWODzgUcf9YoRhyy7rATvB0S/maUrPnO
1cg9OVwne8/++NBRRsTDUyqKwQlYQIaipUzgi3gGZ7KOsVAETILzKO3eKWyzhKsQecMAmVFllKzJ
la19iBV/c2mLM9JA3AIFajaRkL+LAkYlte+pLU0+CGzzdmpNQE+2RoFBBvjxU943mVAQG+89rhfj
LBoMZwmf2QClQKFe0bDqt17z6vH9YLbOW2cn4DfOx1drSPD1aJJvlNhX5OP8FTgRaSsL4qtYXUbr
2D/flAwB+eYb55dQwy2HFymvAVQPq9PmfyQ+r3jJ3YHHUXCSk34/GMXtRxUX2xol9AzvYAR4kHX+
maDbP9kYEotJE2X2uOQq+l14KDBseYKATUIVTxV/+xLaQ7IhqQu0NyMmgMGtD/RD1tdp/u1hioZk
Mc0g5ARXYV6xxrSK7qcdwA/rLWNbqSxXQxxfxF0LfXKixZ44LZqsbEyoHTx5BJv+cwdmHfyQs/ce
2js53yXx2cn2VvRjxyQ9J+RhAk/eXLJ7Xl1CkcZLNmuY4pv9RcIUTCiiEv5ejawkFgkqKAzfmDsW
rH/uQIuErJCuYTDEbVA1k+WkGnKIxzZ6cfnrsGYPoM1bwOxhJN78O7zdyqCLgHxWj4yvxBNpVAGB
0MHoD6agvp+eL2VGOZk6vJJU/Z9WX31kxxe6RFP001N7vpKE2zOkHpm5TYGC+riRj+JzncBL9gz1
zi+i2Mb/y4xUYUA/pHxuzslvbfQlA/aZywdbPTzIHbW3ysM0gtAJfO17weyZC9jaa+cgsUIFHEIS
hoMHW7NTnN9Q+20cMwI7/KdIvk0Adb5q6mUif8872IltRVebjolrtfWO+aNWQfkd1j2duzJALNLm
8AZISD//LXg2P7P8Z+h+AtBt5D7bGrT88L+zrZGYmrWudzI8xKiQYiq+dGTcacQ7ro8mR7/FToCn
yqxzzxY40Cs0SwZDwV91xsa58Yr3ic48ru4EiubohKlWa+jclpnVdzCJX5kb3jyA/3xoe5+RVhgS
b1c0pvMsIfrdRyFZ9I4eQ3JjYBOhPOd5N/LRKUc4/lkMRylANIdzJjH3z7pWLZWBjsc2i6bRW84H
WQtUoAeuN7BaYW5R7CH3XeLQR1Q4cP8/NmFZp45LwlzlYTCPmoj0/candM+pYKnpiw54q83TUNPW
DHqWX8LQQpLicACGEnVPU4GwPe/cF6cPoqkn4WW6GWDhLYyisqXHqOAfWo5xFa512Ky0zdPTrGtJ
AbD5Go4R4PXpl6m2OqPwNwLHXT7IGaofPlZWCpQLHWcr/rBvdTu9jBF1NbOOF9Vh5x81ukackl9V
BdPThI8LjzPWTan8qM6VpYKlJ6XN9RxHkhbZTkHlBjStxY9nZhKd3Qe6ADg5RQkPW83xNjCderwH
pgyLK7z9yNglGuVCdgndN/YZIOOd+/44vwb/id2j1Gm7hZTpz+wZpGYB9RgDXKRxuPYsdZjQhwoE
1jLYifVEEHIG6eBfOQC93nt9D6onYQCRJYpr9TyFO2rpuQywrxsT529Jel+Vgy5psaZ6RGpCpp5c
CTp4tcHDczlpfGFMIrNaPMPmDn7NCn3uFeYEqycL2wmTBe5vWIv+DFcHSPmZGezLBPq6f4f2bNCZ
N0wGKFIqW3jGR7tezmkBAIm/rQAtTfNgTjLLJzoNl4mRqYvzvPqE2+4sp1PbrgMT6rLlS642yS1k
Y9Fta6ucDpVAAPjRw8IMDxSk8KhmnT/mAjp/mV2dKnAB+d9sGI+gkFLne0C9yx1Qzfjyftu4y0EN
Potg699fHRMNMcSBPs9weA8xxg0NA6i9DxXwYokjkF8AF/jcwPmtTjH2cHybhmfZcEgV1kkLuumX
di6VYrkA2U8mqIIDpMZgdTP78QPK8Z0leoj8aijFjjwpfgun02I70kNBwGNc48ulSyRuw0YxfR15
9DglSgl1WFbdqhYf/2WZRccvz974Ka0KTfbz04IA1pGbpI+mQZjvirJUINT7xvquK7VW2k1LQEu6
KWGztpnhowwQIiSHK67lan9HAd7rzt/33rKsghdmISGAMhQNjksMHeSo3VAt5MeYopZBw7ukaApK
WOwl/IC0CQVLMOqPVwOJbLC5RFeiGnOZpKvM0WMMoCjRjsT6+7UwHvlKfpWPn+Cg/8ZNXN4G9xFN
Rj77Czw00zV9NxRq3Q9bxHGJwl3Aub0zo/hfTDaAp4RR+LcmmD6H5dWFui5BvZvhWY225icvi4BH
KaYCZbP9sWFfcQ6D1hqX6yd0BchfYV38gcUIzJdeak58/j4xt8Zud0kZwsUANaJr9jI5Ia4H9pMd
S5pFJKRAnJ4P1ga/Ci4F2D0d8zGSrDVyG1aasK15TbSmgB6TXwUuSzM3r4J9SNhF+eQDS3uwynWZ
fuUJrxKaHeKJ88Dr2/RvpfCbio+8Yhdg84kQbe8DqdjqWTXUMJGyjndFHmF7ze167OgWv1yaIigK
cF2kTWnLejfT9jJ39UdY3nmzxoANL5QriVSUAWuhJeUTmpDY2CwJjisWzGjOi2a+4zS1xB2C93sg
P19eAo2rW2QOAKpb77Bkh8ArMk1vrpkwqS9Ma7g9eCLHiFCaIFb+wk+heQt+dPlUc1zcrxz7cUT4
SZXMNVC01eVTmP7dt7tCygXAoIRtDrsPeA4b8wkJ58VPT1/R4gtrn151Pv7XtiGo9nYRj/xV1gSz
IMevB+OLXyd7/ERiz68bhbmnKFpWE6pYD1xnRM/O5aqDRhUoBpDnzPqiCCmEa7yhM3f4+pVMH7hO
gof5ryNPmlGDg72H0FjlzK2zbCmvH+l/MwYYSxxA+f1YOrA3mZyXuyHKorlx0IdPa3y0zfreH6e3
3eSqx2l+qggr4i/7UgEIw5O8qExdqArDmTc29xk9M9anNZ4fQB8dX62OVUT0RaL9pKwvA3Q4MGmV
iBz0pzNvrwA5UipTotdvqQhX5wYIQz3JiyG7xhjrTGnmBoBijyartn3EtlsIgz4Ihp6aw2Zdf0Cz
C79bnDzsjzkt/eyG2b4Bd3MFqISpOcActKAOVSQN4Z0ozQfOeLSlU8iy4e9zcZCF5KkYwAhEeUH2
T6XShCE2ygVGw5aZ87fKDgXvcj5Zjov/nkyAmK3lBi+SnvqqdHBreA928EuPqvNhvjRmro5TlrK/
ihXWI99OZTeg0wco1Dt706+fbJzZdBCJAM7NDVX/cg+NiY8saReWvr6CA9LZrkQhT8LgJilYzYCI
3ikminjvBCCvS6qJEE8n+2bfKXHDVNTYxklr4wuOp1wpm30MrL49rVlaIGnTrQiKqBEPuequjZHz
TGaHLyFgmEcBxonRu2M3n8SxhcRWYO56iS2sBUYNNz/MdUzM8FzNV4cTCrg5lKnf02aDfpoImd8y
lHEZVuthBTF7bPdxISTzQbw7mrj9ow9bWwmXo6jYQ6ilKI+5w3oU+oe1DE0pw61Q4z11uOgkPJXC
45gFNdBumxFRGsgo1c05Vb0FBUwGS9bo+G6zr4Vzto9sry2G7a+C/h2bloCjPiginsLaoAR3B70C
89R9MJg1NDh1vGwwhfXwsbtoNDiANx1L8zEJxYDkdliNMA7zpbV1wwbBrkHfUcjLMBIRo24D0hbb
E2pbR0PUFlb/NHq4P3YK+AjGGZGUYObv0LKmoE04r0uMVyOlpmxMKUw3FjbDJRPQLxiZtHSAsag9
0lsxZTde0g+JnvacCAIaulxulCUThEUd6JmXUGPBrU/JOYfWifcjw7kOkR0+9zqWoNbm5hMeZdCm
N4pRdI4cZpw//Dp0bz9vNKS/QWWGfnXLIZtPrC7uwE2uiH67wh7bdnUsgVaoJp7QSm6RRGenvg3y
VWLbJrI6Acz4IR0fss4Y0S8GdKRRbHNYMS+a5zb/Y5JV/COW5G6Y7pVxTcWFsA6hrYgHzh/MiFkV
a0mhe16ONNPvGljiITquvp1YPwHXKFGWUvDl5xjL7qob8cHRSGAVjwxQVPoz8vPOZkYHDxT+EeNz
wZZvGnR6QaarJ8i6rs/cCWkA9o+D0hbcSi3A3wbHi83J0+eiWmr/CXgNFIhdvt4vnWISes3cfYdt
yu+JQ0Hyw+kgDi6v/m3XEDvrXBViWDu1mSsnMkseSST6OOkjtHSE95Bmv9senfffQjxPtJs+4MPC
sroo/+Km9gVVbwUOobjKfzeG+5dgEHUpCVHnAJT4xp74UMr3MQz9ICuY3o6pkUo+xtmJOispdXEd
cdx21B/QbYe/OPZ4xIYY36r78nyop/yfuZLOPxp5Pqw55IvSuBXlxcaG+uC46YK34znWlz3XVffh
9HSvsKN/HaPucbu3tEYSgp97ClcrtotqBwFUJVxBLzo5+m7on5o+8cVOgh0w5iwJVtycjpiKRTXc
cbizWHMPaciOrwZ/sRAK7D+Ai2XjlA8NUBfvsK1fh2R+K2mB7VDQumhjj2F0bY321QzUF8FJhgA4
f98b3wuGsRTergnDcWmX1Z4n6SzvgF8mCvF08CqjItEo9Cz6vNKb2LdrnEMeaCz5KPQq93nYPSJe
OQ6lhsmOO2KJS02Os59ytEug5UkDF+49eK41kTwLam35B1W72D/E7DWmetXqzIqbeBJ253qiODl1
h5zYL1K5rnxs1WYYrRXFZeQcjLzzZTDVCC/TprjE0AP/g+VZr2cYkVHPbIEd/ef1QfG1QaL7LGEE
0pMIDpSXcWsvmW847965V/ta3umF6fQ++N6UG693LvJ3fveQ77wE1aTcaWOgeKLuFhxhRUc+efDv
n69GDyT4js8n/ppSIulZmESAHX2MsLVieU/RQZyJT4D77wi9PE4+pxvF51uPtw7KhzBu+GHfiVUC
pBl5BUEPXZyJ24odOgSFHtagOgHFFePlQWGLYOMxlTtEByRo5prCAK+CWnwA9WLAK7Bwc4/Ib5w8
kYxpK8u+wE8jq1E2xOv6qSjZp8GBF8Gb5fhVZaY6aBbdXHPTlk4/9rpTfSmdalP4bKdymCAWhUNc
D4t/pTNq7p9vzFv8VK1YQ35IG6WenL6X1w5X84wXaQAGjEUYEBf3VUsGBD8/gY+OhmIrpgqCTz42
yMovKBn/IzK3wUslpr2mpLqBYmcXQeCg6aKMDYnt6/a77fjYm1ZVabAIp/MdnCF33ci03i8piZAa
AOwiI4K8kNJLbKFEF7WqeElv1wvdSiKRfS+EnHG+lErDsP2rhvhrpAZe893izmY1LwMTYKNi18rN
O1TL45KjMcagrCPoG4BZMtylgv2wcH7HZq/q3bmj7wrec5x2Roj71nNBpAPG2q/SN8bUqB2x9ofw
8bpMkv0ARV2A/wz2LZo1x81N91DrXHQCCAhiH79l/Id6Mi6PF5sIdiaixq41//bKbYxBt9cm623x
9Ejei2VjPq9lsZ/nWWDQ9Yo4RXqqv75s5m6MdEU6bfg7wavjsH0m0ovnNIFSrVlKfEq/xx0Mzi6y
ErMvNQ7wtEJi/SuXWcg4qyolcAPyLcPqWoZ4fvhamOBN2Nr6P/U10mO/E2yQWN4BFpvt6ZyvU1I3
SnpiZygYUTEKDPMrc+G/MpYIrxEjOkHu/trQMm/0Pw6v4bNANQkLpeh6869Y7HAK2vDQwAYW1TOC
Qn9VsgByKWj4IVWXvnvAU6U9CRGy7n9IToMuZQY11KezULkr44O6WUcPfBi/7wSYFMBAlxo023/k
0sKM5OrO4rrVlH46qxWT/9gzZ3EitOCGsmnNyJcKCHPO/NG8HJ0zXdJa1fqLxYsnfec8FYdsDwvE
gPWHdTFAleE1tBAJhNAASESABb7NjfLimvE2fhpGmqkZ9ops//ZH3QtWl0X9aV3h/Zyfv7WX+Jdg
qZwedcNgPMEw4STgQX5pXnCokEvyNeIESQBq62YwzNdaGFijKOSSewx2/uK0x3QJfajMk091fjKZ
ofMEudpw63wb6cRdy/B73Nli/hvoz1WakWN4E8MSAfztWHFWEqhuVFZEp2SY9eFmfP2Nq0STevus
pE0v2G6p1X6AoyyUsDLPace3ERPd8jO2UTUNRqJlZiHiu7LaLw1rQQlQt2Wckm3JGkiZnV7wxvkX
s6K5CKKDknchOYy32+Yk02w8I/YJ1FU+g/W9GXkCUY/wnMTCKYjsMDZygke8MbWbrlAtbWtmSxvG
Px1GlXvw+aNSV2UIkalT+11hu7wqmT2PrH49YALrBtyrFQForUkLc9/ftZz7/H8toxaijgjwWQw4
jSyEbeNRPeyv2hNwXXZGuu8SAYvQteAdIkdYBDJZMcCilZbR8OAC2h8+bj3JEyIRWv7ED5rfEgGl
KKFM6CvMfvIawx5bSnv9mWpHNcXz7E8J0gj8J1Jbg3BXXCnbc/14uGQ/JUUIRLJZLiR2kDzNAE9s
CIaCfH5d7oEzhVH/3/SERT3/yHtrh8fcc5Xzi/oEeVGNkzQM4EbJM5eAwHh7l/G7HRXZo4EJm9Tv
LcuhSkaUXEEwIfMO7eLO5PpL7JJbIIIDtAs1yrm7qcp8lNxdELAqg0VJjpzMuAVEjTjJCqqEm8NV
RBOPdf6ygkYbrHoZKj3kTxeocpeSjfxiHIY3OqLyhniW19P5qVfx76SY8UY0bketb4PrG//6GPTl
k69sY5vLHjmZg7inMOszW0OISw9i22AuJJBPz8a3SXOlrkMg5ZiOtnFj43j6Tr9lXpkshMVYOBCk
F/dWi+bDTZLbF+zSuHrjbIEI7XhBPlAfS/E3yg1ty3E8F5P0JuZmE6uP8WnGL0nvR4tMUEEZqEM6
EtztV/ePLVQIMLuFFKZoQb+Brl5/ksEe2KmtFumdo6TIDT8SIRfrbyjqMiCHZ6ltJxm3rNAOSEdM
Np7l/Y1BXzjtoeq0inFVhjqfnyjyqNKIuSYEICGBcvCGwFOy8RSD2yp5U6d33GZbKR9EHNf+c6Fg
LK4LO6FYNk2pSV0v0T3HKPXuvrZ7VArIpSiypwsBuw1xtShx+kbwHyRPyE2Hfeg/c/8nCvmQmXYQ
xHlSt0Ok9mKS5ia8EjCVbVQZYHh3D+pIO2yMRJZJxATTXY1YkfM9XlNh+Sw3kdRlogOz4Xfl9W0X
oDAfHvLYW+zBcgU81OWMFS+kdNLnkaY+xO8VYwp8CzmM6bCQH0cJyYc3C2+c66MHQnXOwQSc1Aey
y77qRVVg4Fwkoaejw654AU9IlOGNeWeih22OyZBudjhIiS8JkI4+F1uKR41iSL2p7w//e74riTIx
V8X2KjxdGy8sEk3PD9CsvrvUfM/6DWlEGvYKSFviqO5iDhce5DgKdxbglWzkHk02qGnP4pGnO4t5
qNEFjek4o7oqgZ7cg58optKbLoMv6+t9hMpJwhcseCIcnYxjFucoyYvFRN/QZpM4Fl4J8i0dczya
yDDKDFmzYKaOfMPzRPDxBEoyU21CR+aLTLkMqmGOIE9q0AfQFLNmmXEYkEcrL0JP2deHpsaS65fz
Wv8I7zHhxcZoL6qF2V4bu6tDe/ROwTTqCA8PnlWJW3A+Nsp8JJjYDPe+DA2A2eTNUZXCDRfDsUkn
wzn80MgMOhKbjbJ51sZEuLf9jLvk0LwiLkA9huP614befJ2E72uOo13ENQFp87bcm23WOE8SB8O5
pKJtREw2U3EDM3mjCKNBJHQ3mbAqO0lV858GxwtfifEcY5saPMxK6OTVB3OH+mCVN/M/vwU40/5p
Fmg/nAfv32YX+vQK2hQYZa0p28OsfuUuXFFdahFH/c2r6C1iiU1SO675AHtBlyKPKKkdzakRW3Xw
Ws4P0vhwoJJY3Uk2dcLedtwCfJazNOexToGA9gvBX5V7mZnmMg1mMM4WKs4sK2BUO0/BqguS3LJq
3Ai1/Kt649pKbtkSOwwgfvMT62GIN+NH3pak1OlV2tG2MVRz2CYFgq5IQc/LE8qTvU8TgKqf6hsl
juhHqhFRxQC5Qntc6SxX4l9lUvYLWq5ly+K5AJygC2RBpQztalDQRp7EgM9KeZxbULRkLabSSSrh
m/Dh1qcc6klqDKmLp1TJ8UQvaXIYtGikvBq5nVYo5zGt6K6aTrgpjwuFsHAo4/zye9bf3nj2jqcj
3cjISSpL1tcuLAi/nxI4uKQYZqacFkzasmficeMBC5CyhK7zfUOAsWhyhaPo4ZAegXP1/luawdgL
x8kxPGs7Rx0X1vU5I2HgMlDtVToWx3wvIY1i3tz0yJwJ/fhnePQ9+P0o9WBF17RKoUU6cIvuf9ph
spMDlYBM+OfwUdR1DVBmQjok4WzqVRsDOLd0WUeg3kqzfm7MBOQYHzbT5rLAVMLOMPHDAg/wfkLz
O7NJI7zDj2gSvK/r9u1T/4WQwFZVdFiHkW0lJ1WC8t294sTDGF39ueMUDLByBulxJoG/lUcJYzF5
PQaTJJbQKnGKylM/25I+0hOWUdQOrtWP5TfBpBLO/Sxs7a6KzYbelUVVpu7XQFkZ3KSr0qm9QINY
IkET47GBVZXqsiSDquozJXmp63W9cfEwYXae2M54SNU0h4Cb8E/TQTnfn4dvFxHCv+JfUVeL6RVE
VKYZwGTjNZIGRcQJDSXqgzHQgsly5w53fvzRh5YL9MvqBiYx6iA4XNXbG/01LAJx9QvEsHibPLjq
jPKepsCd9xxYAsakO9xkVxVhW+XusU+OyDDZM8LsBJeT1mGkWCWHhzPCLP3oIVZi7b5ISr9uNKI0
ztYikrRIi+CRF8Ydwyo2CqgK1/7z/6enbkwO5EkHgWWPoVGkatvQKTxt1m2ZESHuKYpkgrAf7cQ+
ebQSW55nJHkQTueH1eGyEPlOac7pfEvS1iUl9oBW0z1S6MeUjMivxBrpcL504QUDAdhujSda1Lx6
08xLT+tz0lzs5pvRBKmmg6XcmjohROZxRcGQsTe4O/iRp9d3MO2OMthaKiq1OlTON7eAs4xpk3Qz
Gco4PHu+LxuyH+BNEK3Wd+M5u/DA3vnxqQnJxAd0nBrjDtOey1wKUAqBQiglSXkq5gSI2E96TUMy
lYPvLMm2LkoWSvCFFHROXwpEEYPD/E1WdrAcwFMEWcHFFN1UROFJwoIXFZ1A+BTZRnZVHaDrkJ7w
HLlD9CUvJM/4xuQo5qAGBdzeGK3bGxgAzzQqu+JpGFUTHLX3hSnGrIFxopzeKRRd2c8GguNs2rYi
H6ayYPZYZubjQlPaTLrMG+t+F9ZY2d6phNN31g9dBxEdeM6JJb8TLYQ0sNFzqi3ILlIMrzETdhtD
kQmrQHnQAHDJ/+EyEF2OjEA4xvcqgDw2RdPR4CMEdq9efjxAcXJIi6UvXdTM9URZFWn9Vm0BW34d
Fmf8WVsruR8645dcpbduPvVhMcg2jWGxhwZ0MAOWxaFXgSbm2kokN03J5vI0uCpSvg2x69WXH7tH
nkBMdZBX4EuPKlfSaxl1hiph42zQmD+31aQAaU6vIu5NvsmaeQzSVikKpcJhvo7ttZGVHOzRWhgV
w/Lp84TEl1ypz0D8lcFTYQqkhNlIEMn5phWRzGMb1VWh/TKdQNF3JyyUQ9mAb/xjWioZ+eP+mc+V
4euyOp/+W9VagGMbHgU9m5LwiNlhyY2OYR0IW5ye75QfrixyHIZBVemyA26mKdy2FFYa4LLdgvsl
Gqmu4zEZIqBuyifS7lPYGBAitJiKsPJVZg9JuvvbLXwwQ6ha/iz/a8EjBhV36nfNmr/JmG94qGNc
dPY7XIRpWoj0SW1nkJENXtuW+92OdP3jvGgaXb09cjElmfGnXwza7oXiKmhTOdR9OWtGLDF7p/Tj
EhgM8vkHwqnYnHlGZziZUB+XOptU8v8JMzI242DT2uRck+Tjky/Pt85O5RF1QZAO7KqvRTXwLE3F
BlsCslrIOBzM3wj2p9B6lFKTtQV2X5pqGFKfOZ6PRDvyYt4LoYa9d2whXqpUHj/xR881HiOR+LZw
Em2hJehl0YWyukxxr5MNwEuCUIaB4JLn3wou90MetdGRSMl3QFR+W8Y14Rdevp9qjbaJ6L/UHDVy
ZbEeCpBoc38sGjg7bARyAp5YxhpL1HLgGA4y8oDDLZAZzTvVmFmNe4lkJGAnxdEAZ1ZkGhqdERVk
01BRAJpscfMzC/xhIEC5nUavstwgtvVXseBJKfW0xLQ3GPzSBxC1TZ29noz2NYNkD61eh81Y3NTy
T7hH3KTgLAe5o9QGTbhN6kcgF1fFqgibZaecMN1iQeGAHqNUrQvi3Mc2vVABe/YWo06oJLp/PDKM
IC1JVF2o6fUht5u1CO8qPIrk1VeEBQH8uJ8WORVWmQaDbEq7kYD+sOi7Le1LC+4AcNaVnM546CWu
XtIsEWkB8fQbNC0cGBXxK14rEduvwp8sto8ESoZ81d/i8dz7hIwazeZeQITOajNEgrL3K1i3ZdH/
O+NDlr5cLWUk8qXKD9xhDcnmSBeov5vCFHBpuGLke6WbXdmmB/6HClOHLn4Usnja0T2izfW+BxYp
oMSp+x3cfvL26qXiSNbNTI44tftRSNkxl2aoSY0TkKPmGfxI/d5wUHAli8sY7JLzY0fLBEQqXANV
lGKRaIt52wbFt8SZ2IWuvuDRxxdljBrAU+TG5QEPu6iDsbPWM9UiFpVuzLgMpK8KrdVli0dDSefL
LVVtmg9tfMeVIhm/gdt1YySruLzsRBctiDcMhUhTEgY7EY2+aaRKSyuncMbCi+Hh/ulBkuhNtseS
YJtBDU8TdkddNU8Y/6p81IFya1rKFdzzQTNd+c4x5dFmWGt8uv0Zp+jxjZN7lUtN14ZlQPRY9d2y
mV6ERFKZrR/RFhat6Pz72bXlMOMpG55U/gS4nPt27y0U7wj5VrZzt/XAKoIdecbi2kNb7RutocA3
Q/bz2FYPsZPbJdmERLkUnwS/FJXVpLscYFQKprHvAwH+542OvbsB7mSIT1PyeWXWiVvJtiW/Ph4M
6UamSPjsLl2RlDWSJcBoa9SbpDF+lDoQasXILOdl26OqUbnBpzEQ70TUwLt2hWbGteOvMZ2Gxacp
tZfd0y9AXpv7nLzfG/ci/5732JxbZ/hCQATV+F1mjL+WEYRcEDbhH9lj+02cjobTtruCtKWyaVUr
Qp/5OU1uYpjE0BWjTnL7k24DMuJE13Fb4sJbMIK1FULMsKY6DhvFVgtcfBBq3cyiEqQ9JHFS8k73
XFRq0qMf44L8Bwyxjiu2qyzTRa4h+YaVIqQ/mJ/4t1dxgAu3FdoLLm9cmC/3T6cQ2U8MSTpDpRb+
sy4gIXZ9Jbvb9LvySW0lLuctlWyHgRoGhdTPH/ad+8XFDiBDwTvvzm+uFvtG6VcKRiHo7driBQXL
zXVX+fnqmpcdNsJVnlur09e4kxy/QGyEJcvX+a0EzEhiOmPC81qw4fyg69mhwF2oJ1J8YGXwiplT
Y8wtVCJEIQ8Z3BIMFRlsvA/g2+U9DUtr323XA0plfyNjrhP3WzSncwsiEvEDQzsJ5JX1EBcxKDO6
qJALY9/jk9QuIwukhnlxShBl86uF+i7uhnd4pBuQLicHDenJp3wP5l1DED1bhHjBCbn9BPXQm8KD
lo6M7R6arXw4x5s5wXHstyVtf/3IrwQPzBdQGXhLrVZE3BuD53AoXAGiGlOPUt1cWEBgH8NiZNd1
BduAwpjnlzg0AzhnTsrCcLWHcuLJ9icRxyaeOtne59fi0+0gOdboOKnFDwqDikrF55clinYlxuFr
HFRpCcSz9RxgDr7IE1E1Z8LDinFNJy6v20ctjPthWn8ifx1KlMWmClqQn/YGK1AhZ6TfgiLLs1h/
Jp0YjxZcAL5FhUAoyU4/cEQhm7SqcKbLkg5YUUKzgiiWiGKwt9F698yIdwUGzWn+B1XhKjTrtTkh
eyKjC6qMsdPFMR1UkYEh/5RGY/r0PXGftIF4arL1GXAwoL54EJp1xePfg/1mJGZNOMeIlYJyrpOi
ClwQZxCoB4oMuTSHsM/Oq1lW3W531UzkuocH2uy1Uqlutixy9rZ3haoF0RehAQhlhqEhcYXpoxhI
l1qZESJhEEvl650LPVFdkN6vA5pPByAzyV5+rna7G8dtzihPyaa9TKVJCJIMdPIuPXJMFdZDVGsW
1Qn5w6U9IqvZGkR3Yc/V9gu8Tj0QLI6QBEvkQvvIAJPb0NQqJJnYZP/7V4ARtUK2m8e60VajkmRR
7k/pNhMxZojMaqp1aIzOWvaOxPP9sHzdi3YRkF6HO8O517RdbWFOZx+cXY4pr043s8lDRdGcOi4k
lcBqyqCr9A2rwcBD2RdRA3FpsL+m6RCCXGl4++p4+z/nQ9gze+hEB1nmT6vDkS85ZOygOsll9Fhy
riU9NgD4vxMLGGAR7qtIFVXPjkMZayIEYpPkmmN5yZI4IvjSs5OiC4L/lkLaupYYNzex5IGozYQu
afR03jg4X/0HzQePMygk3W3NKHWo1AByVKS95ZCZwUN3ZhO0XNhPQLKI1XnxMQbCEntcmv7OfuIA
+RQNFNqD5anI7FwbNfWTwXHfDtqi9vnRHSJ87lv3QKZ1cRuEFdZAEFTfYtFjHY3hiXksmuhirtxS
WBg/2n/wt0TAt5FbDV0FR26BjGSPxvd0W77NmJNai5FJF0jMrHVzyhY9RaNWVHGRRG5oKQce3tBL
le5x2YIr+8DDmqIZXfB9Eo6RwkYmiMkJyl+FjuBR0DVQwoEwzSDe1xWs4TfI6IDCC2+PI4MCuOfe
QNS+iDEvQi7EDTVNshFy2i+3nuxAkGn/6yshdVG9J49spo4Wpb5Dbj9BYOz9BgG1cJ3TSeyDXEGC
7xGD36hg598qbZNclHgNe/gP4u8oZtLF+Wgn+78SNC5JIA6GsZIC2ACgHibprPs8cdmBnsSfETKr
G1rdZKWgCbjH+qwHadnyemjY9gZlGb+OeV0SIiji2xOyz3GdJJ07AILVNxGKSHgxZX1ew44UlnxE
nyIkhyjhR+jXk9qSpZiNlf2jgRiEuc/wwGh2U01g61ZNbzRP412ivLj0WtN4iQf8hS80Fpx5NU5v
SRuIXkRVMNyZh80fLRF/ZkpfflW6GGA/UTFXrm/Gl2X7+vNXDtXRLeSZq6OM9NVh6tkQ7gBE2fBJ
NEVgf99z42hrZXhs7oOuud72nDme1fCeQXjuIMyR5o+y58Uzg+9+De6VLbnssrrReWVQ4y8D3+XS
BSML7HLsIvj2FpQ1xru+7QEfZlO7MCHTmNz80liydBbBPLSQqREth91f/5sRKHD+krtU2RZauqNM
z/Kf0wGeaQ7pclkxnEdsbw1oWohP4Gs82clROa4oDqQ5yBHKnIQw1RmHSHfPpUFrKQO8XOHncp/z
DGU5P6nrfSQRcnneGXhBFGOX1rDLzq0NhDU4nC8xxqUVT85HdWX0lsYs+bwFI4zEZyN278JTXJco
FVIbQEQc++vM3Rb+PK7BlB4vIw40qC4EYxk5N7gEkCStXGgjy9I6+rIgSkEpRHfvK8Jw4MYrhudd
lGphwgwvJT7qApsxb5L5GjwSCaTdCuGFIIOSUawUzmJgH9CJcd4NVVMInD5f1Ivb45ff78PZoNa9
+7oIhP3fyxPhIUDQ18bZSOPHLhDBgUxdsJ5me+o4My5mX6eYhG5xUYyLHip1gE/wXnoT6Hqbr4d2
C4Mz/iCVhWeI2B9Jng2ycfmdY3xPPo17rnsyBDT1NHWOjvuc4K7sG7G4WX4J0HYLgld9jzXr2Gm+
R272cBcf06Qur4ZlEVPVcOapICznbhAvKR2J+tQslaQNL7ItZBxmOAKUYZ867FwfvjTna5O0LC/e
Bg3u9pMqpqwqmUqff0H7vBdFIC/gYP9itO0YG+HRaf/H9B/TnzVkX1IMF2zUPlB4o7Hj0ct7925F
MR6euCQp2UOWctRu1h1OKePjkTNwzs+LrEgzYENnSie1v1sPpCRCSGNsaRIYXfiQTOXO2UoG1PRm
q+FM0yj8PkYD3pTZjanzuJtlywiOro19iCSRI/WykzVhuQfLEgO0S9MWEYg05XT6YIZAigAaB5eL
m3y6mzSERmpxZY9OtFa9f+xrIsWKtV5yZdOTDNLXbdv8y1iBZL62ONdNiIeFLpnEMT5CTbkCxETy
BXGM6kH/kbNouXm/zEIZuibAwkedVP0MD+od08E1RTzDOL2Ub9f5TBD/eBYsCoMekyhvP/27uF/V
8Zi2zJo3YiayKGQlwYOjigYsqVI0J7GLJI+tYWOqYmCAedQ98YZr3HYliiSu/lO6FksopAxQLOeu
y7CcWw7NL3pE8RmXxMfjre8VhXND5w5sBGbo7DbULnu5f3zd7DvZTPyydYGCeLhTy/ozrLXX5E32
1+aqnngIjcxwHPmolfd8/OXBPPs68ZYw7rS8p/YnJhd9ixlmwonJvonoMuwfKFQIypJLwvTSN1ZA
U6cuSLmX2ZZuCWY9Os4ZTvLQLyACfbw0waCZl3YmRx0hksV4nBBJtYJS7Wl2r7qxCar3y8C1i3HZ
H5R053GAG4MsMywfJy6sVJ5SyQ7N9ErqOIG8MfhFtl8M1VIGhciwo8EefkBWlO0nLppFPZ9lSYxN
psU9KjhdXeMab6O4SJ6BvdNsijb6QBIV4laeUubjBvZ+in7ZJ5QvgynSkeFt2ourHPuJa1PpqDzz
mpqI58rmV6Z609h93nxPlzi8AFLOhwNNrTMNtxfBhhow0Mo1r953NHYtHI3qIa7D740jCoDEc74E
bXsVi4xZ0HIYEi9XBhAODCr1/cJ8sc2dMkpt9MYK7sgVf3fFLYKbkKPIwo8gU0mwz8jjgSHSe3mA
RI9ohSmTrT5MCdsbmf8a5xoC9CJRyeb/TbK37U9cK+1NnzQg5TCoFraMrwPaIHFDXLajZI6SvYIA
ZXL8MkpXwmeSbrM5Jmr1nCd3irQWzjV18ASAJNGthZLcRIurGOSMXXw/rjwYdiU+oS3ljL4ASiX2
o8SmxfrHGCK0wqgnz3dWbUoQeQFfM9o5NHXOQio0mLa7MBtslmMCeNWSFfa7rOZODdMc5+sHdp7s
QmjbV9w0bR5R2nRaNaZ5ZzELeSKbk4RMFr4t3El2gU9nAUbiafzNMwkHOQc6rJw1yNwOsLz66mMv
VIxw8l+SQsoVBbwlRZcH1vT/bw4zmpiNko41d7WJhMYnRattbhSuoTeq3kRmuiD9rcVl9NfSn7/w
nX4Fs5ko/hCalgZO2vzVCjrVGgqxUjkgR03d/BuXSlka3Dd94P/f32qZ+YCIA1ReTYz+OQL5918i
eQHAiIRF0/j1Fla7PER8/M8ErJLqo9fNTQUgOx9oztr13YGq1hS6aua6FPDoNXoS46LThJnCDVSJ
wVkgO9f01xO7JlhHCkl7EFnPA9LA3jhS+IUDaV6dgJIP0HISfZyz5+ImlnOaYPrm8ikPgo9Iq3d6
nJuPSuMVNji0MgL/wPE2IFF/B9ExwoVWoaH9PU8pNDay8O2v03BfscMUBsHCHmAd55FWC8Rw1zJv
VchyQcT33PWObl7tnMA1f4K1gVDb4Sk8hsbKX54WiGmf66w2TxbIHgU580reG8TD2GZUxKOyhrUY
snNrU4xPF2dFy02crJRHBCyVd0ahHhkqDhwMtmKQbrKlMW/B0+i79ExlD0ckwzOckONVcJZTcIJ8
ULcacZbBhQxqPgZXJqbCvg7RbSIruDICi8xnZL8+FETLHs16JRJjwP1jq3yIlVQdcbseGMPfjz0K
6AmXZyVJQyPcTgvu+0ng8Es3TvT+OQ8QolkaSI4q4GfeB8pIp44WVx4idXzsrL39BPiX8y243HBi
8BrQnnLGGGF1pdOFLlcmC+ALhzfhTakq0qjpydZvjWTyl6sZ6CcqMCMQMXeltAy8DH3VMwU8b0yA
eeBA4TY09kmL9SN1oVQt4NrIHtrAI/TsBU1X3pkRxRG5k8ajsdZXcgdGetS+OESA7862yP9/UWZ8
75NNVKVVvJTiivGOT24Q9g8649teqRZVTg+csg1jHaTNXIU3uptYxKqfYxGEF2doczSHu99ijDwx
yqw45N0RyPAENVMZcZ2Yrg6gxbGL/apdaBob1B2N+qHRI7Z6yO4qJFb1jgbiWP9PvhKjBg088eBd
PcePSMKW4evpgxKd3j96IGiZcVcnwnwWlbw2aW3Cvjymprftp4K3QTOryyKsMzTzKP/UdyNhnDGA
FvQDlI0NFoNv37Wu57uB9Q4J/czvzAsHbwojQ1HN0xuNZ0KlAKKUKJJI4fwPCFlWXYVi31g6sdou
f+yq/uijPtSE+R4un0SP2CC3oTX2RQU7xpibzQPMM+IVhcSW6OFS24Lwrs/3wUvwYGzAB5iMo+X1
8/ZvY0hRxncMIhB9KofKJrikwwKljHWreQ0xJUzYtbM6/d+eksiHo98soefDCCBPPOGvJrF+dbNO
MNVpRzAVtySYrABC8txxylP0j4Ts/T4X4kb9/y8ypgfkG3aYc0D1ntC+o5B1SeaaUA78JxzUvNzo
/2XqZ9XCNDN1BuJ0Bre/abYC/9U8hGcSr2smtPovbyR0fw5UyFSpM0eDcRrXtdeejMPh+d2O8BM7
rT1AFaU9Gv/vRcZePic+4csYDyATkUoiQSL5rhga5iXRqD4gfhwm9bkZPKnkJ+45FI1N9E+CAw4l
W7Us807VBX+IQO8fOUwkWyV9fpcBuTN0jNjCZkRK3lYxU+lzl540a/R+HjpY7RoQhMVzwWeFQooi
n5D21JSCg4pY07aZF068sbMQ3OOUGi1NOG6w/ULvlN48C4QDMDJEc+EMHN5yBov4yW/l7AGwLIPE
ZhAv9FdcGCGOP89vrCdHBO0eJpEV86CFdEqvWsQvvoSFgn8RE32lr4GL6IWrbB2vCx3VNHOQANYu
NDS/YdX2O5UqMqKWxZ7i10H/RvGE77IwV7D0KU35aMbHz6BnVWbzPv5cYwUe35lB/kKNi3bMSnX+
NG8Z1aRfheOY9tD10KKF1ZQrDSk5FtiuGKzX5As3dmR9qcIlCLWVSc7bfa1abykEabTJdVsCQZih
twOXiIMpZNno9qqE2i3ZLEFlvcSoxwfWvlOWiOg5YvYYn0XaLO8yQ189gXa5rL1xBe+xHhqaHO7W
XQLrBTgeg1FlCCto7VcAQhL5GrcpJJG3CWdytYEI7CIPw6NqbXeGbZObe3vM9Wqwr/0K9CAqu9oS
I0dDQNv4gKwLOscRQ1eVxbJaiaqQfFzTz5BwOiTNKcPJGTy8bqo5FP2NV0Gl8JN4BC4uEkoKTZIE
0aLmTLQwX+t7lHmFjZse4rrYNzM+XtaWH06N4NRzUW7ho1rZkvDvBFLA/eAL4sUq+Yujsyvbk6A6
fZpJC+E6w7wA1ulMP+6MCW+EALBsI4orHdY5zEomKKXVRiF5uopglnQ8KYubvSL8e7nZ3RN3UDQY
esVZm7GmsTD0iyoIuLo3gXhlVmCB/Yw5nkg5BnAUNW3UCkjBGaQeVw1cjwm6fS3xgqQAHKMl8MeB
JfbFArWinZQwPlqCMB+A75DHypuWxNw/rDEHFX+nBR9ogMLMKUgeCvTkSLdf1gimBW5iJTSoCYnj
g1Ef6+CYQ6yVWXJ6VQ0spIZrchoV4gfSbQZSlvoe5uEvwPK1A4CIxcYmzDuUHyCmKyO7eHG615ar
6Wi8VbzUPsqTmqr2Bu0bBklViznx+YwBbnZF+hXp3APTAPDpfHdu/oR09tLl/uIAwq8cOvnVDDk6
JtUjBoHuH3uNUbsOzemxjGIvuAO6SRdFkX9jC0tlu25H3jL3/cyumHwRFnKcqZO5kblW+Q1xoLjD
yUTn3g7mKEo68chexinjhgjZa5DhSXslSAttmrZF9Vlt45S8oBdQNQlH7NiCJ1B2SJDRd0G4bShm
7ZaZBj2hmJdph8JL9ro9yrdATHbOWxcoQvCfc6rYUTZ0l2biJbD+qGnhBbXb5p+MeP/8mK+ZNMBr
3iQ8GKigTt1vQQjXxkPL4sGbI5WkHzKzQkt1ndM9wrRkt0i9Hsjdl45tXgu8GiCP38B7R8CLumQ0
PSBmsPSeL+et6meVdCGtuwnftXQPhIGPz/cVx6JNwxrLwjcfYQ9jW/+vE0qNnqIWe4ygvSByeEFX
1JZxJUlDZp4P75xyav1aplw0pmJoj3UGMRw7L/oy8bHE30eW9vjM8PFwhXNtWvCJhNIp6hhtD7hQ
Tg+/kMtzEfhZsclCDwB4pYTnCk6/9SO2/P2SWrRzsGfa+1nwGD84Ev4R58Nu7aPMRpsPIVlObJ+v
3I0t8SV0p8+zVzdrsesgVRAQzhlP5q0BmYNYvnvxCKu9w03/cJ+xXclQQV+6s2ybw4h2mF5YQ/YY
iisO8IePdy3V3vf4g6Sum457INtO+lfCjtbCFCH1Lnkhhej4KQaLVw4TOmrwu9F8AuuGJKdMtXom
/35mZ0Kdri1f6qmDCqJOm9LYyGxFEEjR+jVLjO82GRXbFgDm2GDJm99qZFSQhSaIFTqGV/r3rrS1
H8VQ2DNYdS7plObcSXfRnMqS9FjF0oBcoTpvn/3ist5jpqBxxJyaE987YmEDArIqBkCjnpOJvPcC
XHS03ry0MmS4s+ijMICWoRyL5eltAhxZamTnmaeg4DSiBusgx7xXUln9zV4/Lp+xiXDUuPGXKET0
OLSg7+ysDNGA1G05dQvWJpoCVBhfnjyecn0usDymtsR2Nsd8nTkPce3O9AkP4w6QcS/nHxPZn71H
ReT0yGYVR7nazQcFF3AikZIq/gc0P15MtwSc0AX3kVXKmhTGBSoHc7q50Y147krTUF+YkQGkmb1b
R9pqeMOXmNZTeCxZ+xOnb9gPh9k9OWzr/25DHA28Pu1we+u71r6cHa4+2T2ABKUNeQgMFpalyr93
6kMx0+UOjya7KlLsZxtA0kFmBIIQpmlGnmE+/hU7vlYAOihw6XtQBfAIWsSf1iE4l0XWsa2lK+/L
A/SK8IrNz3npRi3pAG5phplcjLlSXlCwDRiCZ9trOgxclHGUZNAT7SWFqvlX8u1EkfPQfwIaK5Ix
SYaA5Vkb0XJtyHv1xqtibxYtH7eKaq1iuQxKJqvSLY47hA9i+Ds47ye0WdZ/3QYb4AJoHVCoW0/Q
nQRKCG6KZLCxjyEpX5NFzEGXtkBnPSWKONbX9rBLwclQc9yb43vi8rjf5jVjwb6oMwE/PMCgDMXU
zujdGQvAjxsxCZb9Wo8gapfGasHyFy1pubyQEnBnG4OdK2kXHjjDBamhAM8PI2q97GAf4uPW+9Rr
LWyANMn7WFvfwePehFF+H32QqUsEVNE04vLDHw+f0QH7/6W3MlkLLhIbuE27VygIhW2enGWLmIcf
ezKud0jNTmt16SHYxN4tzCYTt0iOL3Eo4TGOmvCHKxmvlmqBySKPLpxXSc4UW5t/fAQG0nsMszqv
BCjGReerPU0f/7cy7cLRTg2lAbVfVZC+tmrU+VcJ1Ps9RIBeU2DcVEop+UXqPHQeeTHJgr6p1KZO
LieO/woC7VT+UH8f65sd0gT4sHliIonUCdAOoX4yVQxA+V/7PW3S3Nt18RNk2csxZEvYrHh60uev
HI4G32TdtTTakFy99JU+bYUf42dfZHYyqNJ96o0MFxBNaI8WDUPHFabz/DSHPpYVhh0ayW/kQUNe
Dz/HwAca9nsatmfBCWONq3qW8ztYpNmcyu8Wsu8ifhtJIh/dz1oSPQB1+icqM1mQ0ld0N7CbhmqS
z9abNjBwCRDnEqwFt62z6MwXB7epLL1U8PNGjd2mqAwpybQTSOXtmdDKhK6MaJZYZ8wsPUM9GVnz
n9kyrmRXZXCNR6YLBiMsIVwGrJ3ZzTF5dD1D/y9B97fMnA4/0fIobEvFZuyIk0kLvcBh1Y/JCPUL
Az14hEfdu3d8XUNJf7UgzhHQrCDZA26tHIc9TAF/VLN+I8+BAorLKtWZJg2R9uMukcHpozhZisAG
lD+waX2vgdkF/8fm3MXb6ngI3+dGiEq/xXmdsulnuw07jTrBm9cc6qM8EltxReb2i4Ywi1QEzKS+
5IikW1iP3TSvZiu3k1ugZqlEhbpoTa2CqhdcmJcMrlHWXaPTFyXRvTOMnTVuD8W9Q1lFVgIIy6pA
TXiyoSBii8h13vRIHbZUhXNtmJeWqOFSMLUpXvaQxTmzvmmJBKc/S1uUmSnBzLqVm9dN0hGuF4cI
zxHcUhrBBciV6IT0pp12bwrILoxIUkknS+xSzzRgUt/cFr+Hpihvzrwrlp/axoo4WAzADUf8AlT5
MBPyjGpB1gzyXo29ikJovXPwK1LJC6A0Wk79BBi8ywJ15BiJS1bP/aW4700b/hbL4YSFVbM8S3oL
BRu9Fh138B2+zxrR9m47apizNEhhgm1ZzkXLgnM389aCqBBtPTfE4zMj2bU+Vjc048b0zHYnAPQd
B2ChuikSyyYQqy9nbffK6HM0gxRHpgOGjoa1KXv3wzTNtmvZzMZwJMh7urbjD7KG0PWF0/XPFjWd
g7BnlP0QMcVKTWoyUrcrxx+0cfcTXhmcoNPXlPIPMtWl2WBXj7oY0FtT3DQR/iOilXYXas5rGLai
9GdG5FxJaJoYDuwWVskC/uq2Dq+AeeK6NKFlJzOxsDaWL843M6iNOKiyTrUdzfcUE/wH2m+bz4Jf
izt5nMMGW4QjlBXuaEJ36izbv5EnvDbuDAo7ZYt3fVFwdEo3SZYxuF+CvtVxDYgWOPMkcSoccBMp
1ahMyjQ/2IKcN2L6gr31LL2q6k7MeWVVxY8joTAT+ogB4Mh1/DsrAJx6y38li+en7xKgByCd0Z15
wCLBxvVFTXMXnMBM+CBYRBaokl+s7TN/5KFx8bnnUbQk2DJkW0n/7d/5q8+KSMBe6oM/bdmqvgZz
3Sv7NyOaGh3FratBzh/+tbN+ygxVKao/Lt5WXEY9yFH+UDjrB9R69eSY/A36sx9i+GIL1WBWM3CL
/ZZ7eJHesAW463JH1zedKlYc7mMQu3fICVS8lJi95ag9iojXOypg8wPo/8ya11pJYHD1huj/kcqQ
Hti2cD6SA+BdzE2jVzlrYTfIvvOAVJ8t0ZR6+3QIAIn1dpDmgztceUVfaIO/fpb2C+O7gp4iDg8I
PzycjTfzzInKkZ34uZhW/lB+DSeyocbIGmLkytntSPcszlAjm1P/ROS5J4uONjjf5QdTCxmvCpfh
/48RoOODW8fOBsRQ2fz8fuP0AoYQaso/O4P0T31A/HFj48Ugk9QdbCe6qlxNVszBhwGQuh8obyoB
t+qCEDqdWyPth0kkXWF3pBAr8HKUeH5+oWTDwaTPUbgJyTAGnNb1DTr4ULFjcBmm0aV20DkZYY0Z
tnDiqz/VSziNbBgXkZRhvk4R+w212Qax5mheZjqjtra+Tp8MqcS3iiDSXtRNKanwm4D2u1vsNEq2
QJfOnIawdQndVamLGwRop4uXndHIMttNI5HzEIjkmau9DNKQSL+voZA3c0+RqRbdDij+tPEVJL3a
qe97GktZuwCcyP44t7ZtWmidhsf2P2MxTXeDYz9ZE+kQx5dFj/qSv+sXbwyc3NNZerSGgKo9kANh
MFkjvItwqeHclOj6j+DgmEoWCzU1eScezFL+A1F5MH4+3lY+uwCKHNMcXzt8E9iQzIErAVGFaA+R
zyrvePutPKMlGNs+Tu5wFEatP764Zj6nBNhxQY2/zEN9+aXF1wgcpxyYO72FtHGbfnqRfuIHd34O
vjhsf7aSMsUClXuOPIy2XcYlkAXXuGc0/z3ez8jZOgYFrSmkW8OsO/QEgRhNA0UeWpvviWUQrLdP
KrBVgk1hHqko0fd8VRELOl97scUSrA2kUNrX/Il2jmFThY97iBY93pT/5bsn36sHysxhAlbejowY
bQ8CqKYsrXPbhNj1FBlzi+EaSS3vIc4Sj0mQTUA/6zuQiH0US562qq6ni2sTeVKjTZOWSvkL8m4C
22X8Vg4HGFSUNjl8yBKMb0dRNCx7VrJefSATuqair7pAYEQtd21iLPa0iGAtqAwRMeJDHhG9U9sL
ZWSNQpS2ypPxWP+kydwAK67WvdnbZK7lJnsj5222D6tYe8Fyb5wdVMLaAe+txJAosV4/xV1Zgkvs
Up0OWealDYiGDGjYkExVjwbDqSa+RX20TMDs0VJ0oy3M1FQ5VUtCtXlaMmfbJmm8eK1XPMlQVkWA
Etv0x0O1L6HOuXM3iWHs2s4lfMCkh0tChzm7TLnzKGfFadIHMcL3UcdxtJGQAfQplx1ypITJpAwT
20ZnKa99/YegjR5KMhOaPtBtqnd9RWTYaWgrVuM9EalPVqPqOKFKFuwW6FKVVX3XdXhFn93CkYhI
wNWlG9sjh47GXlFzutzssFz0YLWClcEUwTZtkauzDtUlOL2eD7eVZwBXWnxb4tJ6AE2Bc+ot2U/a
uuCPdcd9tDan43dj8rYtxFpXY++MjXqOwvpu2SgPUS7zq462RuKALlUmFr8Z0PyjZNEQZxpBYaOL
ymBT4KYSNDVxKlDWV3W7zNLv5I+juxnLXCBggofGrY2Hwar8Qy92Afi9MKz+s/VJ0iwtG4DV8RFh
Z4OVa0woWp6YNCYoejVTuWWhWXWVnG9t4LnuziAHviNe0uMA1+7p+bQQi0biAZcTwSZJH3uXJ63n
Q35ZUr+2PaKZW0aV+QdmttZps7KrdXn0gHDOob+Fpinst0Pz2+KP9a14O+pGRot/BRbuvmaDJcGQ
peMeBPVnGQ0agcRSZfO53+a+BBtzJ8x6xpj7+lc81PNaJqxTBLiFaBzx/GRhOh9L5QMxeaYCZI0y
3Q1kxlkUKtgVT5bohc35vVUyZ1HFpfeY5hnp9TYKIdcuFoLzHdEMeHTz65aJG7L9aZKqF14EiP6a
Ueu6mqd9CiDiBmpPNkIkA0Dp9OVPKJjjm4ke5rm+IeSzkXd1RIHw67YXqCQ6EIONCtNB8ntj+FmM
XYBQf6Wv9R/dVdZnigeWOEoRZnkvj/R10HzfZU555am1f/ir/wMia2bvPu9icsc80yzP/5L9udSj
wx6MSMaNFmeAEncNX5Bet7OVDMrGWQhLsm97uGziPTFzXMTQRTbBVySNLopxnMYqk/tVj12YfKc6
0ko3GgU79BDFzl0qQo33tscWemhMELEeGVQBpPrgLRjd2USH+Holvn4HBxSx8Qwjahjc7f6V+9xG
Ic64mehrP65vFU22h3acael56NP3qRnzE20N/p+o2l0TbfVboZ8oxcJWbNLmwxgd9iMJrEH+UEXA
00Y98dLjbdwAU7tWFchvNO0ONcUIfVySPxBex62HgP4gg2qOHhh6+klBzxsQoHTwJwGCdf/TwC1Y
v1/cCq6+SmD6vnozDoBohHzDHeMJxBwqsbY8NV5Lh5FPIM5WLsMYqiicDZa628lIBYh9T/g4S8mj
NyhotdCb2+UzIRVW0DzOqrEnyHcLp85POpMWkDcl414rX7oNGxealpdL/Xy8y+Vl0rQ5n7iQ1Z3A
IhXGCOYAGhFzvpY3kPgdGoS4WuSDLnPDiNT9GvxYCZ60cev4F5/aqBYf1wPZUANqsF1NZI/J5CYy
nvQBlyfP1/OTOySwwm0uZC9g4k/fYvNeV6LtN3JbeawYPqLYhrCOjedFffX5mbGN1qnJ+dvVagoP
B2KkErt4SzlXbFtf94VDiAliM08tMdVs7wMxtsj7K6K0/9ktprhXFVzGLdvPLlrhRMQsbBCxhVlO
XD9icJ6BfKOB08cNRY43ULZC+8bbHt7Z8OzxB1WV/Rcla1yjhvC5gAqiH2Pu58MkM2NwhVpPYEbi
2Q+Wm+d/l4L6U03/seWX1uZePSdypGlmzCLW6RRz3xXpgnTXb8ZkJzEMJS1XHOnJOYQJ7oFk4CMD
TZHajwYLzf8vyb/lArewN65lRyQlnKJSN+yMKhCC02HlloEOvOhLL5sH3A1yTgMKdiA4mI+37T4w
HKf0pUncoSCkoNqspX4YmzLSgQ3fzNoBS03B8owCevBrGZT2NbYIXeUz5aGgt1uLSHMLn6YFaf9i
TL20aClAJa4zQYhcMQjwPqTScc6ePsXs4+WkgOM/ZRslORAS5+iCDnM0ZVxSrrNVHP4uNjaEO7fQ
qdYYuLSYSz78cWtAqWvO6VO+ABIpH78WWEZv8K6/d3JJR1x4Qh4FHow4xQ9HRURwGTb81hmu9npL
55VvF/iTg5AF1piDGN1BA8JbRuTrAb09yFBBoiQlyrv+vFH4venTnNcnO1nzh9TDBVVIZiwt1l51
UjBM38hvh5gk0lqXpzHuryhqoR6/p7i+ub2AlhmIEpYgGdEb3lAwZJCXd7zmhYQf1V5u4jAJGdJp
8fJKjBn92yP1oCYNDOHqxtORRaCW+lvMPlXK7Gji/Qi+xshXI4k/oDF/1Ni5RfO3Vv2atUt5WGPm
3crMBpbKW6VHNDLuh3E7uB2oecKExJ0Fqrry6Ghm9ehoqIY/9jOEClk4DT+N3PHVL0K1l03vdi6N
68x3IuYjfkl5ewlKynE0Wxh/7PP2yYhrx4FzBx3Zd/KChhqUYiqNDppYp6fYEm5IyuE8AZQK1hjM
kkzP9LNjKTdNiYoaorVRm6M6pPJqh1im3JqOcxWvz2hrcMoK/JnyvdE16aqZ+nww71BjcDH+FsGN
woqqnZ7f9QVYgw3MhF9CHPi19CHF2tTORPKq268yRXdSQ6+RKOYXXCcccUtW6BTKX5/WAkdj1c67
D6bRFFcq11m5lhI9QVFXlmJjhcrI+Lmr1dqUG9I4rHsGXWmHeqA6hlQ6j27vN3EdlqhiNuYgVdrk
dxPUV/sFCpG5zlt2HUHCvKFl2v5iHUvMI6lsqiETIp5gYHbvV3U5O/NffbIIhqLF/ZS1Oo4ODgpw
X0UvZtAsmFA426ocG59uon1sGwIvSbUmpEIDsFGmZK+IWcOuZBmI9YXXkaSOLnObWJISzDakc1aP
VTvOI/ATNClA+5/rv1o7UK3KxqQa4dXWGrD8LlLOO6xpD12YFmZ+1ZahWyJb44keZZpSCf9Z5vJ/
o42IBgRt0NTmwNYhf3Hjr5ao8ZiY0ohrFFJ+TVp9AQNjisu5OYJW4EJaraN2k9Qg2JUBTth6YgD/
xZ/Q+rZswqPnb3h4+IHHF+gOY7TECl3aXbt6k7m/QvCx4hDN3vAJqXz5RSdtrO81MDa/C+u00y9y
YC/D9WQiVGjbjUu1tTHun9gKjCggd8CI7UFObxEGUMwDka53iaHQiPQK99CIFLQZtCBF7a9nxC+y
jJ0hucxJzQAVfSzJ9Keq/SmQBArPYEjyflM0i+wWRGw3qjDxfWd6M6YgR3+UKYbs3qfcCc9WUdrC
XUfGwhD9pblRKCQcVGPID6tLUgH1C6/HQzIZL/b0C3DvMnGJKGRsPAlHAAmnG0FXMW6h7zhKtzLt
FI6QAZghNYFGI/OS7q2mNSQ46I7vDowOHFVeZ0e6q0txCI4+r9lZUDXKKsWowSSXqLFEcRXahXzS
Jt2BXtEGsdPfG9pygTtX5Oohoe9V1CqJdSKXaCuvYSwBwOkNZ12qOZn7uBDLWOcevzEAX779Oq3n
iPuFiCtZcqL+Y/Y7PanIWvjlnnncr/+qiHRQSsYvR7qsgwKH53NBTjllkEsvybXQYLrRkt9UEQjB
oV69qAVCi7CXTxFzf3FzPoEcrM0MITaav0L2900QijJBPUvkJmD8IQtUX+wg33oxtOfUK/xHvsuH
+99+LgrHwp2CLdLd6+cszIEW7P3R4hQemLxExwAAitcL0em8hOvoxVZUAQeQWLI8Sxs2bNKKIXYN
0Ask7PjIkICE0m5AK1K5lODrLj2lSzlhEU8ILXbs4ZBVO+tJbkEXZADG1+MlD4ROd51+xWtAlwtn
Sd0OOCoDi5cfh7KrC4CFiuS8EFP2QTQ6CtkLi1f99eTm4KXFoUnUiLEjZE9788znKgTIJHyXVgLU
g1g2yt5wVMx/5mIufOOeBLE4BqdTQyOy79u26zwfiJ87LG54UJsTG8AxwBlkRR+/iqgqGaFbjwd/
kgk62kfhKUF4TNtDoNtGkk+DDJK9m12/9IpcUdI56CSCnEO+Ntcg8YTIQpQUK2uXsZzDyi6LBtsc
QvSRrqua6kAZD/1hx/CyF2i2YRisQghQpYyie1UPKDq7IaEMjtB1Ftc/xsyL7n8hUU9sj21iiJPf
erleg7tyncxEEDnbwrqMdbK1vHA5IEhpz4nDd3sSugCIp1u94AniOL+oz5DS9h11gHz6RbIAxHFV
vPYpfvjC6O8OgF68vSmxaidL2bnn8zdScpM45vifgrF1OrnkyM/4W3HwrtEijSftoy33xHlW5fqi
rs1JSNsFdQkc+wkLU2i6Ve2m10xIFH2wNmu50hyNKE9PPbsjJKUHWUd39NsG0hxO2t4pphHXdZLn
K6h6T1biEUbmmTmHzLbQVRE3AzFoJT89Z6BB7hgWX0L5r+3eNGwDzYwHf1MQ/1iemnIfeHoc0Lmv
FY3CFSufFGYsvovtBOygu94kTiDGR3f0oqJF4qiYiGVEXGOUMxpOhx6JBUn5gsZ7MFv0Shf3R27y
G0z1QCz295H2p2IDuIvbuhfyZHMzVrJV6AqjJ2doisFctQX4etpvFhPD9LpXt5OGAu2tV41RSNih
pnZ/1fTVfXnsinA/iUZjR+tdj8lrP9YEBaxK9PE7VEhnFQqzZPC2UC6Fv2GVCbQtRaVWhetJiCVJ
miTF/LK+tXgJnhTqwjidhlmHSz6XMUg96niNdt5LNCDvsOM/MduN9+HARbQ5PYflX3OL7NA4TRb9
etMm67M+3uVVdM34drPKBLYEWZpDU+WyY+jeb+o9qDlsqx92CK1bOCeeSDSN8ldswL5vR0f3jlFR
P22raJjTRJh8ZouxtIPU1ANFSzwf+QPiyPfl2Wk+myA7QCGAWt1v4rYApYJlLyNSSYNaBbTiTQJy
L6SbCOOQfm8xVXFLjrByaUrCEfMWhKAMwSu3qXb7B8eAQ1NdVQTw1pxC68HunSwiBs408y0ji69w
sksQgiGRkgGfrgUBeJaxY/f3GA0r925lNlbNfao63OtQLugVfSG3eyAgsKiqtlssbTPjICK09aqc
+FPcEekF5xMmMEtsbg/A1dow/ypi/xv62AKg/a1sXJOaSosUWTkyJuyr6rFfqvKLXwhYGduY/RLA
+iZjvhYgxPcw9FLylCdLpC7iRD5t9X6KKTunLYTx1RhLVYzfwU/TXguyA1iO3CPGt8v3/Ye4gvQV
dHdrxccPBKUU9gf9arnyCNsBPcp5/W6B9K3BDuZdBYYDxD7N/GTsIg8e679m0S+z9hDUo39ucotQ
Gpep72NXePV+Tx+zAgoSyvl+uZITW7UOneKBuZCkFXDAavRVDOEuGBphpa9iUMlz9wXFv7zMs3hE
cnWmo/b4VG6Ql3RcreQmki9OH0rcWEKB37CQHLnZi1FjqaqSXnH8DynAvHfYRs7Y6CyN0TXn2aoL
K0Dclte64VynFIH0fOnkEQlcV4NzwepmXZvDl3k+KPz5srjNWX+rc/STnWtur710ipexCqaR7wpO
7g1XNSlnjwuPBrFiz7sTAGr6hYDYFcPY4+Nea9i8OaXajrZeEUPsfPZc9S/xRLaQVJCDDYN2sxcy
iH1ZwiaUmOSd2f2u3kKYrm6lfgLOd8Cca24tvzN9Ubhe9KulRc7el1FWgJxgRIHXSEliSWaVg5wT
mgIC+ZArWYQfdDiYR+CQWkqh2Tp4qNyNVxcz2blRG2lfZyqHQcVVurg+BuGDwzVxo2io+ko4PLWF
jkoyvnT9ZeMdueezJrAbBdzV1fNZYwHrgel+pqB7bZyhlNdYjkgBdKcFGdVRl98NoRPQ85RExNhr
lzBCXYSRqj2MKJI1DKrsGEh4m6J/TtNzZjrG81OBEhwAlhcBL1QtldRTXCm82Yq6dwVXWVR4IYbD
H09cGvCkZSpl/b0y4fpc3DxMy5y/IefllfdYc0FYIn+JWzwGt0fylpwzvdiA6uabpGhi1OlF3jRH
rSdLp/iJgtzJqCGLYD+X/wf0EYwQ+C/Bh9ls28m5ScD0JYlRiFPjbCLD2qdy+yvENH6svfnVvM9w
WOYmwhn7Droau8dRncbfoiWG4ov25tOiycaDlnd1+aLSeP7MOi7SCoptNQDfLt6aGvjLNSP8k1CF
ZnvLSgqIFWHZ/W7BVrZL+oih9b0ZDzz6R49F4Je0SFa88e2aJWnZkY1zQzHgI+qfKAoywn+IJ66l
OKay2eEqVgbk2RmEeQ6jAtIrk5tWfr8N6E8Pk8SlErQQuv9EWWSXkTfuGjedtRX8DD0qyeGxyvaa
zMmSr2e+wIsgatZRN5u5jmpCu2OKFyulBBWk8r4umqwFwLQEsdnVXisKzS/jiahdLNmFBX6zZ3qN
JM3aSgwMCPPlYgEQm6syIl1LbDNOh4olGNQDa4g7XlAncfjh1F89m7doOdxEi/HwUOc9cMFbes8C
d9JMEctR0/zc3VDg5gHDQjao4dl14OHK8O1IQ8RcBVl89t8TQUCcaVitQfz1UEsHhZYwo/gQhNcg
gFergocs83c+o91Arh+EQdyZIOxBEQ7MsEKyXAUBnsI94Y5DPG7o0dskuDmpnNIXx3lL38dKmxCT
ydplEURUXPnLMd028r6spoa5M0rEYsIwZNbE0PADZgWHqGtQda4Xqy+zd9lqAVn4V8h597nXEsnx
0eT5k7B7By+S12BWCjfkaCzgoiaJ2sUZjOU4zUIOoTB2MZZtZjFWA2OF/WTDCUclbCQKy0Q9IV9w
Td1xX7/KGVwspvGp/ldIrPD9Nf2cYqHBMKSMPbBcIfPrNqAHtAbasy/SXV0psXztuR+7nksWPjb1
wz7EU+yZ8U9aIcVh9ZPx53NQyNfsk0vABy7SR7iU3xsJ3jZ/RJ7wA3PJEXnQ2meX9ZqJK7ndPfC+
P0Z9NFGGryj1/sb7XTds90tHcVza/3he+EXeRmhF5t9l0NR/poJFfnkanjJvuaZRhTQ94Mm0rx97
dnqxulswEBSYG4QaSkh3Fp7KQoZZ51bvv84wHkzUCchNlCSvan6/eIXlG/zxJKZWkiYIVvDdp7dS
GHjgpjzwJYDLotzcpjndyJUWIbOID60517z4Kg03jKyxr5yepdIA/L6Yq2ep/8KzKNxTRXO6PTk/
RtgCM9exYSSmg1NbcyEGqAg0TkzcTdbPig+YzLhC4eUepWS9xDOKdJB35LpHun1+JDV3LZhc+aLm
d41xuF0NhsRGIO52Nd7QtIgf+UtxcKi54wztVCgcNiMnJ18JRi8EzdEiwdKWD2hf++bqGQKQElrY
dBfErSR3SgqqLor3E55FuWts+9rZO1E9brn/mzzFO/aIM7HnYpoRcAIqMH2g5BOoL9ho/79INSJC
b2ihi9DtWnUAAOF+EQlBtxfnpgZKA2JvELYcpUXuJrAE1PVkJ/2rlo2emZaOhwxUItazTq80oWXz
7MhdUwOpikjsWbhhYTXAgGatLq8vXzMrYDhmw5xyBdyZm1LSNMJ4RyXpuCtKCHqoMBsRsrp4y88X
VRB51IIXQct7JaoY/7Sv6iIaIsSAWiHY0LNpAnR2BczFIu6o33S2Kr2FJ2THbFHbwqLfk6Rl2IYw
2TwU1CgSRMyRJXfar7je9GNTcFB/dYLOTB46AoEDOWWHLkeZkvwRRQVsOwLLDKWXpZPDD+c6R8aD
gU2bTjRFs7P0Qf0z5HQSKyMB3y3dAKp2/XU8gCPqshBgQeEoOAMy/tJT5cnBqYScI8o3CsoGq8I1
jkvaZJqklhhIQQH3xT+b8rrZ+MJxEv3sfdeGiFGyXHDcYpRTaNL7/yzA/gAEzKKu/CCc1O5Z9bgB
f/1P2qQ1cycSLBatoEdpjcLruABqZNvKR7Du1qnieB8/eXnKnMcfjMiQqwQUBPTPVYigz/VKMmfg
t2dC9kZp3uji4XcJ7h3YVIXDsn60xSUAak7QU5E2iWoMOF7sQSH6KgSKA6pOhAGKRWzTVUbYHfzk
21nfIxes/SjNJVCBEYgFEaZ2oL1I5f2cvnWmqpHoQNWLU0D4JG1wUvY2WLUIiHRWMfGBzTVxyBjQ
dR4G5LtPGfEJQRaz8oYRJuFCbIPGAeny+5gc7Zc1FosQ00tX56KeiuRVXLH2gYjrliRivWbn7h5s
xcwVAHVJg0yZp6NoLaK2j2V/ptGJPFCCwpuUhMLxLvT1XdImog1Y9XUtfbwqdny28nUSCt+yw+l1
tVyuflDBQoXNnHglM3F+EvZhaxL62PpBNkG1L74KaCtpV4nlEUhNsY5SJ6BDPaHy66JfnS3E37uN
9vk3nKKE73dU0qYSLog6PLnAGlxXGj8TJaZF5Iy1oX4020zO9krImZbwQqwUzrGMPBn+gFJKjEsu
LClAfwkap0jxvYCxPcANF0Pga3QYZaeEo065paKwoAdZZ9ro662So8dmNy+xjww0a5CSI9qs4Zi7
jEM5SXDYB7vZfDbsSAQ6zxeDsZnhNEYEkHGZ1XCkT8m2I8Ng82lHyrLxE05H98yUTmZZBybEVKjX
GOT+NioSm9oFJlVp4yzOz92/QbHgVxII5uSe+oWAuvSlLeyws0nyuXUpTDzpO82lVL0VNdU44gk7
c7F0xAspKB6noJGMaSz02P7KhhkYL6LhMirPSaL3OEv+hrZmhOJSvK5tsPReV+WaQC2D8NGDscK0
GxIrktwfIoSNokd3W8l4WybFSjOKnI1fAMLUFJdNK/1XVjvvYQ8KiPW4LInXozF6J6HJy9NS5LIm
XTVN3LDhOKvnbKnFwbdBhI9COYi6PPvaFkASdxtIrfl8HwLXVf6QjRLyklUIO+466VxHUDBaxUjT
rMugYw1tOxOZYxPEpcEMYJqY4pkqy6ES1NEPC+nD/vpCgLDcfNyLTsqmOzEcZuUn5sXNsaO/MYgF
LZvDjv4d4nNbSBgy8EIiPRzQtEsM7fisNFy4PghU5fDeIU1jp0Hb8/Yn1IQqdOj12lZcZkyR2ZyI
BD22RYU6dQroqVTb5oqbLyadPm1rsCrvcQPMdj+wal+LNlcHdHEDDz5U8PpXz4kEorcmR00jRlEI
66NaIjemrElLYBOU1sG8AAOvbaF169CWQOkOHeC39tLM4nfY+1wUbgYv6xr+OZJvhYXeyqBlXptr
+lYgakcyXPD8U3wrqDrZ7qxNgrc9uvh78PVTapy3IEV3EXiMieYYhI2GU4B7AqqWEUBj7BJORv/y
SgYCuvysHPOycw4gyECpEvh3d1E24gbSyXxvv4TVSaOV/l2lDr7qFIC+nQ8PvGe1x2JFPKoJ9RC2
k8qeYr6lRjoc0gE17Tx0DgdNvK9ijBecFVcleFFCfhMxMkdU5cypA89nNoTJkZmd7nVc6n3mJkPe
V1qljfD8U7QLZEy/6nInGKqMLsPLjGKpboo/oNR/cuC7JxPGRG7ArS7jxHr5/zyEghCOQtSOnQqm
iGLCaiPVI99jjSGXU2YXsW7DgrfttSUM4qOvLSWokO8rcKvUoL+1sAxDJHHTtBfC1GdBFRzBEywn
9ooCk07Pb9AjpurRIx39nvLhu838bum1WFrSqGVUGcbg73OP7ixyU5brHFQtrJhtAIzhQ0bK+bbA
12J3JP5OUAKxsCS2ivmuG71Fh8rcj4/CDX7zPmSHyewGtNFu5pRf5GmA8RLE2RJHkG8SolzKW3CE
gXwuizKlqcWD9rzxN+ghJT/R8lD2IkzSanRQCmhd11L0Vo1XzSAdNzYsfyOm84HDQ5ak3uGDgqGD
KbhxsRUjpgrSQJJXfnrxkzT1MHxGcdYDhF8Iff9OZIbo2x7ax4T7f9Y6PIDDRAVJqReULTpNH3JV
V15XCMrKwBZ9NILYe0RzuD3uoGxV3H8RHQ+R4muxdUxXaJXzE+W2lCnt56RMI/VHp/MRW/Ef1rIG
cJdGpmgdac4NC8K/MaDenUuIxqO+xNYQYicjQ902V0hWJ7BSGa07Mcr6+b16V6i2SnDhHIOKYRxG
kFMLMrujgWaBv53Inyr1ggdiViPdh/zP0jJU3AasUcW09nAbeSLiFUtc1XiefRzhGfmt3vMsp6/G
DLQTSMhm+zyfIk1I5oyrSYqyjIiQcKAxugGI1FfwNRkV5WO7x6ZkVbr5Bs1p/4Nah2n5AJCi5OR4
DylSh2i6ATJ77HMMaod1IUC71R5jsONGdHSNyMgfyDR4JPXPQhsqfTunDH3gENWSlRszS3iFbs2m
UCrkdRcVU2p9fB6DRWpPYc513qZx4rMe32e6hYj4RY3cSHI++mijO4vS4KlKnDzYhj3Va3wpFWSz
VN92jKY2YDWYo1XJNqEw2emSlz/JZZH4wY81p8Z8/X3MYsF07RdjgSgPiSuPaMP2KDvZJ2SSRgIs
qQBgt2iEFW3DqDCWtZQPOFixRcJ1WSuuDhyHKRj0Gzi6hZ3cPiMvC5BHKCVmPijk9lNPMCmKaLs7
heSPArF0ZKNuJosnL6vv8b8yocjBRHRxlMKVUk0Qb+Q07RwQkFlA/Lpf97Vcjk1c6LczsBpIiVuT
tWzmpTLZYlprcfl1sLR0xohv1DVXHACJQLc68pOn0eEnN3zQA7SxqkM9xtsoLcTDDVBRUgIb4xnH
JQ6jezC3rN3ZDXAj+YwBHt6zDuHeK139j6kS/EAjHykaFq8v2JyJPXHYCjeOvShow99URmHV2E95
p8ZinEJkzyVZ9wE6tcy2pfbrjUMDoD9w/RCvsHdXpWQP4z8MI1Tgv4GrHcQbovZ0jfaPMcEf5o1M
CLewZB608hDJ+FSASfS0mX5jbDBY5k1G/RhrYiEt0tU8Mz+l8myYW+uE6O90MiCrLYoubCiZqgNf
P7Ee/msl6jmgeUz0EvUbl/CP5tjY1JGQ4ovrEYtc5ztKtc0xp0ypkpeDq+6XB7dYT8bfkeeNyXA+
4RTCi78mtHrnShazJxUSsRZuW2fhzN0CCEbFRGNeFL0599G3iTrKbR5mo1yX7St6kyZzK5EUSVfH
/2dJDHbqFxtS/Qd/R6jH+wWkVvSaT7e4iu9p+/J4GanhNPG818SgriqWei+iI7UHHiHuu29IMYl2
W5C7b9PRO3CPMcQ0/Hjo13ykzfIe1GI5btQ8z5xv3sW6iQDHTVnakBjd2mIVgn3oUDlkJJrXCTBE
3CZgxAYaD/QBHrZw8+HV3ENXwuF4oWm8DJ2s8o8DVQ9puJKf/zEdlBSrXD7DcZI7moxANS80wKSz
S3WqO1fLkQoQDQ9pTYmyUOalR3OIeGZSY80FV2zuFZjO68CY4IpF+937kboVWRdqbSvrOUj7TuF8
5d3+Le2imsszVEcm1a4tK6Uy2KetOKJenbhrvPJq4YhlKWSPMxCRtNGM+5Ci2hUbnnv4VCW1aOlo
cT9Z7xCzBplrzjHiJ7C+ZuMIJeUCuBChSUIGib028mV06eBlUeE0gHo6C2fRrhljMpUriNuz/xtD
ZLIML5+LiOVuw/cfb3KNK1iF2ZSU//ifxLXD1lU2gyBMenia1RgkAo04uoXJSVuW5i8nYDL+wJ9L
bSg7Dld/jkTEkVclpcvt8wCYXSVWmTHvdKQLWS3SVVpjGmVLVJ1vA2Qo1C7G8dPx+tTWzF0oPxNr
DktodrtzMn7utRp77jB8YAwvue2c3MIUf0NYObbki24g3EIhAPTIYeBSyn0cFHYAjIhCRLqPkOAd
//YBh51dlLW1nvsxn+hJ6OrkHcIbiM+3D/MyFnTsVr6NA0Bg3wgOXLY8MCqa+NlNx7JjD7eZP1EW
+FpntLJfPiy715hzKfELST4fdAF8XNo2Ta5T3btUsYW3nQrAP3G9ToWW6vDLZpK1RH/rrKxJb/4k
qsmF1JWNDDofQE96oqB2G3r4JL7mVr7rFy4yLJWJstR0tKEOxB7XTxtevATXweH45ort4Gx1loTA
k6HvCiix4Vhfbfv13mg4NACKufP/3/cU1XQG+zU5v9P3149Xlo+fbSnQC3FoMIu/VZg1Fp99vu09
uHGv3wiFxsPCkP63xaBtVTmkgQp0kbGctqGQkzhQy0bVjpBckIwYf7pH12Wo7bwn0KvXNSBcfVrs
xkbg32Bvgmr67MEPJvndWITX6XyZOzCYgWcNuEsV+vKIHoPOnfjxM+VFKELtW2WcW5FzqT8hhxtF
/Txhq1Uk+msUwJD2F4NYSSFgat1tX7zQl7onMt1PysAdS/YpejSufrWhVWRaVxYG9WeZB1i5rzvp
C7bqB5OwPvSILyzZPYJxz3/F6Ave9tW2hRsLJc+kBm86UvO00Q9z5w+sYzyALM5fNOdEZEny+6/u
oqnKtP00FSPuEuZKpytr9KTUcz/GZbghDfVHYz0Sb5RwR5PjpH16TecB6jLWcCNy5EpKCmpcBJnC
JiUIOFt57TCG3Ku7W9WH4hMoU3JDFwo53mYAzEsPvmhMfv5J7AYyfV+RvtJ1nrF4hiGQb/xhOs5r
nt24tf88uuh54dX2+/ny8aZkYvEWu94OH4AIubsgyHLjVeOxxvsEfMHlBR2AkvFm5kuXyrnEcfoD
qET3T7DYq360n1R36UWpfVunR3peb+cykN1Gf9IV/GDVtIQpvDzxXhR0whSmTw+L3yD6uNZl/nbm
jchCBInGqWaMD3XNgxmytCs3dUeu4Y1fY21i/WpomS+infM/3WwB0vXF7qh5ZJgOwwS4efC+dO1s
EQKtFp+5uBNyqtW7eCYhs5uN4FYfXPwUQopZPPmKFtYIXh38dyjRfzTHdiW9lK2Huqy5JZb4fgBF
Mg2bDXBl6K9CuCbGWWwnn/gbBzL0GINx1GNea5nQkTNtHxmiYGJLhOOh7AyqUAgvHZfwPwdjw7oF
6OBLvzaoy5+rALXtZGTsCoGIllDT7IRldv0mKRhE0yqsGOI2ZATmpRpbnIM/7Xdv9enywjQes2QS
VM9yVlUzkfJG5MpD+jaKXD05N5tJfWTXE5uYgIIY8DsrwmMWcD5i7WsLhbTKCuTfj744Tar1RNbo
iYvcTgTdFMj6Tr4GrJoQ6PuJ+wZILTmo2+kHgZmGZM/swBqU/qiZMIinc6b1V95AwuRwIOEtyyjA
kI2j/DMIL8JV04Grxe7SOIHsmZCxtfEId3aXERMnYScb7+tWoB5qMI3kTyXMNJKVEFS7Nsh1c2fH
re5ohvKpZ9cbiem6omHNKtEkxPEdi6Y3jMDyRE/BLxKZyFGu5WVYSVu5cPyfhvNRP/YsD7ev8I4G
scJvKL0C43Bxq7eBZl9PevlkUqKDh8IQsznIh0GnfEc+JDQuArSy/1ETCG1TZQ2KszxDNzgMs4tP
+4lZJh6vbke3r3fXUK7vKOeCfJ/2jGRBxEZlckhJ5HhuxsaiI/IEASssKhN8YoZAIDA1rXtBTT49
bMrawTGZZWesLbl+8l9OQVm2VJpJ6MC4vXcK89gcjb4SMiiaD/ejoTQoGKlMa3p58V9b/THsUZxJ
WUhwdwAZKqF0LvvfF4aRx5v86g0wK4kLViOT0snRmzHIW+ZiQLEo9Dr7QaF5+lWwkXe6KXjqyPoB
EoRcBBEkBtzsn5DcH/MQoy7ySf9DSeFJ3PmtndVI+nUF+cWDqy383rC8B7NOlwepjTszJfp8qIBj
VMms/BDCb69UXeKWvoAPfrd7m4Z4pNRvrQWHBSI7nU2SmdudU5L8qyHDnnQm8bUYuseVp1+u+NaR
J1DfMyYP49GC5yLQV8vgFOeY4kJtfDZ8ckq9um+4tBy/heHOjLijSvzSOB//J5yvw5CUe/PhkDcl
BOlCmZf7gPQZSZZDGiAlr8JkM5By4OLPG+JvMJQMhv9QLGf49ftw1lplJW9KsyIgCrj0lvphp1qL
W26fO2x2udPE9wQzkXbhNry6Xmsopw7jJxePFOpq7jdwEfBzV6FbGcNWbI42bo65vHOQB2COFe4C
xIj4t1kRfYGcUe7/zlwAVPc+fh+CYFUN8X6dTamcDeQrBS7RPKRjuC35yPK/qsbL42ZgHWWTSzbP
986lnyO3TdN2ArpAYjwTqKkwuPRd2vs9VtzM7dB3hbw1AZaQalS8cbybwUJFbUa1yAEwwE+1aaSI
RAwSofwlZQOcPcUQ+lZHeVxWQt9Ue/SHYgTnaI4oC0VpCg+k2vgjaKULEmLEyW24XdFStiU2nPtq
YqJ5e1+wra07J69TgGSJqnFsO0nB7/Uk68XzadOXbJ8eWUaMInTHXAtf6aR2r1ulDUIRtklKKYG5
Av7etthUxUaCmdXduF4x4En5qNVRAvf+F0buAeZfzvrPWcCaMIt3wg+Osgxkjt1cBmmds2K8DHQ8
m6awDtx+Y8LCDqXyxhaP3cwSHh5h2wDREuVR1neggMEmUbEhfLgU8kh2EyZasY3ZjZ6QHZ7swgdG
2q9oJnBrzUXYbTkAM7/ttbLmh/LbmDR+2/92/8dPuW/UNY89/BsagJoRe4e6+SGxYWZxgR2wa3Hm
EKXm9p2HV7QjVRxLLhuSw+ArSEFsYhPPuYePrDjtaYYfc/cR7TtZ0c7vrsNAG3T7qTPVzPQi6fGE
jTKpo++aAq46DneN0bDekR/MDP7eFSSIld3Vjuiws65aucuHdSONNYpBqOPTk2xQOrY4ciYyH7WA
+ycKv4VmgsHS3l5MRG9gV2o30GIDHjp9LnOn6CTK1ENWvnERhp/x9q5aoh8o+/SNVMpRZh/StnFn
/OYOMtlwqWycn6KgvRUUk0AL2FYQeNiCpQFc5DvQgVGImF6YvXoVIcmbsblIY6B0BICOzMREdJo1
ijhmsXjA3tsucdo9nE2gDUb5Pq9xhTaWZJbWLvzmui9gGU6uA3Wscmf024BCb4OhyC4MacolGk0E
C6aLpdiSUmNIwkzjDKq1hI9UMxh60WSGTiXCAD1OEN7BYip6021FNtytWZYVBhtr40F6ZQcCS5c+
wy4ctB+kyFp1eZS3OJ+wuYgeYQEc/RgC8Z2FonCJugmW720JZR0vJ8N7b/vLbZKemIgAMYi1YsEE
DU7wAdF/mh/b2ZHDJY12f7m+LJOJV9OXAT+VwK/aeKknrQHYe1eNtXMVyEXecEH5uGcCBAOS6rNR
w5gfB6Dw6dkMQtYc4D5NZuP79DBFA6ZsewUIJnV+4LhQu6RvFZ++/t4KjMoB2HbvLZJ/BVcrMijt
blJCrMRfFZ7tCDYR47lgr8qJ4o6ywbldgaJ4bCFRB8HMi8d+25Z/VQTg5NSquh2Q04zljexAiHn2
8Hga1aHqzZKCJAgfbMXCL6dC23elGA+270zWQ+CxYh6tFdA3vvq/Fm5iVSfJAEZiNkaxp8saP7wm
wW/fJxs9K6B3ARXBDU2jud1hUenlMVqVkoWJQgTIvDuCqklnb3z3Frds3T6L4oTGBLePmlqax4AY
4OlxAYPPm1NuIo6tvEQHAbYRcu0LGuX5IiyJdHAGpardinPsDJK7slcqp88ghQvHz/g0wTj9QD3K
oTEtqdLaZAIYgR6WiSV02hFblYlTr9EzXVa4ddiKU0VWPMVgRCO7DzZYps1nNDI7XbzkAO32zMKS
AMWdXMXFpSkzWZdor2DKxDAPs5FJY506MZiCFKXC+SNtpwNRzNHwKtGPskXyuTkNXnT/CariYn90
xeYSEH5F1Tg+G8S+BTe5WyPOW/KVpt8s2KAy65VUABX9DhCT4pZxzaX09B8lG6G16yaEPbUa1zpP
tAjHtsmGpld96YkfaP5SIzmKwSZ+RjFZd3CFZXs8rC0aaA9EHurJAw5G541swlNDKHQQyBWtPnoF
N/20zKhKjq6fUDjxiv8GgxKcSv2bo72gFYYt3LfVVf+sPFuRqweOH5JE20nAOXhy1If0Yn8kM5vF
IYCxZMoTUX3/fw6ND7bE0uSELWFyQc3l0xp8cB+Jo63o3K4CZZK9oo4erTxdjSm+twlYhrjB1PR2
LmBdjaMkCuAScETPkDDvjIL6ALGXq0rUGGAOxIRYbcfQgXBsLfqJIk6N2TcjxUFePJR55vZpS+Ix
IKhjtyjUcMa0fRpKnU7/fQ2Oi+YFGMZagzCqREs0+kyd4voBuJb11rbbLAHB4UuNdg2RhARiiM4M
ordC/lRTxfUdIHbD5ItE4/SYvmzf0XIUyE3OvJqejOxP5DjHvVJcZunTtiG+UIMWsno5Ml0FtkHg
18IEiqLRECJQbGy7YMmrgsIWb804YRIcUdXKaTQ10D3dgzvpY0ZShmEhwTYp3LiwkrRsZ3IX4+PR
ySwspaaW0OYPaQtxLp+Zw+LtM5vJenWEszSF0yc1JUK6RLpw+SU/l2VZ2kyCuqePeq6FsXvR5jC5
20uohBKfJs66x4Mt/neu+zSN9ZvlX4JQf0fg44Js7A1Yhw6Sj1AlOOE+qnvQDux8E7afJMsCZoaN
TeFMBmhCQux1e7steXOLCW569HJZbS2JYdwlbF8gKp9CEN8EuWCE1WIEm1Li/DaLGEVhDaZs6Rv/
ygJ7Sa7kBgj26P83ToblmIyKfWiZMj5G5NzfPCHk91DdqOcfClWLKum9LglKVb0j+yTVdgO2/YGH
/3KARbLl4E4cHDSlI1R/LeDvTDWPMQu96esSx/f5YDc83+ehazAxlGWWyj5DiaFjRwBVIXlu2vnm
wBC24Z6+0MH5a8txc9w0Ijm+c/kGFN/OjRa5/5QEf3tEglZ7j7zbVHdM1snYqYfR2v4o+NqF/rJR
NRwav75tEWe58WzIUPw/XzPCoybSA3mYxpfIBtYfJvZhtTs+8ApWpIr5s+mELP/lz3iop8UUGCjZ
4lq4BVonkLnmJSxNukpju0lNzyaWDqv7H20hq3wedEWxanDNpFLmao16kmokUJDAM2cwkpGKuLil
2Z+c5Amei3J/jQUft+v/zb98UMEgJ7TMZZH6nJsH5U4mW9Yyinq0McNkj47HtoY/2amQsrnEIq+J
wBFfWR+e3/GtyxM47PdvHjTMDZluU3wYVienFfg0yhMzxSraa0GoZO0flbHLstksrBy+1sjItBmR
b1GTPnt/L58CDhMiSPFq/TM2yf425ixGj8n9giFP/LqRXhEcLdX1p7NWW5ccaQHMDODQHdo2rF9e
SBReJQVnNKRifv4aqm0ErlqHUIE0VBNVuwBhofE/vTn2brjcB/StrOf4Asus0QkG3/o7eiCycdaB
ZYldmNsV65BClkJMGHJCLgBJzN2NmjQlK1t8sJ2bTzm3AWGAWDumn8jVpFZ0G+hC2mUPio3+2eBk
SLPLAtPghrIHAkDvQ61AukT6e2azqH+t5kyxqv4IdaYD1c8ya/SiDcWAOgo/KVhR0FaRQFupDVDK
ROq+HSAa+XBYQJ7/KlmuTsQyn3e3gIhIQw5XI3K4DPUo9jCoLcCRCrqbrDfXfhvO+AhZzwHSIQ+K
VIL4YcS+VheDYNkoU49Wjdb7BQZnjEtvWGyuE1Np7/dAkCVFSGUkH/XyJTTW7Lu32xsb8yPT9Ykw
66kTiNxVaGoV8bpId9bVacSTaaIJn6KEgWbCDlVu8nsor25vq/wXyIpM9GqTi53uTq74ADvvzl2S
PTmmDI1ZQ4YqUvOqwBiWPjpy81Is10yoRwro9BjhqqkmXZ34qH09DqhrvtE8vkvjb7Q7nWV83fx3
qJaR8b96xi8aPCsoFEfA80CLm2W1Z9QQ+ASrdB25YINgadl/FDDCKQSYkRfGck+qd+gx5WxncNS2
K6cOgTCgA/UfRp3DglUOybpFkxYa2Yq5q4M6IfdaxfejBfoqcMa4JYth3KWrJeO0BecE+7zIzpaV
AiSH66ewkzqyD+CJK7vWIkBbqTZ2tvc/2NkSxM4xfCyQUDE22g3D9Nsrspbua1DyK0JTS4nJCUJs
lXzBDx0xt+85NyvVGtz661o2EZrneStliXNTUf0SaCbT8riTkQfmY/teZ4Hcd1NJB3UMYCvPsQFf
nO1VLHxUhw+b5BamtyCu0cZyfdewDMqAQNPF9q//uMp85y9hCjNQNPpKfDL3Dt1Xaq3gWW5TP/T5
C1wDIwXvPcG87ADai5m7PP6jAFoXdGId3yDP9jRb0NHK2/AfT03DrIV8xDUGhdPgyoizyE9yzlmS
qKVOB9tJDe6BUBn4on9QWRqT0GCdVe9UP4LkKEjbsCha1ZFDBZgNKxlPjq8pxD4eIW1loGt2DBVr
tia8YA1XVzGCb2jU/mYC/azabnhO/arYfA7bLjrckuJ6GkZ8LWeizdGebESoQTDmMMfk17EJD6pH
45cHH/T5lO9BzpWVsuNgPyE9f0k3Vuol2yUgWYAc5ZXPr6lu3tXCTr2AL5Fmo9kpblWJ0aqTarmG
QRx2QuJxpAof+p1/Rn4hEPdRTmDfOcdDwaQ+XcSMfPXPtztHD1y+J/vhDIRpPPl4EuJwJCEMhdM4
Fz9rxxHU8LY3gbfoNJtd9M1AWrxUP/xqdwF1IMj31NoOC8SacJ3nJyhlfnrM8Fp9iyLYsA0DsiXj
/k3XZLHLzF92belLFUBlAl2SKsjkKNaNrb6MkZnPWM1A7ucwId8wjyaXSwTLM15ZaZpF6OWzWhCY
C7nujNCF6Lel3hWf5jMbtH9KwaRoJfBoB3KZehiYenYuvlzo9STueNiRJBpKjHnEy4dJ8tQutKeN
WROVgcqIxnZg7sz6Q4MwsHTgn5/9YrsXS4QyXA/Z/dEyRnvGdzBxvA8e/9z5Vr7yai0vySyuLB2Z
PbuPzw8BNtUBWfpS8oAnN2dE3g+wb0lgYAqcRLveLFEeqfS/3qkq7Y6+gMSe3Q0Jy7Z+LvJt9jS+
b+Z5p9SHoGgYb0BbRxWLCCuGmmgyJTaRgvzBjs+gjeQjLeqLbbz8nsMHJ2bHQQyzE2LQrgFXSt7v
GROCAy/vaCohjM8Puc+Jz6uIlohrUugSoEjvEgiobGUm6RH68ibFQ9rgEqKJ3HrY7SmxUKAXvQk7
e8ruKWXsIBcAxO99+pcqCNgTH+MF79Mz6YR0dwsI+T5TfnjFHCtsoGj5QSj2XkrtP0Q432bi/N9t
gxGTsgG2FauJku9XznNj3vIudvPCegt6dJGkiRJHn/elrT87bAFWMxvZjO7SvnafQPB3dMEbBCTP
MpoJXXI6QBneChbwqnVHvAMBvhrFODEEoVdgcsnaifcUTXGhharijfRNA3H5ByD6wOpWlgC6LyyU
0ls2uD5Jp3Cev0LFfSn7nZEaE4VNs5GKBPSG++tGvjxNpct6+YS2yDM/y4/I7DJmAiCr5O+GxF4t
M+oXVDwIKUqiF1lN0YFPCdxt0KVhi5wH79ZTYeBkF871D87HBCiN7kYoR5BF1hrGE/+4wTeMasdt
BNtLt9orezUGh8Im0I/LBwDGPA4/HxTyuR1mREx65UqFI/bLGZPMehvkLsNlTXXmwWQ0uaU7a8H4
8uof4ExjMjGz4UyOw5SUMq4SSozvQPvmpmYSJ4kLdl60v0cIXpcXAzGHxOpxBWu0p3ylod1BX0Aq
3113qJLagpfdyRFMVJImTTns7XmQKxt+fGeneISHL/Hs7zDhdOxpSZw6tOx6pmBWa1C+zksf3tGQ
xyX3+x4evCrQbPOgHv6EVt/Hit0lLVzFAzj/PoJH+qOafVhRJCdH3cZwJOnV1bvBgbFikc97a+O9
0/wi/OFvxQGieYAXEyPHgspPBsvvMmeTlz4FNI5Ra4KlPT2923hZgPSFw2JmD+gJd4xaSfKD2bQj
Dwa8kka363TecW6Msw5SdwvSFHXryMBj0xKQGO0/wGqHQoWMvYKOiMlF/48/x3I0T7fTPEs+sYDm
4TxEo+gjl1wKIpVOSuqMXkywSbNqxWM05csgOAchc3c1afHYOkOwYp/QXjXwBhoKY408hRkYmNmZ
6a498+pG2qUQsxuhEyQI6KjSMpM+5imjmJHlYahKLbQMNp4gL2VUrDPrMUjOK0kW54MMcRcGZ7yW
5T987OmD4LBhmlWRUFfYuU2FHcIUV7e/UzIT6zyteS4T6u1Q/OQFQVkBgRSTtIVKhTXCYUF77MBo
G1m7trS5TSfuzetsGI+X9uqjEwjfr3z4uDL8FBd5fTZkS9KpHqJrUxtImqrqpb+KjYoZj7r2AiEg
ByB2raXEmEgUIdbsj4UsG/NwgfLBl5gx8pdOZ2sgpnMZIORUJhMkFXb+fAc6DrnryLsbDF49Q7Pl
KcOgWDK2bG09TLZYlISQVULNS3Nq1fWvfMqLq5m+6GB7cAyxszTjwzZN3GidIcpw5rNk8ugVwuhL
VzR6i3o17y2goTaY6bJnWcsgZ3m2ZyJHJs+jfB588iru6bkGcQ5l/FM2jBkmOn7BfNJmnXVZLe20
PvKIQh2aKK/RDMtYYXPJUvm/pSj0zOgEuoWsDO6MYBbyDTgfcdJMa1Rh2RZueIyKySj0U/eOzZvW
BIIoSz8ILuvsp5nOHlEl5UbNiQz2aiPjwSOmmrYNkPv4qvYA7WBLuxQpMK2KkH7m7vnt4aF/xKgK
LkYfxjarVNiNSwe+ZygvGKc7+PXaRD0XGD/Uhm9ao4n6hI3vQe0uAlAjepeYCdEaajypPm5dzssB
QlFq4s/dETVdyfkGULvlnak3Z9+u6Asm37loj0DL5Hz1hU16RDL6OOFfwDIM/UXPnd75qiMC8UU+
e95p8NHr48l7e/qOt2vqQ1cfpUJwqnOXWE981DSp08hkfJNiyC3HyKpzLt5kuJeqb+SKw4OKipbd
++dYbCWL4izCZu9qX/QLy/MTRtuCV9rfhoJ/fb0JM+/6P9rdYmXKTWDCbbopspDlLBIeYkD69qPU
ioID3RZ9qN7Z4KUQVMidQrjvV4gtRRjGGtaUvmYB6jkTQwWD67eWhvJaf31mDg8vmK6q+cmlz8sb
CrnzDniWJQblSxja9BMQWii+a0KlRYZVfRDlgcCMKX0mKWLiqv8ovcm8h5nssPNtjJEwkGjXaJUK
D1z2IqcQXYuHssYbZhK3CGl51zxYSWlzonh6wO3c9SJErolOEi1swZuiHTRZiyE/lSAtTMCb+fAr
4yysJp3P6vlitVTn5HA3Fw2P03IZRoyqdaNmb4WtNhIrvzhnJYwyg1v5fSumx8/d88wiv0VUN8UU
N62BD3qmDhWAPLYAyzjmhCkbyK0UvI/04EDikvzdqIArYqYbB/ibopVh5Yigd7B6ynHXuVyaa2kC
Sh54OpuOkNKIgUunKNrSmOMw+NpGPv4kN7/UMc9ezeEVK1aKreDMknATQfyocQSHfhweHmYJUAvR
W7yYR5DrO9b/2i50Wag1fZMle7slnlkbrngq/CEjLd57gjKubdXcI3Tohqqwp09EbovXW9lgsoW/
D9Ka+QCGGzhEGqq543s5uCnS8yxbv0qIgzFAvl/07AlEv0V43rWImo7d9uCu7EogG8hdhrtPe2jh
T/PBeeJvYAsoAxrgqF9HN4Ca4LQkYM9uI75clyn0UU/z2IEIoDZOFOhJnJOZyaC6fLmMU6L1KfYw
7sqFupjKe27vbSnZxz18yyug8z5zOJHci7Y0kHqMm/dN//y4KrnkcUSqubsoLrR6mqs1asyf8Eim
r/K6ueubZCVnYAsU/IadYxEo37joRKmbB93alf1wo18Sw/s9emfVr/uN7QozKwt4v+l6HNhb0yPe
Nx08Pnkp4i5VoM0uXBX5xFFY7DIOcV/hCDG/P13gng8/Frgqcpv8KiZvUhiFZkkdqW0BEhbElkPW
k22ZeCZLQQt/SjSlqNmqK7ZIe8lFNjFGtWCAEqjVnYt7Xm7TfSez24KFN0/QLfCBXiMfQeZUc1vC
ppxFZVDG2matVnX9bkF2d8gsoBk89iV/fOWVxNZGpvVq2DWAmGOGH3vZy06/RNLOz2hy+8xrW8Hc
1igICH+r3gIGyjcwJMTEMKERWcuwBJYviRUNZrrKbjy9qSk/wElA/EpgVz0LsEv/zb+SHw6KdiSy
AlZ/nLbd/pnBh2aXl2jxg5y3RmotPJjBDdOGQj16XzNV9OdEVgmLRJaf8tUjb1Dh9G7sjm3Nb5vy
YOx1JJd980zDOG6ip+SWzb3KWMXGdQQq7H4Gagh9oCVJqJLxizapbOg1QkmqY/viy9If4+EALJTn
Y1ZC/NSsVsWURe1H558jQwYi8sqdRrcEg8blPTD7sMrJPSMPBA4wOIxeV2PILWp5QmpmApVs1MZm
WJpXFCbBIuwz0ZVXcM4Z51Qy/wc1ydkKQesvOw6cwNwW8LQeDrSFCP6VM8GVFN1frECWj4FsKosv
ir/I6iu+Zy5Jz4XmC2d6ELbq3phizmEjnC60K0mJK81ErQqpLWi/HjNbx/X3HJdxpnokDwY68tz8
rANJ1Aq/2pEzT73u3rlsLKT3yY6fxq3/AuwhrUJbeUDuEE7bYs4P7sk5BM3hkruc+1H2ibYvG5Nj
nRUB5zm92hyfKJ5Mkv/ujQWN5me2IXucvUizziJ8gcOwQcPDKCgsanYnpjQ0tR3Sz4JU9R2co9ae
+XkwyVpeu2zrBjvh/dC7+lsqncUZptmImsV03zcAN4Wx6SBCjh32oBwwJzTCrJoHNfRF7Ih7dIY3
/FP0KTVIgj+qKWE+AvefgpCHClnz+puTEKu+bCvU0VzGVE9YNRU/V4YGt9JvsyWNWpg9nEhoLtMX
LBWGee8LtMGA0WSGmG5jMeLdLfZrVGKzOTO2bJ5LjPprSczrH5SwgU/o/CL2mVbQ9ilWh1qgbzrA
JJLlo8vIX6JGf54vOSre9jfgnzIrR1TCkYF2omsYM1CpHRDlCymOQsfT/S3F/WZwucw7a3MmIE2j
jA6zMqeSwe13wggeA5I+ksBNKj5hMBXhpNekv0t7Bgj5bof/liEdlYYe754DZ+fdUxSNZHb5JzPI
Qx/vzej80wOi5N1yF2HvB3Bx2qm1IpaLLfu+Q6PPBxVqzh/J9TOupfKGmODFwY5wy2/S7I8JJoRE
otjhzioP8rtIvmUCd3v7EO7rdw20JKbdz6dmmbtAnBZdxANZbZLYvHN9OPu+w0PtDPceI5QL8qDg
GYOd7E63CYCKK/EN+eFajo5IpigSa6n+ezOvuWAx7Ls8WsV9mWyji1Pyi30sttWqUvHZyZzarQlw
4eRKqlRyx76t0bBpJjK7Qa9PmCkHztQ4mYr9Rd4xU00zgd4gX9JjtLXoXRgBXnVcnwtu5NJWIXzA
Q6b0+gB56PSHw5vmjz505GZMAjJjJruQ8avB20e2NLyle2M4unOhVDUvwn2uHztqXqgil+1+it1X
PjCjVaw/bjelYPl5zMykeKnO34NXEyvMapAGNXUnteHqG6OqBgnpYpW2tQwAeTNE9oBYIO1ZVm/P
aBDyGWyyQNAf5pFSunpmoKjAivCfemfmAWNMs+LTbJq+sZyvK/8qwvswG2TGsWrvJH6L7LG6jrUF
HXUOimGOiOLg37k8hPMUXL+wr6THWrxbZd8gomqlP1H0GNyedHkMTBNYcLUHf3UX1qB1y1eOvnTR
gx3R6XQx57/uN9ZBZcjmJ+94slzQvRhH4vaq2HTh0T3cTA/eYXQOHDlx1fbjeL+8nLoen53vgvKu
CRHaoxBa3r3KBTayCiDquBQgcWcb0S6pJjCatoXyi4lJL8LvZSHDvD4MbuHkP/aqrv1dxX+gEIGG
Yo/wpbvDuFxFxsE8eQ1UeNB6ZXOyTH7lfPzGNdTIkKZ1sya1Bu8R/k19cf2qm8523Qam8it7I/Fx
PzGPEcvjT+7A+KKey6SrNvlAYCnqjN+L6Cv4R37bClIMd/wWXHyCJyKDEsTGO6RQW+dxdC738JKd
jVyUFpLjCbuNSMvCDDSNgheXrEyu7/vLetU/o9fbQP4L1cAa6ErFfqOUtqp0FyxdRIs2nISW7VIx
zTDiFVqo/12teIpAbSoa4EAuTMZV6J1egAzbIZB+4q8RpPPKVhdccdlwS6Ji1Cdjae2UswPjrvGq
e47QyOiioOR45npwWJ4hSAsjX+sZrnYFTc56VVUg0eVCAQUS+Y1bG4AzPbNZL+B+iz7lotbNcvLA
uA6Qbjh4zwpnSlzSVSc4naOJLJmKjyUWpHBAWjOw/PU0rH+bHl0XGYR+mjzWmrBMXgeeyefei+i9
H3nLy61c00JxMWffev6ofeju3HXll183eEKfPXDGCiOrKytqTHlGNd9UEB7azuOoHnp64VMttFru
+hGmE9TU0hxpXzN1SCm9TkUj9TScZ5+H6AgZ799w5Gv/XgescJI4RynftBVc+1FWm0nLOlp96KAe
9NUyrS/JAhk7KCdm7nNDzrWZJtX+lXxmQAdHnP0kgtahq2Y+6TAmbEzq9QB39vNiUX7pGEiZF4a6
VTQGH/7woQRnzEydMrh33ceKfHH75c+SNYWVBgcYFAwGPn/t1Er0U2aZ1ZfPASWok1GLplXdfvw4
q95n3Fp6hVZvVf8Z3JtsH9XpHdkqYDZCUohJCVU/JHD7L67t7TUxnH85rDVIAfpOn2/YTU90eCJf
YkJwKuFSgT42S5S0TUII4I4Qkv5lcbkN0RUEoSMU9y4IhENgfGhCLh2rkC8gkcX69eHe+DCNE1Fp
BPTBPNrR0D35XvyoS2eaVjHUZ3wRtbtIcTHVGmp2G44NQRPNT6FM42Aj7YQyzKG9EAfb2uvFmqTc
unjNGuejLL/rUUIXek3/BxWOpD9kMBErI561HjH65xy+OxbZuKqxA6lENxAtb1019yWw8P/VWdJX
j/17FNts4CyLFeiPB5itfzjti/PJrjmfUryfpodpwhFGPl+prC3dg7AijhXNezZyiIHDNQhHtAad
GBf0roK41cMxQhMWJ3xyV6aqhBrWiZcu1ZBukB7Z+GD9iundulJ1tu9tsQ6YTRvoWf4NCrb+0bmD
wRAJAnNpSp528fMFVJ6lD+xnrPEERZ+hI7MzZqWnGGxUHFKgFseoblq7+XNau8cni0fz7PlwU4x2
dBLv4TBI3ksbv7YV5QWQ9WJPE+FNmqMeyt8XpOKL3pX2BR1cR2z6WqnMQxIrolifQRDbIePaXgkL
ZZa2sYsUjDtJZebyarbUUuMEOSjXE7xbwFLSJ8fva8PerXVy64E8KT3b+w5268nj8Tf8bhquQQmQ
JZYl0LZLJb2IGBMm+r05b8WLKBgZJO72qaJJFvj5FKM36wf/oPC6fkpkPKwlc1fN1I37ZeofWt5w
MXzLDL+2MZeDZ9NtLf0dKfSo791qL9+wm/16COHDhF9Qsp+DENLVzviYaqswBRgLUcrpJs9t7S9v
WZyA+f/AT6pUoeIWwYN6O1JdzgHE16r58Lp0OisWpuOOolgy1sjwEd135wAC7iFYSmQq6f/UwohV
tufwXCx/NmOhvtb0YHn+DI3nn0f0mTcsk1H1ZRJWX5WUKmKxDkyARTsTnKqbcrIkj2AIs28e+Qu5
VqU6D/0fHIa0Mx3nppVcTVsHgMtC9y4/pIMTBGxGDLwfTzdcxnojTZq3MrycXaQDAmsp0Vi9YpOi
FuWS5Adc4E4BkVgQfCK0MFz3FZ8QSoCCdznhf2+T2UBQmwSu028tiglGClsOfKmGTYeVXOc0/Ru1
uhB/UqhT6jvB1Zdr1IbOw6SGIrwln8PAtzDweOjtp5QxyjC08PxPXXx3qHKzlQ5kZCBJj8UdacxI
2eXSiMs3xBJOAXz9HgP/lBxiwKHexAEdqguFA1dFSSXronl3uGxm0ix+Yd2DP/YtmilV6MNg+n44
8EraaMFJKQ0Gdd6abUuobHByB6lXX7HIOd3qT5N+Z1hA5CQuEz5YPIHMjKFI94myTVrqj0+9myQo
FRGMPbXArAhEhF3wWsZlCMch/noSWnzyX5sK1AKzdLzMYxKspxq6VwZBTrqXpGqQ65BOXA93gpSW
jCxM7xsnl4oVD2+TYWGhSOmyVnPUMixDWQ3GhyJ7GEYc81Uh4msOqweoPv8VvjWuTt56JH7+jOAl
B69UrfyAHlkZSNu1FEDXvIpqwHlqsaInjpx/2BKMTxR+1zteZvneuOm6Nx7Gkq0Uf0wArH2lh1O1
ZWbddDrBWij3NxqIfHAzdVH9iB94nCRIiGgXs7Gaosp2+/5xmS/eyIRQ1hlHFc4m7kfd9fGOnP2S
+BO1iadjwBkwSHkiC17Bd1XN6eE3nCJZ8IjS4QVkB9DK4IbB3kfni+NzX34mR3BT/VkmbQU6nFAA
lf+TXCHp0LXsAGSHpi5M4bbciSBYPbqUesbTQKtAJEQoUHpYvLNjWEbCqwGEdKTNr8drd+uoc3m2
4/p3BY9iOlthRiZ4RTuR0ykxNvOlNIycEwVO9hGu7QjcidXfvDC8t+WSqxPAjhI0E33xx766dncz
If+2rHWkxG3f0ORy2FXdDTZEP20Yj5Oz0oSOFAN9P5SpcK0hjTn9Pep1BoYjE/ZoxQsRqaeVir+V
6BFTGugne3ADnNcEknscqJjQ9vqrx6kDNznDJEOPZweDfv5QA4NVuYuBDWo3YGU5H6WkyR6KqxKd
sWFOa7mPNBLnmQIKJo0PIXdjNphM5ZRBJ2pXH4CQ7MhPyUB8BLgbT/1IAvTbZQvYKHelg1ZcHNwd
9JqQv16X6zX8onv36hOhXscNh5SsRwyQjCIRBbBFZleccxHrSWzi21QyiRhLisBdyK8fvs/nbwl9
AbjpdlAFDX3ap9GaD1/0ZOoc+t+QbkgbhLuhhOr91K02zry8+HbybMqmhbOL5zOnsowWP16YZE9E
7cYHlN43FGHuXrto8xyRT/mCOmjLAqCRrdtlskhdkaabrLB3cUlKys1OhKjgXSdsWY6TARd7JP79
6CE+vzIVhWXSbozZeIBoixhbbzwlhWvfQt2iCm41A9xRRTxQnCRXj1lAJuolRmHZiiT3dJVyJopt
yaZ80sr56o27/P1ngwbNBFbsqCbbHe2zFGwm5GtH4d4+Iko32xdvnMjseE+whNUqj1EW542Ep87E
PRwgCfpGDDKELXAsRs9X016J1DO+DCMJYR312owIVxl3NQ6CHyeXEndcxznEJ3cSAcO43GZc+3ZP
CtWOSJr+fmulX2n0IGjaapXxbo0LTMMflzQSn6C06fJeUkBJGjCgO1bEJLVc5c/Mb9QfI56NFEde
xH6Nr8o+bDZloNjWyZDSeHS3pTZwHQgxZDdFLjCq/F5x5x7oiA0CPP7/HZz/n6TlHjoLPNQBa8rF
DS3Ue5tGfPF6sjQxa46d7wdpqlOxlmulHfi5QyPzFE4xnwJ5GUyMtkyPdh0y48GWbI+Y2pOrqIVL
/0HwyrB3s+SmgQ8K8fARz0tsSXFUwmx4vwCzuIJYpHXwM+itfT5nP5lY90AL7r52OlUmrrsDZJNl
I4PnNVBx2Yii6kKJJb6GVPdsqNWbfrsy8xcHPasY1yL+57kDPRcpVOIfIOB3fN8YXa2UWAqowS6Z
G428KrcYenHmzou52MpCd/My8I5E+hju+8oe5qjwliz2fjthU5cT/rRal+GFKnMra6cxY8c9JCex
+t+dBJbAB3QXefsu54tgSd6C1YyJJiYCmwmwF703JNNcVf9APXoV2jFqqRSR0edCKKJZ2IOB9O9Z
5Wh7lwKUDn4IckvNWerPJgH2wBWnb0UAwwql17MYU/gcH1DXEA1qtJvQYaWpe3Q4yk6ZVzBuxdFg
m+0XKUrdkEbTh8d/iKCF8l6W+PwYUftHPViQh5DPtitsTGsGGtxAV1yEWAtmJmEdHQSAT/T+GPWh
l2Agkt9UX+oK/JKhQJs0hjmyVhmIxbGdFzr+UEVnsXgAzCz4RBF8oXLQSEzlEPr/UTUlOHGReJHc
ofTsuGyXCZwXCq3fQCXIYwcTD0TECgGMI8RjnthBIqKLeA8kD0VetemMx6uqNzVFfBSnzr+zPivr
+3P7sVkPXv1lXFRaKli9F5Wq8EArHq6a+fHyJJD52dfB2T9qTCDprcjhZGPhO6XvhEqXQW1NavFz
KGWIBHJk6TNlUBziqx5n6ai/llQhOMVao9ECgEYCocRX6a98/2yZBV7L1q1e3xWYBFoA3V/6vp1g
tRIQy6YzUDuAwXvs9U1UwJANuxwzTnw80oL5o0TCoAiN7C4K2vMFOGf4/d4U4mgeGrDyk3MXGzeH
uyr9m9ou//nyKmGHXWeJDVEr50xG4KU6cGyygkOvluj30ItxUIAJnDetBX1bxq+mYFvAsQtIJM4n
6SfEjzxashFumWhpOLEZ7PXXZ8moSYLccqistY9ZaaBta4WGXdQRFIJd7G838SHEU1ILFk81fA32
ZK2M7wFtA9VXp+z/a1FY0kKK8PMbJbOXVxmolwr5PtW9wRmRLdXZ9nhETwznM4NJLP/a7Gkvv0ve
hSGE10e2MOA9XUr4017HQWKFmO5YwC6ep9q2wKGaOFm8+i2f7gROXYE4+hXym7bBIgK8kPSMHqT3
dSTJvt6TLmK/dT/Y4cQVJ7pIgej1BgzWdTjbwL5FkXj3I9KIHhLM+S3uLQugyN0lpNwVJln+bD5O
LeptLodn/WTSbx1zrHtGAauuhmVee39Q7MhrsCTpeXXcQQEStJYpPswU/k6JgYRY3oQgRh48d9nt
mmykM3ob0MRBt8Yg6CQdw5nvn5jjtQfG/GZC4d5PBAtf2suVHo8v7WZV9nM8Rg5kqnzm8mMKphhf
lzymod9SPythnUQA3uUl5X8YU/+RR/VBBQehrq68eKXd8vdDVfGILKju6djnpXJppB4vbsGyawHA
vh5unjjFEVZEPxlUmGTUCWczJaYlJZRL/YD3L/VPqqzy5CEaJGuuGej04pMa1YzXHua9C4vDLlPd
XY5Q12+Lvyh3hfgdOwlErpB45QiRfXlqEVsyAp1E3Iu6yGDZ06lLt1RhtLWYCUarpgSxdzmjaYLf
fO6usWAuF6sHlRLhD/BRdIa/SGn1hjGL9Vyua9bQoWsha7zqaU7hKX4f2fYFTFvi6Dn8zd/gygYI
G6RJWYtEwSWSEWwfiufBsjpi7dvPWeqSRIgyoAdzr4+WWPo7UJIpT+5ujo4dxUAkqd9xOD6aRHjQ
FsFJhrrQiR9j+P55uRxmN3PjybbAMR8yfTr26tBcGpK2G0HTF51f5pZA14/oLvQi9WM0i/em37eB
0UbaULl6ti2QC04CwLjApveHPqNvX0pUlc/T4s1ih6tD/FwC6cldieY0Wr47+eB6dkeik3FEDbGj
oux+n0g/fuNpHO2e6Ov1OzYFU1SVY2ZZG0b7RNOfRM1ExWRyRUQOaJSse6e4+pAu0lKiwdwdO/5U
W4Om1KCClR6eBO8y1qB4KkvCWBFhIsgJ6Ctl3BXyMpCxnlvMEKjo9uIkdcP2y8SmCP19bcZ8o5wy
IuRwQufUfXt4Aw7B1G/lEliczJogVqptb9MUMVwuzNc0b06oAQqY2kdqAWXJOVgu3CgZYe4XApon
tAivFMHJP/E7yO6R17fe2feaQPqSfIXin5/nHqX8LWXEvEZh5C+rtEpdaz26B1yKiOzjfRNzV+64
RehRpfVjrrBhxwhdln5vG5cgj/Q1A5raWWxQ9ucZ8f4a51oEs7XQuBLe6Yo++YR9Phf946XG0zsc
iEvpLkSp6rjpPHmtxkdKDrxZAK63p1MAAKdLGI4ivxbqn2kNGmU2ayArQaHrMawrrkTWlI/uorfi
t/OQdW69q6sjGSOif5X4nqYfpdHkSXzZ4TgnN/c7R0Fdb5ryFjMVTJ8OsgRLQ+pXGfUvChYMRDxQ
E8/+RWKEaH80zmBMiwVQlGstaW1TdXlpN7Qn2VdUzZ3mKkScm21PnBsVfJJHV7q5JaoGebsEER4P
X5pdYI9ybeqR/V8494PYI1HQ77MhdByIr7BnnJIw0osDBz0iSW1NauPNBSWq4kyUfotjLFWbVJSS
L7VVSJbSKnN7VTLwoawUwkdhJEjA/aPEK24N9Oc2+8Dz93CGcq4sqkcQvdflSTfZYY6ydRRb6NyV
REwjwhwaqjERGjSJtQmMrXONWEeCxxaRZwhppoj0hzK3kITx20I3MmM04Su3mnTtxHCximX5b0fC
xOwo9tIC46BVdIV56nrtWD5MYs3n4mmzgr26k6EnVTVJ0pMZK82cs/5Ug7hq+07CMi14lpxoqUDl
oleAa61+oB9LzVI+v9kKMH0MPLFb+A6ZfjOOWeJKNKyfbD8ztu87kPawURC1wzj3j1XZQE5Tui7q
9q25YXMMNx6jdsO7oq4CNSXfWyvN5tqILg90uFwVlQozCMrLeV2GSaS+0J3PGemqTZ7rNgBt4RQ6
xeXdcD3mOUYsXZOKOW59ulxVCeyf9BYkDlZx1sKPy6KZVdscNMBPWa9huR0I03IxEXQmoSDuI7ke
Q0AHUKBKUZzCiDCiTyYPec/CNnzpnLujOl2Agray6SnuA+rW1r0koHtCcQtQ9h1CGbSnN743i3fm
wS2NxpAw9bR/+NbY8oOidNQEVVbqcNaugcgmDqe22mEiSvFK8LSL/T5J7B5MhhGUjezbQfkHyIpb
NYUbcVoASHiolPf6lsZa5GoR/N6tJjKIDu+/mh/t30JvJjK5NeNyspVOl95tcqHSrt8eDZwvyLwf
EqXLdl8oOY5ERIybF5272pc/+TtqNo0xLCmTsNOJVMxFw1eRLVFUxtKbC1ByDTkGxrv5MO4g2q2b
LdC4qvX4/FLHZ/VAA8AU+IQ5a52MnD++FTVnVE33PmRvjDqhG53/s67jKV7bzTOuBnXi5C/OoYTe
tTzkFbfNCQgKifOe4IHwpvWCiCllY22KefPbSGMRhcu4K36+dkZKVaapJfMirkmZ7LzsE37dbTmK
eEXQy1NIpiw6LUvK6i3wg9uE45foM4EIFsqeK+yeju3ucKVp/tXuhh1jLhQRd/yRNuE7yQ0wn6Ma
h1y3Embzeq84Ur9CTvniAF/+8oD1u0uDpu1HNiV2JJRZkORBztv5GuN7/UAOVvT83SEuzqlGqnHw
pRFHZJPC+dOjpGUH+GdcUkwPA7AVYOBf2ps57/4Jgq8rRG26vP8HgdLjeo8+5YatleWIB2nPOmTw
iwIJfmnbWl1oIWxpoJ/mmjo4qi3YdMGmRs/p+tW32Pne+6lI1Pi4C0BdGXvP0WWD08gpPbtJzsfr
82ezcsnpKEvtAIuH94Pc7k6JdGnl5UyAASSrzi9+yOThHKLZHE/t+B+QbVucS5Men5XrzTu+FQ5p
wTfQnJJvB6GNTE2KpCgtPko7/+2xavZiXzI9rQ8YDt6qzGCNATcUhtKQrcwp50xvaUR5og0zhUh9
dRbnHnThdiQMx4CmfNkRGjVNmJrT0rTpEeAJB+U13dtMtXUmbX1DPrdEVDY2l8JQxGEw3mn8PqBD
hiZs3Ga6Kpobs7uy7ON1NLNgbG8tUS1tF0fps6M+kouCC8taZhBks18mhKYvdBaZc/+q1UpVIyCK
e0ouVTCK6834XZ0EP5NsPHo7g7Wac+x7Z2jSm2HY8OfrtQut9LkGaVb1QFILXhsFYM83m3wi59pM
iQtNN5SZbbpErkEE+mmK8SAJTS9TaxTN0L4h63FIUImqvmTAX75qCkGkhgcLCncN0peYNL5niX/W
NPjDZsAu+x8HmvKsZHXUV+Qp6lP7toHaABRrQh6t33tKxytS2anSPhkXcMwvlKSaUH0uhjJu/Tuf
WRZ/U0zKIxrNd5jXqNREEcVFw+HmW/i0SxeLhBI2IoAV8LIb/HxEgAP5zKE8mspb1NKQQuR4Sijp
VZGUrR2YI5f6qw7mft5RfF0j+xcjsQVfxvNzo4+mKYRuvifA4TjGGqX3qXhIm6u6h8jUJ5qf9Ox+
mg9TKDlgW9XlgEZMNednTo8UNtMDZ6w/EIIUJXcHCfHgSFHwLsBK0qYqKhQ2RHLDXIloBFibo1P2
IyA8PxgP9VAOfBm6Cq21wlfpOVMeHRaEONUEZX8ec51LUDoGnPkbQ8xWL91JVrbrxFwlXOTm0FtO
FtdRMqxbxknc6WVHrtgGcJftaSSjI22hv5+ulRfN/32tUGVPFSRoYP3yyMRbayDeksJoyND4+93y
ttYGJeWA1inO/RsfrrO/Vjxymnk+vuC139TnCd1edF92kx2eMQoE2CisaXq40vlgtIB7nRWI8gJ4
u/V86Ql9JFC53R52wegOjg8CZTdxnyuNmjTJgMaC6yVnfP/c/oID6K9nJ03hD1Z3pxm+ZmO7oVIh
RxmmL/TndxjzfGoukBRBkpFhvYBKIMmw52wfXrLkpi31InxPx5eVY8lq7RMFhRJsuiurcboi8BtV
J+95e9tsTMqtLp+fr9fToBw8e0laketCUPPQ38jVZvzS/J6oKoXijJoMtJRfLbk6lNgJbpVAReGZ
8q8Nc4sGOs8Y66EoNCCvgUzwRF870c5KnLIIWKjCFGK5p1fHHxTmGISEG9UdNkk7w23zyoJqCVdO
dmtZ5po5Fz+zXGiZkLRv/tEKO9vZGs732oDjkR6fULTASkpYGZNjKrETnhfifCGf1L9xCAEy66iS
1TMBIb2jP5zxCLkQuapdId0TMmcVmq9WREfI04RwgJHgUmxBCWGswBW7ZyU+wtsvje6ZCifuKJUB
jAWPODO4wj8c5AJe3QxXI3t/f7ubDo7Fo3gBpBSPViFPqhYxmGn4asiaNKFl7tD8RtFLA4lJl1xm
JRXfxc3lPjvppb/HM/nWMpDHJpau+KhqTYf4TNC+mhOQer+tIuqiHJ6zAuKmHS4ED8s/PjREyjY+
+EnSycH5DMhgp1r+sBLXs8vfP6eaooqpf0xxLTSZdYGFHzbdcJRGiLI/Zm0mMISCCvGk8RNuGyS4
RZbCvtku4PorwEh1aAL4bnFq0VGbkLjS5P2gYeAPcTjP+gMgsT79iyduv9njkA02HT/ft74TF28f
6wOvjUr3r4S7R8sFz4D366i+sD7Py6L+S45RliGLTTZ0izm9+q/pYWs6tPuF95zhNE+MYzbpj3dA
4McQErOyFAU0ZjqwhjavyE7ZKLIKeG82WdH/c9tOst2FPFGQZCPGtk+74WJ4KCttIgTC259i7mEf
DQlqueWk9QzBKn89tl5UuIeYgaJtvLFKcGTVTP4LahPjT9cpkn/8gdW6VKd2VNG4THQBhmyoEUqj
onIuG7u2/6XcUZXcQ0wz0GGyP5fQyNCbKzUSI7Byl9GHmetv4mb9e6YLXQ9zVSq2HHsjO6t0NMwQ
b3vTILNBEJgn6XNzTsKILXE8Bwx2CMFhMmm8D/HoEOyvmlX0YpVD90L0Ez+1ewCqvRj5PZ1VUjiW
8UFNMpPfmqiyfnmK5p3w+AuBH3tI3Ma4hgGE8cva6g4lYT0Qh1cXB+Caz9Lq/vbqiNN2shVWg0ho
IvLq7YFgkNK1qcvEs4TqMw7Wy3S4YQf06T7qCYQmlJ6X/VwPPFjsKZxTP3JTvTbqidK4Ed/mJZGN
sI5FpP8FKJzoUjL8N4TZa+SJ9L0BMOvEOBWPLi/vHyGGoVcSC7hF6VAjpNDjuxj+Q6s7hOl3iycV
Y+L/KflqR59VC1KdMOpOFlagpT80LtV02BfTTl6Ng6JpFhAMjf+IHkHuI9vrSbAomCsvx8TZvIRc
zkDhqQPT3WFrN5Y5Q4XVd07CE4aAATspU+D4bOzk1Mk7U3FYj4InKoFXzwdyOfD8VDfFVHisLCSL
1kMUp0wN8kLvnyJb3Sj0XUr8PUVXUCDqVKjjIDhdpX58BhnYjODMqi0/O2aYJbJDKOMOEzfmMhZh
6rMTQbQdSd5n1GaAp06g/8bWzeqc/Co5Is2ZOL7LmWF0KPL0M9UoMrjYkPgffUwtkSGYwPmCL0lA
jLJb1uR9J6h2cLCPTvjyUunlkm3AuyFZsiGq8X+a22cYD2zqpWYnhqN+LTr2LyBauzErF+N7e8Z0
89eftUB1SPJBI7sE7dwEgx2EdgKTfLrcqpJYdOZWUKLJu/cz/j1z0RquxYKHvRRLYKaYJX9wVfJV
frIy5xxWeK6EZOLfIZtLUWyN5vwCoNq7eUrsSZ2Kv77zjwKpaVo2d5bxHYQKDURBs9Lr0eXll/Sl
uO4xc2dKsuJYaFu9XOiMd5oZF7Dcf+w4z/6iT8lxi0x8E+Q0zgLdSWi/Zx2LuSL40pyJAGwHVvRW
NxwWgS7o4JMTzC3kxv8tSWtOt4vBmM2JAtgLoW6TE16Am18C0EDddZLt7+nkIvKFxnzsQ+nGMUyU
KqnBwS96ZmojxjbuX2tN9PXocLCsVt1VkXRqYv9SvaqFHCIxb2v5DpLnpnPGth2GQ3oaYNzjine3
MpDio7RdNnqPa7P7Og0jjON3H1LayBkLcxTYpTEXxLfTtcbfNmXbAVm9/28kJTzrcsk3zgmmby/C
ezRT7OYHorkbTR5CbNgwbojALYf61Fa8XUz+8dlHBXWOlkDSUrN+GB2h/J69WT7D7bZA0EAiI9zj
rzaF6JWX6vp2TvV/YLwSG8VilJYAizUkuF7hLW9K67WeasMsVPc9Prk6hiXw6pcaJA6tbkQ0Wv1W
hp3O9C0UQv7HG/N34WWJlBjQftioObc8D0iQS1b+i1VnqtlUEkhLU6eDqC6m05Mpto5RemCXrvCC
UbogkJPPrXq00L9CVAvnMHFraWMj/ZOzk+ZIbLrTP7If3owmSulM7sgv+ZwG5OcQaFhnE1jw+ctJ
ZBYimhFzynQgoLkAKBhSdFtGa6v9c86XZD6VLh4XIZ4OcXUbq9dOrAkKVV6lx/V3roPiqlQ5VsBr
+JwmZGzAgzLSWyEZa57tbhqqZX4S6Zzwe+Ne3gp/22fMfizbCxLuhiKi7scHejKq5TyfjBipIrjv
Fgs04TC3OCah8PVDnsdU09Iekdrh2t0JcyXUYc1vKBSgjuLPei2omkXoeJ3SIgmaOr4pxjYz4zHO
7cw4mIDvptjj88riHYA/k+rvxiNNfGwKf7XZz98WJcsdEOk+KPeoFH61XVLqx4bx0QVtjRL7Daam
jBayBnMlZiXAAvB+bH/TF3qi2HVXYSu6d7zZz+eWMjveIt8atmqW+CqyYN9xDTzDZkr5YJPnfIwy
Oaxco61K7k0PuEHbiffkxWZ0OwXM4leGHMAxsOKlC3aFMqWhmqGPchzg79+5/Sn7zK24T6AJ6aZW
jnVya4Jc6day0wM/aZ4n3trQ8zsIYMeXcDr0ZVLFkLl703ly1EZ7pOtpFuyiiumgdyCRB05PQ1xE
O+5C6chi3mNj/jj+z5iqlKNDm0ZnLcmJanxNK0b0o9yLZYuYN4wWn0SqEBIkX8NMxbwI+f5y+9Il
agFugrZmRJnTNPT7kg3oiNb/r7mrNxf5jxhmgKAABThmzobV99yW0ONlsZGmfhblTdMlysEN4wBW
uu1CS9MDTJOziktzZ2sAvulxseWdLzMPRhhIaHMsq3sUykpWIbBfWfeOKYPQawDdszjUOn++uyRB
BAHmSwbNh4Mj8b0mrzl3kHWAB3DE5uQh+KsNNdaH0i2lcB0oT9bDTlnW5qmOZigbcILOlmbm/yXq
fFUgF2nF/YwQBLfHYZMgsLTtgR4rBByNJRt2ER7q7wukx/UMJLgH4GvfPpNZGM8XltW0aj/rtGDd
Pn5qL7USC8ooyRmDLO2EIoDGTRWPMHPODv7Wa3kwOAjHW5jHqy0eev66zV+DeP8wkcN3dE6xqsKB
L3J4+xD3tUZ9pcDHnrnlIl+Bc/eltGkrtlZmfjOD4BzaIia48xnF9b150GBTxEe36SQX02WTJUHi
rcUXAZzbbGSTz92oupZFnK4jOIQ1d4ZX8hOKypyMqFGXp9VI0OZ5p/sjx71uDgtlLKi4Nn+gUcCu
goljEyiLTv6h5/Tbz4a0bPTbZ4njoO0T0vEPi6VKMMXI1Lo3iZ5HXVFVuhGWhUkW4BKcTOEg1fWV
u0aVrQzbsc1NxtJ/v9xU/Rr50/9cvU/VspuzdkjPug9fuKELQSBGkhvrx3JnAZmslgU/Ag0RmKu2
CNW5hVOXztR8isv2RzBsIanQVrLgld9k1xX3sgmuBcdLBbWOE/swD6qiRfObJQRpjEdXvscq/XsL
vojbBNkaMaz2RnuWmpyxe+LydyYyBX9u2q5vQsSrjNANmAInrV3FrmyIlHpj4heh3T1XuX8haKzo
xq6DihApEITArnm2BuOuMfIMH5XWaWlNOhBhNwX0ea3I+GkuxWg9yKhsb0I4jvwtzO2P0+xg34MV
B1Fjo1buoCIpsXe89GO9D6/UjyX92QIZ2Z0/jpLiY0iKJ792kMy0V22SMXov/kHrm+Att3Wzfllh
iR1OmHPVBsQlTn/xevFXBl5v8robyzqHwvCW8fN8W6ry0qbvu4M6jgFVuXHEkh1fYDEjIhsqODVE
EQkTZqDGMcZxrmJ/3miprDSItNcRBAx+7vPHgmgRL6+tvhyucKUIu7Kf5sKwJS/8Y1rAuP6Z1CQj
xFzUdG4P3U3D2P6EVQQNCsxSk4Qmn/S7Bk9RlNtjaNJVwH2fMgVOBt7j54RkxT29n7njzEZYMhjb
xYcdEkdOhMmV6e9YhjultjIzBX5fGs6RHIm40RkDTERzFjvpqn3DvvE9Z6jVcyzPJOizX6syD+JB
WiT4w2o9zU3m2zcfwHr0zR3R2FZUyBI3Wrbdbe0dLml1Vhg9CIjJPKAC6Jb9AiJMGbuc2uD9gUj2
YzgTgvFmD36y54v1Uj9/sFVWknxDBN1MdSAGdjBdKRgANIHKtOMPGk9CzX64X3e0PzTLee8ceGGO
9tI20JUk5Jr97BPy4MHhYmHHEnNRYwpAg6SJ4vHi6RRb0ZVORKfUQA13RLzTaGDmRsu6pKhid3wc
S8wGnqQZN5qxHOrIQXqMSTBq6yEuuwSuayAqFJDMGkrMfjfFQUG8kpNoX7KyhKZrypEfOcVRVYNJ
SrJtx/1Tx64h3+TDq5xVvpufrxFEslhaa2D8uaZmcw5BcryeAqd9YW3zJxSt/BWXG+VH+N9S8xTs
E0FFgKYRMGsiFqj/CoESr/vttcECvCwJwexDVnTbUwkH846vouSzqzYIYomf9MVi3VnLCOYeIlgB
+4X6GLYRA+gYseLZAI/BfRtSE3u5q3XobQbwOPieeBGrgRV4EWZ9dHH8mfbfsgsVhsFcg1YYjQkM
LUKrPUvX2/6nGIO0obFWtofCBTISWxQ+oL0Z2S7XLInEOrd3NdtqphOfwPN7L6fymLu0+KuZDZRZ
WynwJN/CZLE8K01K44iniGXJUTvwcTShHaYAUNfwMFP0qzOWBtUQKL+fUyAt1BkAJZeL+LKY3g5A
ajIuFBIQFFnddcRtmUkeDt0TQE50x3WHJSQ7jwCRq0Mx3nuh+lmFODg3rJQdQtR+f8Odcqm70N6O
kIdop0266KUhyI8MntwIFSGCnlCYnjl2ppMVb49/2sXGLz6Nfp0LZTHkphy7vQtX09WGQ5V0ePqn
Z6Sh8vjVYMfFjxzLwQ1lNQeLMRHYGmPEiqLMC2eStx8DPf/K3b0ysb//AoncmfVLjpia4AF7y7mw
Ml7ZVt8hYl1EUhh5rgVbUFennZmdIDmeaLRpZhqzrvrALaiOzk++PMzRKz+Eew2Rv/PJ7MtHn2Y8
AiU4eHNyOqWKza3ONed53Sz1VyVrzDK0riIEm+r3qoQIKrxWGoxPyYoocog9VYR7LyhsXmIZYbma
iWywBRJjMI2kL18zNFH4mm9shvpsm1AESYhqWUt/eLv5HTkb8yrT7fj5NgCLCS6Xb/q9KxBvRA/f
u1hH0jg6/eHJfCDG62dn/1TMsDbNXqqwv7GRVfCjwXXRdQluz4dzubDQLIQsq6q3We0sTcOG+pka
rJUVLEuqFKqoT5NFBO/hTlMH1cVuwlXtLLQbVIYZYXwyqXOwpAzVBuHmECJiyD20X6j54Iwfc2Zy
r3jlKzqRjaBF/ItuE1SRDFfXdv/Nuqyi7jhXeR1quRWlkxyKduuhci+GKJOsecP9t6DNnhoTbg9r
Fe58hmQ74UMCObu0bRHsYo03dW4UtogM13SjSuQx69OAl9Gs4TE/U18DzeUk8wNbYfhqxKz7Zjuz
sW713OUjMqy6WmkqwdB6LaJlvwoN2G/+KGl2EGs/wPC6uONfK5LVlslrEaaRw0iEQ6KbK0Otc35D
lk7jv5iE/PXEYjeV9iWq19AjJtuy1JFIUxEWRkebjTDq/PznrJf9I+nLsDpsvc1tzxbSf8CSWZLV
y7VFkw1G6E6oOqb4JyBboJ7eEDJVuPGT3VHj4omDZo9LocJsCzZIKszUEDDl++oGnbad0AIE8Vz7
+QIRxfLIznONPwFOJJ/v6wTW2tXsX4NmR5BhI9S4qjjutovWx4W93OgLPZ8xLBOCsFjX0IIA2dW6
MUOsCYLzzbRsT+KjbIdxgZGcm5jo2+gAlscHElhZKgQSHkhLtAX9lRtFJPERu8r7hDrtYiUKYrNf
AgSFhIcPybMTsVqd/RPzKEM1LNyclY9e6Cn7hhhK6CIVCE7vWLRmj+OBogfCHAwr1v2nmb006qNk
QJnPx0HByLIOBYMy5GlIos3DIpu27SI4gxpfnHxKPnZS7kvrt0YVCNkX4+bKRlH95OtBnm9+bxRW
Vs15ZrDpTg1IDH+PtSRGt09R3gLnYQhUTFLZBHLLI3jDVdugPIk7tLzwESLIm6dnRfgjiZmhvbNK
Iduw68KAvIhgW4Z+Gr4JNfHRbxtVUKqs02HmPLtva2KrkYJ+9YUc5eQDDH8dvKM00wPMoqKgOBj4
CoKjWDCBcKpyIJ4/e23kMxeUV4Ykvd9Y0d45ER9RiKBeK6uTNK+8DgAY5aT8+z7pgaNM87MeJsVF
T1Hun0PFMtHwX4QKWdIJgLDnGvacWsNK/R0dUzlS3psAowlkkb4oxdleN19aRmHfs2WgNArxCSHg
ONnLi46Rl1+yGgVwMMe0BkwG0uzoyEL5q5w8pzsP/sUcPDmzjahfxwfN6ymWO9nmygrInKFDWXos
XfG8O2rE1yv5XcJXXYeN07nR8eoJAFQ11s8OD0hwGeKKLVxFxZqV8do85wv+SlyPGyp9Zzg6Ubua
i2FRoHInsoH66k7tdQVRoZq4r3zWZi/WfBd6ZmSkal3T6wk3TG7vxVbvw89Bzbd/YfsXONOCA4P6
cUrUaDj3eFVMacLVfN+5vSTnFSY1/jkFlaW2ox6FdcB4A0jVS6hTKpns0JVmQlp11BhRDWa4AfjR
Jo638hST+eRxeC8QzfQEQBq6SpswTkPt1oKl/OshbbIg1asKhkdsHQTKD8HLSnqFkG4KW4yQw4Eo
dsUFAcPR56pqqqyxi8ujjw6TcAB+zLjRumClV2GeVOU6YukaDkoGjeY7Px+cBRLVRqRT+jDz3nGM
mrpcmcXbtGXC7MYPBAt64fddP0k5Xbj9N8L+myxSrtfizlMbxhxTDPEjzcJA6EJc9CMfYMILXr2+
VPVFeiBo/4hR2KrWVUIkmxrWHyl5DtF8MNNIH3uDIFxhvnWbQkJ5EynLkn7y17vpGGLWX3Y/OlL6
ykZ+H7UOfeTlt3sS9Px0OeUhjJcSi6kR8/34BNfg6HVnYW+aRMtCbOnH8Qbh9/S254QnWh33+HVL
j/IcVzlDv1HlPYE0MkJDEL1GUNFcuH3ceHh00LpUCDbWuzBUHcd6ozlWdRqvWHKWicLB0dmCCSG2
JoA3dOCif+ff4a+JY/E2oqqGHSwxrN1ie3YPSGjEMDz9nLwvdTFes0G2vrY9+hPmsKTmsxv3o7s/
NHxlWzj15VtDVGJwxHOR+H6GxkeZVLNFPPTZVjSN1b2Wj76pmppgwtUUwrLlatKTjkMXpK1oyDi0
+qxsCKiwZ2zO6VQ+Y6P59/Mc2D6k62HaF1RiIMfnthKKI5H2ilUVnO+KXbucNFcl7BZdDfNt8+u5
y/gVbZcq20NV2mNxKgA7GSGMJaZyAjrVpMMKp4WTyBMqeeaszPjZ5AJMqwSpcSe5h3g5LsyzTfB1
/7dXHj0V1v+P87FcL4XrrAIM3f9ejhZDCRh+smng0RaiewhEyYcKY2hHnk2BfUGM7OKjx9sYwvCI
YbPuXCsxw0+Pb8awYPFcScFMUDMyYBGT9TI9acX934JsRYpodWs5y6dJ2wKrtUqLT613WDVnOKgi
wDAYKgaGPu/sWLjR3Q5tsE+L+G81Ag9u3s2wwjJZW/tqi2VMdGl/yjVJYcjx04zoAXgLLDdSt3lu
8g1rsleZX/JpJlVyPNpPSToWFqBceB28TtBFGyjS16ZxnTsut7Xz+Xidi1xd/Y9PZvvdmc8pWdeW
K9fpEx16dY4wgZV6GmU7lVv4sMpdkRqrqpmRikj2g2oNMQbOjqxe5dWNoKdSPkifF4mnPGWpBehM
LzSg9FThtv3EZN9Yxv8d7gVUcF/xg7oqYZluYyTpAFuSeTzVnM5QgqjKXz1tjxyl2Q1DROstYCmP
5nMm6KaBXKKLMYNTCvv+W9GdLb/TyTUs5/cb7MOWfqixIONICuM+7Fuigr06akO9+1eCKpD4VyZj
ucE0kr58fs0xUyyJrsF6x5UoZaO4TpKD5u4YbBqA0I3JLAW7n/nXR/ugf/eyTGccbRsVzBA6Yxth
IAc2AD3BEJMh60cpMySYcOFSrOpqCKCEYWDztM0Pc1sBi7D4+ciyvfkgpcKl2fh1ccXf31SvlY75
L0VyUn343qVu6F5M3I/s5gYELXFhJtf9UfEdrnhLrkRErJyniV79hqxCqsHNp/iJsBtAF5lAUcpV
Qe2gL6d4FTmkZ7LrC6xZpoD2GElM5h9s0GMa4Z8/1tEBk42DJqzTtQwanRpy5WczgHwWmK133Rzh
2XkQ38w3O5/WaqUcEDdZ5DAEAiBR07EYfl5zhoxDM87F76noozCqGtneVpdQkRPxW6dvTCVWtzMh
y6pCjDZ5U6W+SHuKTElstBtIiEsmntXZcX3efUPA+2uvXLZVuqHySHOih23RPcHsVMqMAUOWo07V
sYeJydKnvT3BHNcI1fv6yzsQnIph1h/rCcyN6UTZU2pcupfzBJ264AlbKemakKCA9cQBCo8rPMik
ff0s2ybsprLcw2mdsq4YMlzDO/slZJy/Iz33P03t9MBCgQCKibA2ayoz0HaoZBYxzG0ZeXMRD+0N
rJaU0xUUgcd53QsA1k4+jJulKkjADkF0FPDTkPhhc/z90rkZoZOj8pU++tgJQqvgmKSjG+auk9VN
EnFhpW5oKSRKOJcRKSCLnxuZ4vho7vn5u5NV7qaBPX81VtFnp4cIbgTNMD8FskbdWnkM0tmWNqyG
+T8AopQOzo9vK4vFrwOM+aux8Z3JdT0T0ZIxNxZJxQha6krtddFmB2406LrsNRLaOVnesdu9H7OF
9zEB+O1Mfbu6fzVZl5n99o+2UJbOy7U1zt/WTRDDlgbnN03atPia7mZc+gK1LCkpNwhgWy/uSvRh
9ho+pwpHU6XAYZ0tfkRNQ6UVNW+vcPAHs98K/qSgAX1xpkBC9ObnE0WoK7xgx58WgmGRvDriGnVi
AzxFh4NNxWrpzyEcU+gpRFkSQ5Z3poXSXdleDBmfPTwyvD7EaaXGD85JgrI9o5k9Vw2RlLmspK+c
ADPg+QKUTfCk8VaT9rcLN2kpk7QJ7HUdRkm/upzPL+rNswCvD1WGqtaOsBqGBPvead8ajBpuvVpO
eLfgXWvkELrzJtDMyYfNUg6mEEXY1iwH7x0SXhMEBn1AV5rGK82fkM7O9uNNe1ijOBWKJRPs8t+x
grcyls4s7NiJrLWeY+bJcUvB3+scKnmezJGncVp//an7Loh7To7GDhOCgAdWqGH3kweqA5p4UEQn
oQrfWvZva7rCLlFfGwok5VxXSTL4yJYJHktpGNhzfTFeIUchAz+4v5a2S3C8bCd3BgFjSPu7dipD
0XQp4IAbx4ZM1ST3RHJKDIfv0edBqzLsNq6PMkTBJ5Qd8ZCkN6BrGJnZNritpU0XgoAZyGJs9r4u
1tT28rXspoO+h+nJzS8O4GnbAEPpLwDPFyqsgACZOg+t9slaj80iVzBR9aRlNtf6mAbOlh/sRprC
VOYiOe+j21aijqceRtVzcKgoiGEMKZix044rs5YNqMlLVk/UHI/kzpf+rbxhaj2oqOJyhgWez7fs
RAXMs/6UD130h36aWoaRdJyWnecVN1Bkm7eCL0q24LYDlCcJiENhYufkYv74UXnZuQmKbHTfDk1v
jtxsexYsBnCw65pctBmJGM5mGjKySBad42D1EFEDtCRnDxXPZ8SUdi+tgIrDL4to5+acETT/8UR/
FJwoe3qJg37qIKBFI0Fr46p6LmV0pPTuWVabnG9r+IHEnl4gF+MpKvu6/64XjE/caapW8q2VOgIY
YpGsWw/Urq04ROE+tBDzn8fL01rpQapt+9Ht3BMAlFgF0J3bm9Y7VGqnHvB+2j9+ArKxtFj2N9u8
J99L/qlBNTzpAzTXZ55JJPjvqUTVH/Outw44isl3Odj7u8qR0nQk4UI0jiwxPcx4SLfn5mmOiCqj
U1hZNFHvsAAmY7tzu5SrfViFhlU0xyO7oG3vojMBtZy/Kuy4eA7XGspNMXU/Yl1BRW+ji2wwsTWF
uF7NBuZSQGFZg16I8+ezLMc8PdQfnVJ1RmZGZVS3WUlZ75wbzByKeCZe6Y6h5sfRegzh3dZ7fjWI
XCLEyzamw2cvSyPlhEpkUnK4OcPMzw4CzQM2zqij8LUBxXb5kXCK9q65kfbveky0QK7dBHRK0bU6
R5X7+08+9y5gdM0QUvRvcFpNVrrIF8rouvFbplBowMUFN+WkRGjjDj2hZP0WdRd86kIffQz9E9Cx
yfVC9kN+gLJ+d5LaOXY2zeuCp4sN0BEkcjoJihhHBy/YXdBIVl+cv1l46be/1N6cfkC8EkG7FbH1
s+XDNGmXCEy0CDK8NsXE5IndgQeFaQrKOT6ifLs8TXj1EI8OpqpciZdnrCEHrgbT3FFbiKrNPHPJ
2Zx6N6bvxifYINK8BPydJ12UGFOswjyl4FPPyM4UgF3hvSblgZO4HaMYJJwARCmpfKLEPxlTolCi
pvM2QEC4JdRxWVf5dqPSUWYsWbFZnruMBUQ+ZwSXIBuRcUOWBxlhOtliWoPH0FI7OLNVUgk4rKEn
mUdVrf1N8Xe+C0v+h1U/+9jrvRpMG1ol+/R0JxCZvquuSh9kswFOBXX79JDP5jpAln/FmsteJRDe
kBgcY3MN0ZTBUsjYcDu3gsiFUm5W6h2OqCXTvE9XpLiQfd5ruuSkEJP3JWKJcwZtZpz2nW2MWVkf
lqOqw/FBHXTQ1qrWfHHzW/ltG3xZ5UrjKjXO81sWQ9v+Fzo2b5RGtq0nyWbvpZ037j1sESLjXAjy
S2Kt4lI+sIu0YycNmkQeioxEiVBP580ei1MC7wTS1he2MB4AP9D5PdKjXhcecy6JJKj1arMomNDK
Pv+q/f/Rm0TIuE7Q3A4hRTubEmjUAfP4kPORAylZsP17OVZw7KGjdWx5Vttmmp0DO70ZRj7g8yRw
aJQ5WD5NS/ohLwEHhlY8P/xQbLzzUokw/YB4ieE5ADi/FudB+VJ8AKoXTWLQwj/WjJiKFrPn55xH
Ay56G8Y6mNNGPoPu1+iSnrkydUdne6DOFtvOWZB5cMRPLkLObu3SZPeA0azv569zoccIbroYvKOA
IXhltln7Gcwnr/GFoF0Fzvr2etB/77CHiHxLu3wGWLAZT+YTmBTMjn58lSzX8f4TGEM4ingi1s09
trteppsmXmYUrzJfivfXj8WBjltU0lNGYFICzLD1W75otaO6fqovg0GDf281gqTSK5EujxGhiGgn
Trbyuz09sqJ9WpIOH2mHzDaW0OvjkdiuKebDzcUJDapbYfo4ufJljbTb/uP592pNtTG56+iy2jFx
PSbtRj0+TwT9rlBnalzTPIENVEe2VK/OW2dLZYaz26ZElgmWvnaE6nnlCwEpdgZQri+2YShQmlGF
4wyCPc6S5bX64+ZpJdH9QqQ6CIah5R0FidZLbiHRx5unfiHYb2mxoWIEGWcQR8MdelWR/CBTj901
dZKRiEHXB4kvmVFrwf7mRM/ABBi7dzVmsu34X++GQ4tKlteSPTdkG3X2ygP8okuAa8IBxh6jg+xP
z3nW/OflJrbTCqUUM3lPEPFN5+pfy8DmcBgpx5InCClrbI2XMGZ64OnmtfIKB6lFIvszkhu6L68u
W8sRT53q+InjOhOHOiQq9W1/diJSnflnzLJaLzosg6KVGICfK46/D0kskzrspXvcVcBeNxsiZ+db
ux+AE0qh0pfEgYmmL/X+GDoGWeyvJhsANjNYMjAjEJCeapAleBnSROMrwiML53QAdQZHudy4nZNq
2uuS4IJgIranq6JeKBpjLtDZsDl2/suRzrOVGIAmdJNkDZTVZW/iwswZLysLmisVEVcOAna+k1M2
tFVIJI727LXCA8X/8vZwFOZeFR/N8stpT1/reSXPN5zp4GwItw5F3BxhaediPtBv0STmUX9anQLh
5lnQLYu6bk9IBipmY+rkOlyq08UISpv0AX7MOlYCHa1A1CpAhz5IgiEJFBED/njMeQ0Kl/zYThOb
Ho1U0ev8rQqL7iuqZZiRenBzEd/hnEMe8YKnB2do7LWoJ/XodbbvluuXsFAMkBzny5LQF/VRZzUT
AUiQBAj9+FiqFjQWQ5ke6Fgzo8354dGBfW2QnxI4YQEl5H5aY3SfW9M+XtX9seso13hGwHAJsnti
aaTgM6jqxXAOrug1rFUuXXDdMWz2CzTbDliK/03W7pHtwbbDd1Cg7bPhjdCy257q8CvTUqpmHGOl
MKSohSXR5lJXgFbR56e1h0w0EAsdN6qUV7Bagri1GCnK9ZVI8znh0jKrcP/OplIvFPUTA0GaCVhf
tporHKxvHHuh3X9Qz7x0nqjRa7+pCv4x+zZPWKW1IwkHHLVp2e/pRyIxLnsPya+ykL/kf7A5pjw9
4EtSugkKFkStkOSJHZQ0eHW2tVvohpklYrkVzG4NUxQvHRuxHfnn7uH4Di6tc0na4hR2uftUkqYv
+2Tp2RwgUrSEQZWHapyFBV+l7FfZjgPMM69jWvY+yQ08WSwnL1G2gfO3PixpL4IFv5RADdlKsgp8
qBgdruP0ztDlmNhPsZiFOL+ZqWffZLyYgd6+5yxRT82333n2W73RPOF5CysrZvcG5rPRhXE4DW4Q
TaE0Lzla+Q5U6lFUFdq9Ni5BkfKdb+2WHMP0sFTJJfq0S0qi1HX/i9TsF2/yT0yfKRcx/Jz+yb9G
9vPHucppod/ur/ev/Ww2MeCXBWhVtfrEqy7EiGd224BRGuk+6hkOy+gBx6mK++Hrnz7z9Mucv++g
Muk5Eb5h7nKeyzjO0+2S9AisaiQXHq0Iyl7fqe/iwNkrId3oLUdDzLw8o/2cgEw6OGy3pQ4sXQrF
P4Awn/ihOMfguApmXTYQ52ZltzRoWysY9jd83E2TUKZEteqCSZNhbK8xOhMNo1npyLtodQPX1Qpt
DeFbA2rY30liviz4F90g7V6oQnluuv5KO8xbXmclUvab9w6KEOvpbT9i4y9CvntQcAVTLE2veD8U
WKuhS65YGkljUNjqrdNokwhUscQHqhmfpdV9prDTZYErlnWgHX6sp31uzjTs5CvY50uRFGqOaImM
ZMB7tBZVpcUYIzPIFYrIv3zZIEzdqrpbt0f5et+HlhFdevomUFEAWn/MJZp2X1KjresSAp4IH7QS
jnbkRwCHN5HT5tp116FygynnW9iu90NPgzfAYWGgBkr95iYhdVsvHhYWiBRaT9xNBXEY7Rf+rBQX
SrmcXOHHnqYCj6v5mOrFzJqcjS7bVHV4oo0q48cnebANGraks+wnCImCOQnu63jrET2mOq8vgZcQ
Zl/m0QkgUmrjKMkHllPehCjbotq+iB/tGKxm/yjqWUkLS6PHiEp0BMlAId2TIb9+wu5GSQ8MmW/0
XZQAiJzsBbQS2rss0DvShZj00OzdQ+6y2+hZ67BwWVjUDGvFKxgEQh9EEdvAEyOIBs6amcx6BzB3
Kb3CD4E4mpAQYf5XgJLhu+iflpbx7z7hbc+ETlMhblHlzNEt4NGbyCxZuSa1XZ+cZMX1NqmT+emB
zGN0G7xGYanuh3HfPQVbxujuMlah71tzb5CMolJf5qoC8IWnzgt8Gy8ijTozRVXhFxT1ckNrwn7m
KaRVGPasZOhejY59zqXZ6/Ey5kKiK7qz5ocp3exiTwlLthb+Aylbrw+zMlYn0EOHtw/TSHmW9tqa
itlYBAMqD2oj8G93YgNYZzCobqElUaEDUYOaAnIfghvbkOJV2XVxS43kgiJWFCfd/Wy1DDsPJOGY
C78kGM7JvFCy1JbjohlRPJavTXyb7LnmwKUlZmULegDF+amIy/QYCjImHHUCLbYhWugvHwI6dAQe
DDV5eoUjqN73aXSLernA8RK794KqZQMDeYnck2LFbxG0nvn/MuVys/HemMoIySMvLV6nWmlpoF/y
RlfustqkquWIjJVyqizoCH185IsXM9Zo6Tenpqh2r70uXjI5Y65uc1k0B7huVP/dhOnNet6TZiKM
xUejTukJXFhgq33qB92mMkVIApwX0dj0A9vsXxD0YJxYUTCAwAp/O+7d4RaxP3vwV7Wcpb9SdpW+
J6r+J7rFNMKKTJllHYRjWjTwIlzl5k4tpXvYm3PTqRVJMNaVQxXNocvdOjjlmxHxO9pCVQPfB0BD
x6/WQ2KrwA/lp8t0joGZ/QbTz+nhRgLXUlfVr5DfDterlqf+w1qKKxu4iTEcmt2XERfWLh9Y3KdT
VosnVrbrO/20qPbMfzMY7hybcW7hR09pGX2cwFim5eDIOwv0sXf7eBAvGACc6K2jPt4f3/DtPOZq
h3yfas4fHUj1T7UBfOxOFW5LTKGcpHuZpNzTNOKEN22DBgvyRLjOkfh3IhSM7dgEIgEaZrTFiwc7
th7LYoYNnoaGcjM5tjJV0OkqDupHsblnSWhYvkn+3RQXeZ+zQqMVhekTKFf7W6IMFmk7R7FWTSym
Cdyp3TnCfWm6kxLv+tOFK25Yq+7tUIaJfIwkOcxESQhwCayT1um4E2op6ITGwy9iGlDYj7S2/l60
uQX6nj7dCbRIMV6L5M/PVQWRctrw3zrJRdJdccRhry4ruQwN8GmwC+frgyidIBD6LXDB89csKAJX
48NIzxU0IEbAHhQpzzZRv8RIUhhLpqzmmJnRFSPXyI4stbxF8s1aakGDhho6/Qio6kmDe2KaBrMt
bL5AQB2yOEtDQ+u4+PVcDQhAC46QGyTw4+nt2fO3UKqOLz1ykrovGeWJZfE2q0M0W0vvsP7umOHA
agI3hbZnID/roV6ZHzljnJzMZTdq4Qiiubb0/HexRhB8xK7hDvDquz4CcDeVouIX1eAShZExFzTs
OM6pxvqjzr4qrY5wh9Bwzgf4COedhCY8x57tfWevnCy2Pj0qhZwREuqU7nQjConqZ14MFM3kxE9A
5bjZoQitUW9K086xDqQShbSctg4AJIHf5Uj6vjmieKnHLRMkP+hw09rZSo4Toeg/mNKPqQV10t/L
yyLD8i0xxHbFM4QjOD0/40sETHuK9NO6tLjmYyzFZxf51nuo0EVt38ltehxyisCLNl/LHX71H06H
14Q/mA11kI6lO4eV3NV9jtaUm1dPRE23OKP+Uri2OC7QBnGt4N3+fe1ui+1fXiIVrV4sFV1MCjJS
W+yFuapGeTwhWHOlkpjtvhMB1afg0X8ZdNfHgQszKHE6A0rYkYhOUDEVJMiZWow0DxpTS62Zp/dd
f2omU4WtSHAV5aDCSE8BNKs9yoRyWR452sRNCyuJGfjFaV64egWxMCcFjel2P8EajGV2/Fj+kpGE
RdRgp8HftrtlD4zxyy4orLrcpTBxlpgGHrbOk//Nz8hevXtRJscohN2wuvS3+MfjirGwS2xC9PgW
MMuq0NQ1s0WZANv/1DyAY0LG9HEhAxxLgs+Fyx0KoW6egrSY2vbuF555CRPMB3hFAnLxobcrpLi9
S2sjUXSb2jR6II6S8gNjL+1E6tp5SE7gWvzewSwjE8PogI60kDkC4lhB7zBV32MGPbzEEL7MlkrM
s+mGMPBe30pp4K08nIQCs+5HkSkhGVpFuED3KbH9HEv4AX3gEK6opSwO/5On/gk5CLdleUzee4oi
UBMKduW76RmMxaU1ftoctqHPjOgwxj8q+gW1eZ1QKu4DefwG29IKzUnILj5KzX04pMH/u7oZ2QwQ
cZuVn3eGdkSmm8m40rE9N9t6AlBEkWnmPQE+2z84tkDf/m6u2HPC5hFZvaCOKvyJIOWYZmslMQs4
cS+QA6bNn8S6MODy/5eSp+sGEwAE7m/5On/VLFVUf7127mjjHoOzzuIgLaohWoicr5043hwVwT+6
YVBvaWK0LwfU4qGEa+Xq4YrkBUpTQzmUSZNvdP0UKuozlYD0NFN9ks2TFDAT01glyqYoNGfa2NS1
yFtU8+c+tSR3k+uuez/JdKj5UQMuwd3HXnNYVEGOtskfsrLXtndmz3QF7D7Zd5bkazqhXMZlHBUQ
/58VK1PNXmyJaPzypU+Ae+Q1peE8xK9+ceWCQgMwvkQ7I9FWz/X4uvD+H+IhHHilI9npYSgE/yTA
oQh4VwgVbvCyfgHW1yHo1kFkhX8GxmBn5Tm+gyW6FsAvNvmCUwvKWdzEooi6NGJvEfUA/kSizyaF
CaioW2tdjnycaJKCWbGgjXq7g0s2obQJZmbEGMP/pG+uKh40nF6EZHxm7jaUHHCTUXHvPGj+yT5J
YWXNjSOkD3Go6OF92uF1Nqla4WyTDamrrftZXl/jfrG/c/IqPGgGsPyHdJOnsM9nLiRqcpLsWhye
vKgmMFacyDWbWdo+1VCkSBZ15/qkxFVJ9HCD3B+dAMZAPxD8NbdlpFycKkIu/sHj3JA3ArMIEGcQ
uqRICq32dNYnqaOiuzTk2poHdMILgH5oBVs3c3QKTm5dTNyujXiw38j3/KWuSJZpglz+OvDuByvY
ebdU3LqRZw8ZrtYKaKDf2LG07QvXK3snTYYDHt7SnyHrwGMoDbAdj6QTg+ryCtLyrDBVUMyftzfC
BnCGX+s6oAOoUXgkjo1cqiYOt+QE2rSGCj0oAjVgq54hH49pNDALDT7R6Lsplj8271DXx8b86XIp
DJLupSIcL5OFHN3gFU5zreKbsAHgmgK7kVqm3eQgJLxSD1epxzcO9DorMIYYGgUrn9UYltP5Cg1n
uJFWnvbULh6uqo2X4nwU5J/Ce5nb2dbsXB1fWhf0UdzQgHr0xkOyY9VHDSL8Qya2q1oC8siLQlrf
BI88lW8bySEKJrC2FWGIbpV/ug/n8724r/pr2xEOnZGvItEID4ROl/m5+VPAIZWXQDvOQdLme8NU
MfD/dkIMAIY2aM860m+apeJcYzX5Zo5ukCaBYbVL0wC6vhxI1IBWyWySHZYuKGEgBnUYySDYGjyR
h2teYu4fthfCSHLxjTt1p5NsA1jdv0v+s9A3hAKveLTt+f8C2nRfqRepW+mw7e2qZuDNQ8Hmo3Wv
/cpa6of4mP+5jBE1bsvgbFSl/VW/UNK6nFAluD1xPAWeGgMTl/xKQ7ZTtNCqdRbxaWaUCPf0Vc4C
TjSvxLjQlFMyZdSwBrLqsKnSbPGCfnru7nSx/gy4oOoO95vRzn7empaH21/uv1+N84usCcQmbpbG
PN/baKtYPVe/PHs3/Y3jhyB/CPKFQ16quvZiPt58et0gRvmBN44qkgS2/LHfM+7pTRx5Y8VtffgR
uvok/ABdwK4FLNsaK8CcDkCb2L26K1TKngGq2d5KCoDlRm1SuZf+58rZVcBXTVio6SNgTR9O1AqV
F1lgM2QsdxYvXqY9gRS8snodcC5sC5cRWo8JZvEbasBErfYuI1W+zYaN76qUCwM3NfA+L+SMqnbc
BskT5deje5yDx78PO6PeLd4SLQmHIeaWPmmi3Yjw7yRpNdvz45SpxPeiuS8K0EuyOILDxE/WWNvf
jYOsd7ahT2s4K/5v2vITE7crFYv5UIz/O3qoxXyrvoTzbuRtu3mQrOEeR3T1BSde8SFr8wTVRTcy
AS/vR/flFrn9xJRhAVMnzneRSkhSC893Bc48v/I+iN9WQtXOGmHkfg8vpeVLf5dfD5kLCUbIC8ZU
UDG3Jz+vvAZQKQ0ECBMKuDtCGBBdv84ZxHRu+qjH71B5b4/LPDMkRC2y3ZR9lUibRojhz5ARbsfp
l5A4SU6qPbRGAPMAxVqn1om1jeNAEz6pF0jtDMbYPgUoLN2hIzCvvjhGylVcUZ+6HM5/JeYvelun
E87DTmg+tcu4d/vIwu7k+sA4oUW/bQ4C5sJCLKwmtFIFTytfUYIpqgpUtO4myYPiICMWwWklqY7Q
89+7LGnrbGT4QK44ewYNxEw3qnbXDLwB0bMgLF66vZiyLCQ3SjNZCV/1v4qZZMMYRl7afQoV0e6t
A2IYbirffP876Tw9aNh9yPmbwrfd6WkQ1/ZPD1fkwrP9E92X8bnNICQNjDJXHnVS7Ds7xmrTwU/g
y+72a5ShB4cN1jpmuu+IJMXgJmHHTqMXnWthIxXjteKZJwlvJTDSNabp3lTOtAmnHXUDDByXlTq/
GhY/+2RcmLM5BfBqubTcUCeplCyN7P43mF0oKffNX1q0S/XeJr55wP2vyl6PkwVozadsJwYqwwsq
DWnlBlosVWiHSf09SaznssJaGxTxCrF06PJIAtfxNb8DgHMAlgHOry2DIcs1FZs4+N+CSBaDYj2+
i+beloz6udSlRi/LZPDTO0j3jWSGUVzgJf8YyBEdJzrWPR9tNF/p3RE4Nypy7g73cSGjmwezP3Yx
LFuc1HtQWkAA0Rjk0HIdC2vrg3PLLFMAE1RBv4sVgfdbtsH0CkznozF/gKVj8RK8lYLfU/KRm5O1
PomdHNLRVmGLfyktuXk7PIlBDUNSecdumsDRYciryUAbCbWebg8iehIkSOw6p7OoYFdgEoezRG3t
rTt+HGgsJ2qeVPK/t5elnl2uxSn7Om+0kBUuoxuPkmlWSHVNX7UwzeJ4hxwsR4J0ddpyaP9o7vU2
xmEYgN0K/44oy0cyKp+jT2bcP2E8elgnsUN8AJ42LQRuSSDAgse/+Jok4VJhTZTNKEnfTH7ARj7I
0cQBAYGuU5ZpnSBYy9qnrZmOWTDwP47F8ige363Do8VRPG8qBZKUMSURODkPnp2f8/qndenPpvmP
LdYx6mv2M4HRtTvIg/0PRegMnE0RS+Lm54sqHe9lJIv94NOunI6dO5vRayI1Mk9SQXI7qmDnEmVH
slDwnVwvUKZiXzOVCGqBejPyrtTLQTqDQ6vj8E7bdKsmM7Wqf9Oo8ZN557BP85fDLwueUCkZ+5Tg
wOYDvx7IWchxodevlaVq+zpKd9iV1BuR2VqtQ5lpNLvtiEs++nBYlqAM2EC/Qim2BnaUMTSM2Zi3
49UqfmjPuLRGk9D7IPkaCU6ZMU4U0YphwccjMprR3jd9SQU3b/K5Uq2mwLmFWnah9koNDfc1e7i7
JJ/a6ptuZw9VeCqhpZEYLeFxK5UEkA3Fh0QRfkFYo+ArEyc3zSEPZGUnXNW/o4hpnAkbbt0i2a7X
mU6mhXyHNwrBdeipUQogdcm6DhhoBM4IRvrv/3WLhdVTHT1cUwZo4Y+ceQqI2Ig7K+j3kwvg6hyI
egiQJO5+DE3MuxEJAsptavOyuNH5GDk4yZiXCikbeSMPOsheTS7hL71x/ppJ04u86gRr7DpvsQjU
gJKL0yHToHzd/CrJ3+aWShMjAOghlOU7LlCoOaBRmY1UEzRDlrh842mqhTqqhRdz7Jx6sLPXijIS
b0HVZWUoCfic2jNmTLazNcGSt4fq/wiw4hqsrEALIH98ZW1oZY5L+R7ClMZanB0Vae2TGNLBr3gw
O1L4fssnFK7hGhwOOVdNNXwuUpkpYqRv73jCyz4RNQGHs718e7kIwT4LOhDy9CmUAlJngoqtrGs5
U2GiEbgT+tsmrgxqT+/EgrwK5e5JrMR31TEe8J8CK/YdOBBYAi54Xi/+wesPi0ursN7FjTkHJDOp
ZSTjxtLhjZPIfVK5IGzermT7G56hs3n+Bk2fkUb79++k8lkneZ7oxPXQswLqfS8i6Fs9xqXD3Qgk
hJcCyqynLOrvMyILoQtF1ZlmiHqvBbyaPND7n7mp4Tpm5ITUVgNc7ZRhqAwtMv3v+/mG/S0nCewJ
dUlg/eQIiLwgh35m6W13btnZFka3bD00oN64kIbUJ8qoX5G3MLeJO4nv0PrRQLs6LDn+tzzXjVL6
bk+n+EM76JeFncjnFotUBmiqJxta2wBAt41dRk5L1kZf2ccVO0apaTdNBSAmknoVWYpIYS4h+9c4
P/mCUs+PV3Qz73e4d1XJHHqMwJzpu469+6QqOIpij9mkhvJEU3M3TRWF3/mzqjT2wWz7hV9PXNZy
voAAaVKXnDvo4EUuqNbKBMZmjqp6b9iDFQ8fd/su2iIVDUetoIAs19ByYFqnN5wnTjQM1exmpmmg
Xa4SVXQEI2StDpcU3IJLOYD1LBNd1sl8eDNwnMQEbmLbiQRw+t/Uyfyrw4aGztdzZDef/IaD9hqY
97F8wQZMi6wKQx49xM8XaKvc9apa4iFJR0JabdiXMWJDle9jai8PfEl0hWDU1MLTIEHMXId2Kh+3
N/2YgF3RLwKawOqxio8gNpt3xLVSlvYf9bZTego3XyCtHG5CqtxHNo0oy44Gb337P+4irnciDS3Z
XAjFqG5dvB1YKJZqx1uAco8vbalsEEa+Cl1He9gDpj7IlwbTK2U4YUQEvs4791BGmwQxhZh04MzR
khE12tj9z/h1YS6pPqspOb2DSZEpZavlRNl7AEKrlPjt3B7GdI7X3sPUOFjI9rK9fZpdqA4Et169
meYUaYfP12BfdVtxjiLcDbJRfhe2R2NpgjE0lkjN7KaAVtrQWPwQKUe1esfOCoJVlzSZ2vmHVmW0
vmZTWuETlAwXPjH/GwSi4lUIqrEYqKDWcXoq4dBioxYcyyirxfBjOLqSTDom4JYw9EMOxJQjkhj/
pHLtcrSjOT6p6rWn6yN++evlRJSfOoxgslSrPN8U+/3jyxCI7IFAg+I9/lbH24xgbym1xIuGZff8
4hNLUYfFaU7WTC7Xh2acbXQ2t+mm/LltCPcG9FlWQAjtjEd3DH6UzO3hy2GUeYbmM0yluq0RmFV6
sVihwGuRKEIqyTF91beDhu/zfq6UGwNI5BPrQ9k+pPegqZVUn3iwwQatH4PCGlwCVI+X1S7J0vD+
2hhrc1TO38oXMlYjF8xPYZBfja1AgHXD9KA3UUALo3LLzTAhKpEHQPwHaDnXzLaf6mPTyBPU5niQ
98gAm9E81GVlQixt08jH21nrMzGybD/wE6NtGbzb7eT363N0bOkMZi+I9nTVQTDyjni4/GOiv4W+
kBPWsucsrxSgkF19uKscGVAs2idmdBloL/2S18wQkGLgsHJD/EhLJ/QeieEy2uCAA/o44UJOKId5
PmmnRJYG9UbRNg1ByTJvojhejeFfcN83tRNcsSkcAefXKSIGsO65eng8HfzEan/BjuEhWw7/OmP0
rztcUaffnsP3/bgAN+36cV6mEBrsRyYpMvJ2DBuQq7gsmU397+QUL3svcLCnouQ6Lo2kTRwOpTNk
dWFyQ7dy03Yh7Ooi6yGPRZM+iyHIwX3U15qGW/OPpNQhhB53BHzXT7BluHBDw2j0UEZ3L5QnzkjI
lIuedL1xEet719qRckq9xa2B/MDne+aeQPydsD4yzk7ghhwwGH8S9cxlcQKTC1yMHR/CVNkbSqdn
4lkynLHOMQ5QEUDwsiYbdveN0VSOwojwlqN92zvnpsrczQoNZlKEs90xLfpK3uMVKfoqMAEw/38B
sxj2htNoK9bIb4sJq9w1acUgPqEdETMJnuPCKpd5jvKjSgNJcfDHHpLJXtDaBb5WdPiAQFMx58fD
u4QogAwkXO2iEzBHNb8Ll8kF+E2mD4uL3+F3e7ZLqYvRv5XoNhvsDRiA44NXrOi7vdlRtT5WY4tW
jIttA/aA4ihbVEtsPEiywbMZkfUPiRiU3zybm+CGlS3thD4ahumAYj95T5oNeaT+KNY9tcC3tkpk
Mibe6TknZz/CoskUMlfTp00TLWo8ax1Ii2dpclRfzE1/ZHrHlUp42JqAABW1SVkLnfbfcJrcq3FJ
gS413sn/fsjWvNvZgG48mgO4lsCNXnzBLVwLhSw6zaQfWGbMN1XoS7mci5UTmJspUaaHNItcU/fl
z/kV3xd1+vVLUlu1ky5QzIqusdFMU7mXnx7YcP9uNHrBStYYHFucN49EaCR4qLl9GR5la34nSrQd
7HUnQvJQtwphbSVoM33wXRICi1mlU6lucykIbf5BUvfjG7TGQKP/6tWvfU07zgw9toM882f0zMwb
4UqkXmgZMBIYTaKDG4gLQ9l+bLboguGZucRX0A3+pw4sDN6OZ991Qp31ibae88+W7ycYZtig2jhL
G9rk4Q1b0jV4gDY14W3IwyqbxOQRGAeKJN6CIsiZU+H48m7i970nLGxCSUHm5MYS1nLUGGmpJBIu
uUFb3ID/C104DzwMvlMqAH46es0Tiu5zb0UMR1u2WJW12YY5aAnIw6rtt9eHILFQ8+yuBNuNVQHM
iPITTJU1ZSdBpKPxilOuUVNWiobxos1jijzIsS+/TuGYPSlBTuJd73HxGQ/4Uc9tMZdG5L2haOvu
tWOnpPNCaEe3BdFBJ+9mwMWq2Qc0nnQbBlVVXUU4ECaXjKbNaO4faQooUEjgyDMTX9rZm/4Rgrgj
vpyZ2ZC0cxN3avX82b592roexAKcwk5VGOq8uDu9N3kUn/dycqfMANsBxxBRlQNG+NukWXnzzVAV
MK13JO1lU6qvL+NkhCFyeqcR7beqSSjglg5kGVAEDH+l+CmFjYjZ3ZVXY1pxvDFTJnbj/NuEYxAA
pyJjMWujC9HWObh87OmdYIjeLOYGl34VX4IAy1Ke1/I8z2NeAknpV6WMsPhctpJHOOgkOWljdCft
Eg1gOkydIo+DTKSuokPUZU2/oY8rlYozIJrx0mIln54HgDgabh+Z8Dae466ctXF1FE7IDZd58V6i
BpVm4syo3E8Na7Y1U9XQme0+32lY4RwujmmIsqRAncrxIBl9+4LwLk7NrIHaTg3KRxfojlDseAbv
wzAxFDZ0zGq+HBtYs6A5PpDSS5LJ1Gdd4xU6nKmP+XJE1nfWxLDMVkvwM3oZ1S2CUoL9PoLfGco6
B1ae/YvzRZHLj2wBGeWtfBm9ZLU9cWoUTR7bMWaR04yoIyXRztrdsgxNyrT9cExjCsAObRlFO1iD
Al1RRSQz/+LmbkgV1YHcESB4gzksYorNyPjamQX4NJQf1I4M1R9W9sE5x/hA+db3SvAeYWVDhx3J
jqY5G6xWWgaGW3lDfKdFkUtRVSY6ICd6OrZCFp27mO7FmZDWrbTMUcQgOQLLaGu/qa2hvBh+av/D
JyQcnzQPaEjjr9Tuupnek2nqvU+ZUE0UdFRJpIdn1oMAAyjmISadFD5p3NSFsHexA1FFccnPkwpd
BKFVJJ9vtGNuVUxhnZe5blGFf7lWCNTIX5iJiNUODPI1rFTQjvqyT+UQwACqkubnwuYJego4MrZp
ej3fsaFuBR+QMLNJAF1JgdBkYtGnkXIB0BSLQxSWHqfM84+gKd8RbvFL8C1ltaE8Wc3Tez+iPX+v
TIiV1aik27wOHt5Yzi25ju7lpSbHmq5McYvvlTdiXFs3Ujudjpp8QfK27lysku/NzHB9WQRBZOga
/TP4RyAl7JlNNl2yUg5OdZDVnr8LQh9bBBytKPu0fF1due9A736vxrcSa4Va2efYPoxlXjXLDI0V
abAQjqaIw69volFz5YWpcUde+wx3z9qQmY8YK5TYUBf/2geKtoxtxqHDCsdDR2Qmn2+JTMwuN8Ju
VFRhq3OmpoLZViB+p1ARDRazxXJrupaMpN8awQv7O3gihwe/SdDZnU4G0FyyRxBoyMk+7Z/hmx6q
syIUAxfYOlMXRMfC5xIZiT2zWnIIREYV2RT0K9daoUbVkik/U1A0YA9cIlLy7CHfpydDxIMznBVD
gg4WnRJcghUUO6h7gSGqMEuY6blKiTAlJu/cmJIgJyziiUglEJ9WfxvjdC438EuTJoV7TQfaDdty
3PcBMUwOYrCE2pB9ptBnL3gw8d+aqwdavwPWZA4BvjqcgSayEU6Bi9wHK1ormnsN5IuL/cOoJCCV
+VH7qG8QJ0B3lDqp4o2bTtxC31S5/tfrrGXFFI+G7u1svaT+orBRZeFmDXCRZOIb1/S2jgc4TxDO
L10JxagZnUZcA5cQIHxwm9+wlu3a6yASxDL+ksBILJjeozLADqkmas1ENXrl2x2IdKvyathYlCe5
9QCMNSB7WT27BfM5CmbOk0zdYlwRM94WXQF2fjixNundkDWEwK/u6r76zawKwzUxGO1ldTO2BeGr
c/5+/s0pC7szhAqAGngAnEM50ohle4wk+2UTHVd2TShQhJ0B6EzwxScs9M2/nYShMKOeyyHpuFYK
Dbknof2D2/amjVAIT61LZq1zZOFgmZHetFZ0SCQN4gY0QfUD8pjbyoRA86QXdmNVvWRdnKo3pI+5
CIvn3IisJT3tEqqjBWSId1dK48t9YvCv4ZRu9FJOkbuvUoTn/0429YEMIeCdCEWNEEVpIDSg/ba2
iooUXnhLvavH+7CRdUCBjsPk+ge+fN7RcH3gGbVXBqsgvUJ4sD9okPBgAa/7BeCPkkBm5ViJNjxW
y7EeJ7fP0OdGamhilhW0EkH0IoBrYrla3BXAx3j0L/aTyPRezGbI54066lTiN3gDP1brK10UtEoQ
x9MDPF/nKJUxw6tAkFMPmfQiMjcXstJNfsYpxgCD6Ie0KlGT0ipfDwuvDcNrAcp4tZ7pLYDyug9b
fIoV0wbc+kxGAf7Ybvdlz2boZ3m5NbffbjLFcSF9v7h3dSbsyXoBQTdvfUD0fLfC56QhMQ34RZxx
SfHIyyWky6KjBCNBvF04vhPcT8vXa8VAz5dOyeOmOLPbDnk+t1Yil4Gm40Nc8/UnserJcNfOqKPy
CSk8Vbuq3NSiECkcQrqAvQAgWrmyhlAUxBoJ05hZTG5UIxDSAqa5vG2GnXgJRPb473D5x5S7IdFB
0Vh98nI+UHvWzhlv1zVM6XtQqvuBhoi6AQAOFh4O1+sSRRHnmMaXJpIe3EIE2BPTd8VWz8n6AUju
/5cZo5zJ/ZBPs2nJfwRnDbHQ2uS51dAbo2ITMDjWIwKGgXk62Qa4GTMXfZEQCK9jfKMinonXRwnU
R4xc2Pzd556MYXrbJ+DQMFAKCx6Y4z+rYZFWr8i78kUF2dLMsENesjqgpNYxy6H8ZRA02fpL/0pS
yrCja1sWlxQSWWWcp6FNTrqjvXj+TYHD4422TAdutUPQLMeGNWEZoh4MbFJV3md9NWrIPtc4JCnw
TxLLloKBBP6Aub0vIpe2tLjDYJ8pUb6+ZmFsuW/DRPqJbUyVYZqJYSg+lF+r13i0uMCUxM3Xqv/k
5f5NICPAKD/KazhM/JTbPCa6X/phrJS3zoB1Sy/3AUNLVGMxIP+vx7ztu5WvBpjz4mxZGeYlRSOB
hlKkjsZAbZYSPYb1qBVvDj0sfWY7mwg0jBVw/JR6wMPoEMj1PWFgX58L8Rr994abRekIUKJrzL3f
sbesaAmY/a2bi3rEqEWWNNZnAsEHZGdYINi9sBRiqU9J8/SkahnaNSOtW7ioeEvbR3A58a4N8Ykx
/0tHyWYwS1kj4tmHXlYvDZqbJ9Mu+H50tuFIYFQWjNUfxyXxPw9fdZYcoBHaQVFlObPFb8DuEHx6
YkgNyTvftG4GcL+3F0hmwcB26QL+8AR2egNolu5qJBpmF56vGpSpNgCj3xHCD9c3pGhPdu8DkOqs
Y8vfGgoUowHYKpAZNU4KZaBkQ6zk/VAgj9sTXX5kAYZ/GzL/7mpBeo4hbjWuN0yYvW28o4WE8n+N
HITPjSbJwzy9By+nRGg0AJgajAPUdBj7x8vglj78v1R61U8fPRaJrWO5zk2lip9j2PaDjVyfgcQ9
OoBmkYYTfsw1mNWIoa9W/k/Om435abPK8oEn082L0MM7fMNYEXoRCMidn+N0zKLB4xhngq2VxH1G
mT3LKiCnlDu7xhGEXnu/lJWZzVx0Gx5sLj8oYeztQDro+RS1JfrN/XSsZ9gSlHDVvEgivABNXcTg
rL35HsAgRgyUtaSJCGFDzMMkfU/AxYllTu4ME0DiRU1OeOfXitSNgJkRYl6fYZJUYEq8BFThRlQ3
JQMEK3CX0Y2c7+3Fu4JqAU3qKKSRTPQmOrhuP1myjlam4UipoMG4Xxm+3TKcxbVNzCnBulW6qCk5
bAnhQGIDkCFmd5D/IV5ZFcstTj7gpKLoxsWgjpdNz1LmicnQo2aJhje168jsogVvZQm93SggdiP7
njwCg57OGcmgZBJts9WDkq/4inncjnWk7s4kNTIHxSdPbU1c6yA0Flhs45TorR3EzguUBt5pZmQL
jw58PHjuSOIXO4X4GblXGNLtfu+++NtxxqFhyWaQp2y5t1eAEZ11D0xZyKsR5bixwxUkB0leECKh
VqWr8Ed9TupafFOye2Gv55ygpbqupkeUtEbW2Gn7rEoX8UwiOpGD6L/MfQGfI4alIyggtxLXadrv
D/XJq7xpiWf4/tC+hdcrZyCSXErcmtXtWAw/vM7g8+F9YxVEmSGsoQ6k7cOAfULm3DYaGpX1hD2B
1GSPAeh3/LnKW7ZGymTxaYwsKuct8RHrXZX4EN7ZXXIcLAlHChs4iJIKL2dT7Bbr/o+4rOF6Sf/O
iiALy0iRnU9Yo7rLH9GxK2P7EYtKIhsWvijWQPRfQ+9wAvHZI3hTk5Edw9ulzzJ3/2bEGhFMWhqK
5UoBVza3FlTnYZPqXKnkTMnFsYJXU8W6AdU1a/A1pgZkAoWvKu6DiRZmg5dYfaoOno4eH1+IfLEW
Sl5LZHc/zpj+iZfu7WmMTcMdsoPHKQ4Foira+AKdp5ezB1jsFE96FPcaXEzzbRlMz8yI++zM2YxH
9ub7Fc7f+5pJs1NKoTuEqjTGe87F94z1yRGUL/cwuOlgAHLGtvTqyCK2gkzyROEjtJ9H58uGiQpR
Mi9SZeuBGYGd4dIYhdf2SnZ8UgZWA4cHA2/apcj6BSGjKTbeRQwyA6urp07ySMrIHm0rxe9DPbjf
82tP12rXNrvSwQXRGa/6FHTl32pbBCE2vs6TJGDslvq41mFmzGt1lcgikYw4HIayaVnvVTxznfqi
OXJMw77r32ePv/tGSEKJ0oGBjsUhtU3jDvZXVt6A3XCIkoHwU9yI0OA7JueKAp2giLPOxmDDpjBj
7c4jauP4wNhwD2GzXpPgmnpxWhczWtqisu7MA/0tHM37uqCKRZcU2iUsxC+yN2QERpMoJ+4/YvC4
u6f1zkPoPeNuZp0GujwMp/8tP2B0z6OW6fiy3p00J0Q9QtMdzMv2OmwWJ1vaVv5MqvgmAUS6OPUB
qmebwSAKQxkPAsMgOGq6Pd9tgWRFV0h5E8RgS+J5WYxdLNYZsnw4Gu862EKKVTgR9VKcJs9QVKdO
qRlf43RjncY0OhCNI1RpYDpAqNQe6hSmwpEDPjM8Cr1VGGGilKe9OLFC7BGnt5pd1GJD0ZUD3Wr6
epTUbJ6ZeBY8npidlVMFMEKy5sTRwboRyL8VdNJhV+jXVajLjAzzmRHzhjKH8HI2yJ/u77JwpW6G
MNnpVglnwMLOdcMkIrv26ZI39FQ/Pt/67GbWL3itnu6JBCxhdR/9rVRG75PMLEnh6KfB0vflUKvq
Eggjkp6qBeJnr56/H9HaqP9VJc90miBUAq+wNr/jiDskwKVsC4t5gbjjhmkelhAGCQXYRhcs4Jit
SW4apKRcUyBbGOnQFiqDOB+aDQUfSC5UWs1Lza+D02TbRIBd+8nVUoQpqrAInbFvjY2PbA/TsjOA
xJjUSmgnjbHh0s89vYwTMewtO4intOAVbd2VPCX4cWs6d5TtIUQxkXYeieTvErPU86pw8g/rPnsH
mnYUntAX+nNBnRpivo73F3fL8RU7UPuIxMxxdSYEcMFFOO3qWZKi1lDoCQJjY1J570ZmXfaTpiCJ
2KgUXwE2RqRrBi91yvt0rWdTA9bNiPDO5tlSGgL/wsRdgEuEMtaINabTUeGNKakpviwOfXno3jf6
c0Wqv0C6OCYEKlDzbxAdzwaqmRJcv5gayaI3fIlYFI7r2j30JhAObjLktN5vNfcLigl2b35pGJqF
t1Wi1svJ+pQs0L0OA2izOSrwYBwqxXImaOYP6t5uH8lQPn9HsPxIfBOpYPpO25iWbx7RJDkic6Zk
S6TsEFE34vSWL9oc+qdNkCWU5EV7VjkLX9EbX4tt173VM7gnYdJy5eYfIaANqLdknPE4hrrp6LYO
Wya9B7lhdTVg9RCyCzhiikghpBWpNYpYNb0TCzUHalWbzW6yTG5DlwMyF/wPZGY4dy5c7PHpTaY0
Nsrn1SJt/B3Y+Ap7Z04vlypEUNeNKkjWdirXIT2Pa2pJ4wOn/gC3xSqSOzFofHXhW0ijdiqCG9Dn
/RJIcCsG/lB8n6oBbuT+wMG5g4ic3bkhjNqh/UkMfbAs6rheJWfpzaBJcGm8hH5dOHHJWs3nKv/E
oDNiYS7/5haPMWdaKWBc/DWy2+e35b1I2V68zeiUFfMI1aHnTkDTBbthYTQEbjGjsrhVrK5aoRjl
EGUj3lxW4Dm2K3nGsgj4vFzt+KGrzFSCGBkhRtzor2oaFg58CPI+k9d3QuPxJ02iwx+rDhvX4aQC
0Ah3wLUY7EnIITXudnruwggEw97jo0VaKA1yTGnCLEmlrD3Wae/8hXMarRtQ1DFxpP12zmDBOkkT
9oZy6KvS434NFZe4L5m65K5e37seFa3zdr5oil6LCKYeieVteiiqDkfXkV28qMpD+9JNCXth1c2Z
4IgF4MINQX2jm7w4tUV7/EJW2WNfDJHfj6Yl32i3uYehEDdduIJwBXqLHi97OZj6xoazwpUT/MS1
C+Ve+RCNDzNzcORSo1ABR/uZveoW5ZmEqtX4vzaNeXpIA4+uMinQcG6mV/lTh3FVIg5JvQo+p+WM
BNTBujuDmfQVml6Wo/evPunhs9ppaK3O1UZ8s8J30CIb+Boe507jy3dzcjaNhHulrjgcNBYWFIjI
z4envuBDqZCBGy4GLcvJFry4h+cdJLZBy0S9oAHyb5siBa/M1YHUUIGiESLHDbdIa7GCDYfzcZ3L
1LyJSaQu0yKWZLCf/ny3Gu9eX9zk+cC6glWiNi7TjsAaQr49QmoUI0RDiLgeuVeHocPQP0X6xhd6
c/FDMx+8zTvTf4IQGPEk3ZqGLwqFz4Tqi10rGcZkg2Pd2H37SL0GiGqDfHffesuiy6NDyJz6GFuC
V/NPMoE0ZQbE3YXHFwEdPUjaXbDCk9LTxEAB3Ryih9bj7h8rFWOqMd0fnwBfymseqHIY0oD/h+Rq
r3ABgsoqQv/6oFY14N2MLvGe9HU3WdaGc7lRLUG6tJgNzkR5fPUQDafjS4KvErrQQpUePgsGbm8U
S+rMnslo+JIG+67fCzSkZKpE4C+5h8jrH+u5Ez0U0/+KiWaBPMlsM9X2eaN0pFmInCHXERakYCeX
+XmlEeJ8tp27/yFMVXoRKc+dOGwVSzpfgksMKUAiWYkuzNZFKlDUob3CGOoSTR1+tRUA+WPaLeeu
nX5LoIlKyyg07jHqE019op5DsTHHIZBfWuCB03OiCjBl1D2glNAdHh3IU+1qx8psx4sgpxCoMMBB
FLKgsuEm9fiMoVxxvE7eCrfUIeK9R65w6a5x3ldwWxUz/Q+nPl+jH/3ilU3SMRM+CZZBky5+uLfB
tUDM5AmYLiUQozrJM7IM3qkoGMF5MKMh0FJSFnFHWlPGafhFiPzSSQ5dmXJoDeMo3nSSDgpxi9Wx
m2+sa0QG38SDElMMBFcVliEzWKPnqcOgPTIFyS+dTQt8hIuD8TLWdtuKhgvVMvZ4i/J8umavwp2v
16CnUg/ChqzuVMRZAvE71uP2NLr/Gl5x8bc2lwvRjRNUbsHilexEYpTrko4V6rvF+vInUZ6QdRrK
896l2X0cW4UYrwNVmc+TarGlqj77t3r0D5HjTCwSC+7DZ/lVHDtt8hX2gTbz0kTuvd4zLUu6WXmT
QUJ5VRLbz1SfEPixVVwAlCwFk0IYcbXU9E3hCkqrI864oSijo8fn1mIe9ae4Yk8o5cjVYtliUKcO
r6XLMZUvwzSqNi8InGVh9a3JryLElE8+XgmDMZh0/hI5Ub8iQyEjSthbJl9znCPbDWqgxFcLNKA0
mKclJKxblc1CKLh9bqwo8Tiovp6cy3rQC+nEtgv96jGov7utJrUpAsA4ScPLLF0lB2sO8VRr+ROr
qtjSkVOyb2KN165WHWq7ZESAqR9lPRNsxgIQjnvUPyFTRW1HEYXvEvVhafDhGXuFrUfg2K6wuCOX
mf8m7r1MsK/M+kFOXCOvwc/XyEpCwbXkI71YJkR3SXATqP3N0bsfNzFOCIBkU09wn7m6FceXO6EX
/LY+j+vDbowUkz/aBVWXazQxgP0O+K3tuqiXeoS9Op8X2eEd4xw4x+pLuoyMkOeZaqPGQF7f5Wu1
D2R2kCg9IdDJRBpQL7+F0uxBfPzs5zZs2h1SIzvG31waQZDAe8BUlQ9tiYq9klqlCImiPVBzxh2r
Nh+tWsCEdWmI6mQYoya3TgM8BvQLR5RsKWBGGJeFiVeLBya3U5HjfmKaH+Yl/8ucriORJwPcirV1
TcS5TiM5rt9RV4EAQqX0I+1mwVY0GSe/1LU7fp8qFuNES0Xuf/R9skpsnJGb7JDdfJijjd+MCX/N
QWzLvlHGI24Wmunwvh1RjlvXZGHXwSZ9cWQM9Shvm2sBAYJ/BBdkcaZWJtaKLCUGYwEuXlTj2KSw
vkr+MMJXwpia5uY38hYaemDbgU1oll9+KDGYBfSby8UDm40e/HmNcSVv+wTXWj/uRt1qn1u+JkeC
d/9Ur5U9dmk9i1I5mtzJvL9xYCD98uMhnzE5yR86sZ4VyoXMZ/QFYcnPunqzDH4oWt40o0lounpO
sSz+bLJADKIuzLSatBeQHlDmE4Wnm8y8YDlBbv/hSS2mHQnhmhnYwelq8/AX5+bmaJMFfPHYyx+i
W41ujnC8Lbm3VUG9jNhiAznp8uAiBMx4noH0pXU7TQr/0kTtL8Pi7bLyPBrshYrEHO+G7yJVWxhX
f/IaCa4lhiFdjd0TBjkbAnumQ8pKsj5OqCDoUw16ua/XMTwnu9OGod7oK0C1VQNqoOttCIRv+kLn
g5WD5Y9JLUZb/dinNVtH0/eHKh91eFykEUk7DWTJ/hJ+MxmVu7P0XKvi4OMISyDNMRIOTq8NBN2R
t3iODV843vFSf7N91AS3F8OawxeN6/k7Si2We9zX/Gkuheqik2ii2Fgsz68wouY3EB7+doQwx2tU
tmxZyLwJk1yn/xl7bPbOyrxYV6h/S6n6MaOz9DhpFRpluFAwalO6IoO1s12OtD+iL9JMYILcArem
zhWaKqSXtlOKpOfRpk0ExNFD1+Tdc8LrwN+zjF5bMn1CBNMiCpCugibG5jIC2zwpLcxoAfryjSJp
jKtut9zDh0N9d8oWyrmAtkMx6ypuT646s2eYhePr5JnlmlhuQmi4juXBD4elqrMdP6b1Onu265pf
1N5YUqqRYZi5OA8O2wD8lrONc2p/+HoU8iv3JKyNwjRZAkhJWCkO8Nt3/UEJVCCDr6A6FR2klq+k
STmwSX5ziGR7tZojTnKpUh9YeJgZkwBWAZDM1b8WT35i6bLbrqbkdnyZZhoaEaV7c1oNHD90nIJW
YRH0ZQk4nI6R/4IA9EoNhLE1I2JOb57o8d08WftFvLZX1Nirt4B9+BtT3BsyJs/3ODcVaiM0OEKN
9qWhNkARtE7wqmAXoq/mRs1bU8qXf6bhmlkhIq1oQLNq8hS393BHnkqSoLAjHzhrXC3ua5RiNDA0
jtp+ZnrMfo1PZU4PSi1Axh60rNucGay7qPzuDZ22KUGscBTzMTKO5nRLgS/FjfS2kdpC+1sOgFzq
bsDUeAYK8/Y5LxkL7T1HGokqWqClgEnStPo3c4x4QC4usI3zb1AvPlKsHUafV6l7uXdWQBGuuqtK
hn+gc0o8nd6VSkTfT2K2oGZWY9jaUSkzWtOvIYsFivWSy4FWQKs4ca9JKXkcEedGWkLsO6+QtSqE
IqP+WhChSURNo2X3Ef/ErCMqrN9iUpplUM8UZFuhN4rxi9zejnpCZ0Z2fKYROpsAWJVnXmI5hX9X
I2F5YML+N2EktDualwErZRFVGwdEWZ1QjiNcqAWYZDH6sQHXePY2IHkLED7+BdOn6XLrwcQwkeyN
gCbBysUGc/pU7YxrpssRm1GbGZjvsBxC4AYvkvQfcXuFuLgPRBtaCfHjLVHBMQTq6hWwY93gIaQU
yHxv+vkLWyEKBv9ef2ZR4ATXWbeoG01paCNLplDPz3vpJ09CkcLRIlHda/+gch+QUUZKeZtao1Us
SDR9Z1GhuNPfjlCDzh8K5QHQCJzapJBLkqHTsfNAnE8rH552hItlUOhNOwR9zz4DotBvEyuaIU2b
p1ExzmbEmWjJxTPJ5GdFsP5sZqsYieh2GLJbPvjpIrhh09v6xvgLSLgF6RuudzWdMUXEMbGwdtZO
+r/qnh2RgWN059tF8mhcp8fbCPkTzjDz/CX5pR19N0P3yvMvGsecEE7rYON89uHKSyG/7JKqDW92
WCFBUipGUZpl/n0aklWz05IpKi7xj3mRoeJG0/7D+oSP5L1L7N1n9uqv0v2RPSIh0HsBqlcnCMTm
xX1z1LE1ZlfXAUD1dBjhkrmgYyZ7m2kOF0XKHFo6JhtAn2hP40Mo2JaWCPJWivHNxZnyAJ70xUfa
gEbukNvasNBtLpBN+uo278uM7QUqHV2FqP2j+IzUJi5aY4KTNMc7c5/wzJcppf84+3WuEpww3mQj
lk+PogJNm3YMBZ3BHFR4fQgjPkQHAOBm01KUWwbyuuygk6SFTtDwkaQODkgFOJzLhagOJQNUSlaW
CE3W58hZnNL/aSnTk4mSnnXDxQQOMN1XILCzZwMEZFpGH4+9RN6SbDp0jTAqocqSrMPTCLABLRq0
xsUpdMPzUhHNCJ1PtAsW8eC8KWybUoHPcKUtCpVZPXCOgNGar/KT6DGacP+OGnlbsln3vSVlhGB8
1zHbcwP1RRQPwVAFPLjQx2aSwOL3faU6bRzAsMX1cHbvnoYg/nJ3bGbXACNimdPDhLtD6tOdNcZN
UHtWxQk9uw3jtCqtuUcX0t9McD1En5bwD8QCpDNSxpLsx5SXWZNcQY/2whEamPmf4BzgC/+bYmc5
EBtm00MX2+fqlTOt07VwJuTBguUoKA6ZsGEAxxSRrp/NE6wlXiVxfjATEWciWv0KiuC61ZuasPM1
uacnH+Y3ru4AZ0QDnxjzb0xA8W8YcBq6QxfGSjyNnaV5+RTcBRpLoyelKCswUkrCbG7itsbqIFLP
astCcRjajrL2x4Zgm+yNurfGR8a+FyTVOAztzDTEB7inFNJyObgcCnAankZKC5EXTVJ6vvZDYWuu
nsulpVo9eakAxwny2M8tTQJBdOZEAzvk1+kXtm8big58rYfdcxdl1wi3CLXHSKwSR+y5Fffbac2W
fUG4nZnk58ZRFQ4eh5VSIzW+4d/mTNLz906PYQZ1nVG7WWyhqXwu0Uc7agcqDBtBu1nd4+3+CkCK
mJEpve0vIqZRHAGj55p1bzVeR8OOJOXSFG7k0boVV/9KCDGYX95VOCAD2l3+g0U6aZeha692fG4f
5b8aTX03nJYPop5VkqLlUkyyMRzVG6LxaC/cmM0Jcb3N/Q5Azh5nASELFJRObp4q8Y8u1ntCE1xT
ELx81pnKKzcPmleX2bRqrCfwHdPs5/iR3zOhym/Csdb4OU8C2A4WS306ub73E6jQgBDJkNctvxg+
QQi3ldyxM6J8LNQ+GMJqg8F6TT0IJO5nbnNO8pVeLDcvWXUIitSgjd+cm39H1O3xEDbZXt3U6wHG
Woift/iRhgCs6GbT3nxSEAxtpa9xygLQUbt4GsaCZrvCS/T7bYN074k7U38DUppA9KSzK/s4peDg
CuKDR2xWCdPuuY1Z0kovLkbp8gjJ70RbMcJ0Yla/fNpnGLAJ/0rRI+/ztfylfr7xmAMVhegxr8MA
0cxXycGAfNCRTTC07ch62NlmO4j9IOuS6A/FJqZbN5+oYiydCYaP8nQdDSt/vurE9qsLj2BmLK33
td0lQ59ITh7QoJ+r8ra5lkEemo1+tdRini0SM2a3O69FvPqOkp4CytwWc9uY2ORzEnLoCGqohu4B
oY5xtoKmpEY66WPKx422WrDMa4q6GMNqUHIuiVZl/93jd6ix/H8GGO/g6eb4Ad7DRMI7Rq710WGh
vosFbkKcLkRsFzDxjGBhPa8DyIOziq8BJTkiu2bTGtwgyUvnwxshlWlvVDlsTyb8BSagXfuuzTYu
sZ5BnSn8aMWVLn5SPM7R9WwForVGukDAIgzwbD8Y3B/bWYf7HjA1OivJST21lpMq6GVS0rcf1iCi
inOJVofmBezN81jM/52x/cZVz//qEaj98RQMD9ABzL8igeD1IeoVT9Zeu32aSI+7hO5/8BlUYNOD
2AQT3ol1GALDxOH5q3enJetXiiEUhmt9v1f48dW6hYC9GL7VnMU/BGiHr+dD0yjuCFBmtpad4cc+
C0vvs/dCGv8xPHz8hoyi8Mx5qA6cQWcm+Gpx6ZGcuzGlljtycpixwTuP71riQcenHR3gPbL2HWZx
0UIpQUCfM81WOaXfGL+lmsCS4OVMBLSkmZVyT7r9EmjSoZfRICffivu4DMI7zMoskMV9GPR5Wub5
kfoRvzjQQDeJpN775Ol0LeCOQlC7pPTbEqqdoe5MZYjrjpbwaRkac+z65/PMS7DsJd3Zt5vv8IZX
ri5E6L69GGO/AB3feEYWi8uBhMsA52Vp6itqnK3HgkH9uVEdAqfS/7TOv23a9dnaxL2TUmaNabTu
POwCrDMkyg2gU7LE5P/jpnB7+hmXVxm0gjVw0KOe/HyHG7KD8r3FqOvsHmNgMzYs9KXEIMutdqmT
2YBFqQ99HlXYYhVWXoAE+WDmkJI9tS6sC3xxKMCUjG8uNGRxwGKlMNgSXKGsmAVh+6Aftc1SBnjr
xvE66ZkgQBA92BlOYxrUgBbcc+zIItCaSMW5Kj5ODqaf5VKUXbmRahK/YbT3ElkR9JK77Ff8lsB3
dsVW6p6HvkM/d/u5q0i2uKWkW0qYg8KKbfeod+KRTAknrSdZrpZxI1zkjl9eTvWeZ/1MOo+SRTgr
6PPgXcq1fomkB5Kd3F8LLeJD4qK45uaqahXyCXUvf6DJdeoVj4MywhBmxBsQeK16ltENNAmwWKK1
Jq63Y0bup3o/BX937XFqkPccSVwdbrx5GRPOPX4bS1v+H9je+I0cf8TBxmJnxDLq7vnvYId5/ley
jDlLGhM5PSZNKCIfnqsv20K0wkUhC6ONtzQh651ZXIPHhmWxdNn6Fx7fjr8hdxAmPMpKw86jQ8rK
fZL9TcvRFQXYEt0a5WVpZWlAkbXbV07nzJnNVikUXFJp5h78ddgNtLe1Seg0JNlrJekZ972j/qri
FLi9NcML9klbVFYFXk0obi9pnk+/QZNorDvVYG1bY5wgOWSYbs/e9jIoLeUL8Yw/jItcWj/xiqx1
HywQLkD55VJzS4dwe23X07xPtQo4sYByQpPSR4srlUWsOH6TCAXPwm5uSdTMBQCrxSq7DmjKyfW/
HXvSHGZOAw9JKV8H6zLA9rIePovbEPiTx9r//kpoLOLSEg42+KhX06uUk/etCeBVeXqi7mUzRHUN
fwGfhbjKqH4ynvyHJqcyJRpdXVQnweZqjhx1GdxphcgAqZjzE+sEgsEpQWSOMFCAKkmDaRiRHDP9
7XGL/XtsvHC6jUrbHExWaiZA9/boFgH94Ulixj+eEGw77kiBZvr322B1Dx/zoBRD9PFrdcJcef/B
BHNXVFtSFE2DhpGvXUi6pLH9gLnHe+JZAW4IqX8bxcOIgh+Og+tOc8Rj/jElW52eHmbuR/nO6ce/
f1/Wgz4qAvzOetxnSqhV7ph6RahbF5znZA/UEkfX8Iia1bB6jQ/axgSp7P2xUbJZSebcYPF7dMRH
Ke+YWf/PrRVqdXFH33BxTgKbMj6TCYiDr1iFDgZRpxKkclbEaRbUjRFmIwyb/t9RdO7VuyYlVW8O
nMGDqduhOL6ek2awVWx7G2XZtjau3Zq1McM6TomsEdLBkrfToSsRpbLoi46MMBtzkGNh4FwAw6j6
4kWBa3Ds6P4s+7d9PllnksqXpK34J4+g2XwXxObhhdZ8toC77vBrx+/4Op4FvyijJyhSiQTSjuVs
pjmeWEtg4Cx/9x/o5AOFMoU4v+itUXfq2R2XITbt3ySPZd4+MYJRQgo46lWMnSiz5/Mwp7tYBZzV
fNBjEQGSvbaKjhcxOtM7bZnjRH/3LeMrDRmZSyRslUWih4d6wCw+Vjgk02WVwDmADHRJaklbT1xZ
rJ2xklNkB01E9uEuDfuKC3f/Ocr/EBjLnXjdvfdsn1jF/KB2yab21o9T8DIsG70MUz3BPkgFFIui
XehoS5ibzMFg1tB2UXJ/0S+SnMrXf/7u7PEZhsTpxfBf6Yt/UmWlHiVxt2a9vriHX6z2G5gNvnhr
lL7CGqPEc1NjywK8LnZ78SaMmDbfSk/tGr4I0nas6hB620AV2qRRQTLuPB8PkHCAmC7wHKo2x8B+
EmBMvLV4i54/nkqZsC5+Vmr7p21xhACx4Slk+jahj3zFOLUawII5myEUdzduDPFhCyvuptOrRXGe
mN3lIr5f0vXtGyx5IGdbJs4hxmqwORpcS23QPmEpSxIxOBYxLcKmv50+UPWWl37OQHe4g8MW11s8
6kowVngIasX2344NnQCZ0LD6YXGhFjU7Fm+iCkBbFA/Sk6JvHLE6Ov0uDPVdH97cHPci7U5SZ7o0
jFl/WRj2PrX+kwnT07RuNP6vqU7N9hnFjVTQAf8ns22fI1BRB1fZnHUIn/LZxxEJZ9Hxi2/ZRxq4
rOKZD6zYoeu5+fu+/owBeb3xZTFhiF+r40fSC6Yf95Q1wlvDZp2rkLAZnOpaCG5pJEpblOQhEwS3
vAVIb7QbMtrCPHqPWfXwu4bIFnXXrFyXKSvnV6Siis2ZycuGPVQMZAN+qMRKd9zG9tcAVuQie3qS
uTiVBcsca3qQT4nMtEI78lyazJLFxI+sEgPPc1oWPaWgsNSp6oqzJVp/NbH1jfPJHH9L4EJspHyx
C+UQ74qPUCAEZPAzekz09IH5fe/Ju63rTLyHShtlc3pv4WcHWJy4gqfltEP8soebY4xtAWmE1Loa
2Bt6w5HBFbtD8rAYPg9cVp/EBB+r1EC9a8VqFvMQNBHx+cE1sBpifyzAGzeEF6pTmH96wSD42iNb
KJKWkGRjM5/PoszB4/UN0xjVDP5DROolirTHc5O4Y1JExGeyIa9cLsY6kCegsxjrX0TvI/OJ5Szx
FaW+JdWLgYE3qfxNxHfSchGyvQJWdHNTOpNwQp2nR+/x+CHfzR+4FWp768hVCcAMdaoPDu/1qyG0
0W1nSADmb+WXoTYhc/E7GZEsWXMFB4UcCVLrfdM65ZhYZFELWm5vTnlpltgj5beZFlGIzvkgZDRm
C5qzN0iJxifUgBXmpM3QDhBJ+6kvjffyUjktPM0C1RO+ACHRysLh5w9u/lxRgjwcZolUdNm/bdsC
fmlEsoYTKYgEBeWWgUx4WnoePNaECOZelzy7HO/VIDf9I7zqF6usB+caH+dqL6RwUBOpDGVCE7yE
T4soUXuPX9TEtLAuA+fN6tSmwBRbIvF5svdWn7PnvAdZude02kPOwYpczH1WVoRwEM2+quZpb99k
gAuYm9xQtl506aDcm7S8xCwsBOnOnNmzNTxDKjn41R4pCOVP/cIHtaASgdUfRPBzH+fzhX26dneH
hMQ9MJkeF0cQ1yvIgKlRcjHsZcgZq243alJ012CtiTpIrE0yU1qY+JEGHMoSYcoTV9hBkJgx7nwz
v4i+UJdLmt9M6TQCqMBODGnML0PjdOLhYJPyJZvMyVRNvt+8I49BYA+AJpBUPW9trqpb7eKKwFEd
D0dLOdslYAbXJ/zVDEqjWVoqAeq+NUqlTVeTd9fj6SeMLiucUSHi6sKtRKwqQOb8zPMebtJca0VM
Q8MT5F5r9Rf8XcrMtKZJOKvNRQ0qmTHpHgTH7bXRCwCrAnFia8cwZ4I4LJgLwU9nsDgB6ybZZw2p
p9qsqGDjAlsb6WuNzt9xVhPVIT4g+M8Mdr+vW8MkBBEGSb1KPWb/5V473z7ZvqJGAKbL3p+ecOz0
bbe2bsKitEn0I1VD25bV9ARnsiy4VswRyHXFplAxUMbfyja3SKDlQ8T9iwui/KHdozS1KxozS8RZ
BhKXVDk3UM2grZGZoCya0eI2cJpzHg4jlFgrc+C0z0yJMDnrZ3x+dDid1/wImQxgtY4gNFiJ4Baz
+CkHDbsVSOQluzObaJ5h+SwImZS9OzvAzwim5M6XRd2Hf6sgfYTdgjX1gjNeqMP6hp2P/20j0+Dz
Tee4VGsB67x/N1IjzHzER/T9B7MDNPTufKmEHwIOxKgImEKeGL5rJ0dAEmuPtUfJsjup2v9Jpidv
ZGVxIzDRDyU4XtY5QItJtC0N5cOGOX51nvCbt6P/bOoQchWn2ydtkUmrbrDwy5Ox7IV4gHJgkbVF
KbeAA7rFTsNXAQxhyIBenZ0kW+0PSakDsQFhs+QAYafMpZ16WiA8+wBGY4yZi8L4KrtqGX8GgCTt
//P6LLptyBJLZWYXorz8tL9yAQ8U1Ar/R0dfPfW9VTDjwjW/Ya1ewwLuupHRaHFfGA9d0wqENfUA
EF7OZ9YOuTkVRK/aaFuVHETny7xKEPrPL8RSFvuiBYt7WlX394es1BZfuJlOO5k1KxoJizHu2NTF
k2RzAT/nF1xSqxTgYy7kN2185k0wsiV5MnJ5xDJABu7XLxYIB1nRLD0f8b7pXrqkV5ZbxlHHhvha
RRizFtskYbh+0vB0HpT8tLt/HPm7bdOxqjm/JuGKT+gHzAFCxBHGJ2kfDGc2lCnP563JPQOzHVBn
kdW9pwGEqrXSh/ApR+kUxeIsB56BOr5BjA6XMY/BAGt4YSOBUGcFXzdw7FKYKJaaiziz+r7K9Y0Q
6m2g0BrrnnAKi0/NKj+WxVeObxXgBJy8VPnPy8gyT2PcyUlGX6jS3vebPTBYBVKMy3hCdXN8OXhn
XHTt+krtX/NPOvbkr31P0aFQgyTIGVBT38wjZuAfC0Dw0sO9rsAY3YXalvufyMfdMrSp/KMhQ9gC
pcOOmkV0yCYlv3nq/Qv+YP1EIuUHGOK5H6YEK9Mm7pWzcPm7Hyh4HgTlmnCh91zyzi3jFbwUgRiq
II742ecGJnG0P3WOgfv0WUbZxkPIOpx0x8yx0OBCvtTW9DLWX3mKvMGCsKXopWLMb8tzXSeZYfOs
Z2dfowwvbKYOTt/huGayQtu06VDS5rbJpH51XLs+yJKg4W6qBhtLulSuId2ZQFOP2yyayI1wxsTX
rC2n/+6iMB+S38DrnDLxYg3OqBw0ZYBHxmFKZ3Af1Di1SNcDP0o0RS8pDTUSZbh3byc9Xk+MZjwm
m2K0NeMJffJheBypakrCs0Tvvb1ZvfSU2f/vHSrbcS31JNkyLXPvXvFz/N3WaAz9xqfDgsT/lF54
Ujkq1B8TnmNP5g4wRBhOWqrSdM9yYPVwz5PHNr8+Al5kAZiFv/LSIqcHZgM+qB2xSLKD+p3VbFSu
Qqnq9WolnLxb6gZ3tm0gk7tjh/YpKq/ZJHCKO18J/T8zxI2hVn1W+jJaksb4tD8C+Xg8WOKU0IeM
ZpSeL+21eVXWucLii2sjI7IcbZansLzPVN8Y6Ygb0ZrMFW5uvIty1ed3svLj/YkAqTng14lfsxvE
7FPYiLwzdryDeHTFYph5q9hcZPuDsNt0iaoRuZ6PEtmxGeaNFqN6YNezCwEL3Kg3fTF437RGVfA9
/s3fnSrQI3afwT79b8hmRPrgqCjq5JXDyp4AgJ8J5TRHyqP5gImWTp1xw/+lLApXNfpx5xDovWBB
HqfTkP39asJMpCi1N90nY9IiQTTc+CxoKZPbu1h+4Wdv8p+sAGpAMEP77Hl7nedWlpdAa4xKkEvv
Gf9LOa/JkTIf4/872Ze6VpfzaJkIc8s6owyn4UtmNQh4fyEjTuanCOvH9P4WdN7uMvoVKPb/FeN1
BCPOjiV2hhvsn5kTLipR8rnzx5ZT/aJ5pjuVH9zN7748rxwmbRfxHufhq6Vb8oKDuLD90O+JSIpf
Xf7Kwm4K6hPZts+n4IyOSPByHlDbATb/TPtSsXAWyKxd2iXyh66doJKQI78srsmSr+BFK6J89K7I
K9dfByNudd6Up+vlwtD+C1iWQaFJXjpMZxBc/9JE02u1HaNAkVB9F3haljJU+hWv3GU0mENmsjw+
huGeBGjBagaAY9mpWHsymtv1i97R4Jd9aIOfvK904KHGif0oSm301kvANcnYfbmuE5ikK4OyXK67
LXkvTJwS89zhTd9XpPjD+Ct8R6OGmHr7eCfu6/s2G6TQGHLs/pIQh1SxBBbP7gXXJ5yums33xD3n
+Un+va8GPSDV/cisFVOhhebvgjjwGVcKuRcINTNCo4+iC3O+255lAr4mWAYZek1dc12F0a4SLdjz
LkfRbUc7TENYgPImb3es6x1T0pfJIB8tsWpCB0jI9EwvmwCrIzC2FjtVoSfpXeGgol+SkjJD4jnh
+2zF+zqaoGYxdhhjpBOuntCPsy5kKIqEUYz92nxIijqOzxFpySc7a0UQ65eMuBzAf1c3qxRqXkrl
teWG6yYWRFuDmDyIpMz0LpqO3IPnLg3ujMKu/T7vy97I5wYQcJGqIUCsICU/Rt6q2UxTnCGsAhND
v/0tTXYqkVLbKehHec5htLHlE5X2X5HSx5wcLuUzzkVPTMia3zIJwh5eWR1f6XDHU+rSsp+2/LuF
yQclsfFJN0l/lhmA6/9q1e7RcbDYpNlrJnN04csY83omfnF0gXPj3M4HCc/WTHVp9iQOcIhWjvEG
vS3rf81dEr0DycvUBu8SeYClq0DzgcJpC6oOF62LQIaOC138CQSeEKOoGifu4aIN9hKKpUnRKnbX
ZIBkMCRvFgOhNXBM84/GvaPSnQXkbLvoT2a9qkUwu2ld3Dce0BCZC51Sa+c4u/ULO0RgUye4kK8R
P9I7Uu1gttMEytfspLsOnzLdCB/Oz4h2VKeXHHA2a5XGljHPvkkNaRU5Na3b9IptM8UFyE+5iaWw
aOVz5voPihNeZ4kUTxIbnHWla0sY3TKI+LVnt5y7DLbbQRCLtDRzqqimVvKV261+u6cXuU82H1w4
NJ8Nxq/4KORZj2jwIYr19LDgJ0Qu78XQCu0UIBOyhsq4s+ckMelKPxI1fAppV73EddooyI37DguT
7P2/UxhQ7IrIjMDw+LgjUNozMNfoY21ExPiNc5u67qhqpVSpYaC9LJf/+8IB+29PLgVczREI+WQb
/jMVdKJ1wggVD30mkKTown73nM/uXcvmXp6Pkj71pf2FQwckrj5BIJlLCwIABwoW/GBlPNh7pKp4
qk85oVPtBjUA3HeeTzwXuFx0KVV6VxgPdWelld4XcDIRmCeTk1KHGR8sOCnfRVAvvtfFzf1bTOsz
yTPxyyJymxuXW3sA7f/99VeN9YSzyp3bBhmY1GMOTPc6ar25Jd/NFKf4a5L6kth9WLAhoTW/uu7D
w0qObswrAoozmNvr3QXVyW4We/uWR2M+bkEgpL4NXSVb52URuqJtcNB6JCpMCHgtXAc1HON+8zdx
fp0jxD8uYIe6YiUE4HmytQN1D3hUQWBDWP5LBUmzvyuJEmc3po3o4FPGTgaUAXYcm7KXB5d1IHtS
W/sP3Zqffx0tiIduO+ghovaFfTL5MBRFYrcmddbLNbW8mn9/c+LIxRZxkG+IiEeo/pdVOPgfeIlB
JSP1Rb9XBUGJaicMF6gK7hmj3NBDIKx+zS4EU6JkYa/BQ8i9knWgRYVMl5UzA+CqBGrBWwfC+sFl
dO6CLMXZB8DOxm/SXM+xBnFc6OWKkD5xvvuSrfrSGe2MeR6yefuvN2PFAURudBjFHYOdZDv/5HDk
XibX6ebPsTqF5wWUZZXYBURwm/GNMFKzrIXv7FXEdcWNjFgStW3O6XWpCRhiIaaNjJQrxesw4cB+
XJxkzssXotUDzGDtp+CCo1eQd5c9kTD3jgAy2F3GcOw13eDwsW1cDYiAfJjU9GtTAM/0xG5vsMjr
yRldnReu/yDkW1WZjKzQ/z+nN3wiRXzKf2iTkxAge7iPtWIZm+ZoeR+xBU2srRzYRo4yo8jZoujE
TYZH89oxWPmQ6Qp0NV8cCimSozDCEuJ8+llw/Je545TNfrTLFsxf4FNHkLX+BExxGbRAWu7a6ciH
HHvplw9BI/3SX3t+67s+LoP8MbfSZZiH36td5kCMIikNdEXxjK6ib4BhulXhrUE1124Tz7BCdQvu
hsTx9Z0AJJTlZY7AEuyV7rGnyEbGCyi4tLDOsbAZ95bUFun1JzL7DnQf+nLotN3D0tXmrl90rWK0
bqN3Ke4CDiGqj+ar7wW3RJP4iYggvtgChIxM8wguDpNijCNhEICytM7G+WFok7NM4E5ZZUyzH4F6
vM8n998mOvDvIFOrQ9Wv9/Wgojc7dWKzT4dICJWf2A/VE/uwR+l7oj/1XumhZwR7IuSLcMS2BO2t
lucEoHLVAOId+yG21swiPfx0okQyUZuRqKQ3qnJlnle+DdIAA51idbxOQCDkP0hgGywshyZfCfda
ZuQGZp8wAtWya2PEwBjZVOksd46au5ehqCrkXOU34kpwXAVojCxQeP0snJ2H94LyKtcJcDEjX+W7
fYeLnla0Qeof0ZqGdTUCqn4pAfQg5ZeU5oJabVzYzpAsmkZQf27ROz3DmnCvDNMwsLpfQIWoW0uJ
cCupI63BfCl/ll/tor5tUK3A7AnG/OsvwRlnFf9bj98rD35Uq0aeH7poJL3FEA85DlqtC+aOZFjA
jw7l2TNdMcLAuIQz8uxMBEWQuDIb/Sn2+Dr3fNzqjh5ieOeOZtt9yCdWgpCUZJB6ImM4E175gxts
62mXivM3Bhz3CB1mBj7OItPpk/gmQgk3JC2GItEltvTCJ5HF1QzKfXFpdxm4ctkBqJab1uElvpAr
6Eb3SGz3aOjH5BqJ2pzfCdqPfaJIfKXh2QkD29uQnfEyPLiKhu2Wy79kXtJd4QEeWJqbNguXavPW
kv4CIGRdaIoB/Nuu8bZSWBJMoVDMvUzdGIN0C/58aYgxa5Athi78TL1MktIUIvgRN/ED1NqR+E0/
wU+fhzGMrWwapADvWSJAjbnkQbTV62XbitNeBvO3h8pIUFZZhN7kZ8800KUnUwbzcqVXbDvMzPMC
hTroWqUWhNhYN4O/VzR/aBitf69velRqUU/V8X11xKExpumCsQNyZpQCqnCSm2RNIrp/zByCNKuE
sHmTOvs7K/W68F0PbQ6qKIsJSQNmSBCKa8hVPhXieCL/CIkr/Fm42+YnkPEsVusUQmvlyBEnvlys
hd5V5TB4Us98zhCvJ5Z9XvDY/9t1FxTdjYnOGnbVybJ273zJZy0aUPjIu1Bf9Hx3rRIzVyMN+A8C
2Wc6Cd6wpyMA+KTQ2N+KcODXx7e/Sax2+mkfy98ID6mNZQEOvaVC/Q1gmZNegI/6Hz7PD/eKHeD+
BYcCabkH+nI1HUQA4j4wV6kGIcxn9uNQzzhuGjC/KIq0Au7RcECII/qxBd6f38rrcyvYS9TPQFsu
pYn5sZcya4NbPjvEpm72dAeFquJrOCXyMbp+Q5hqDKhRdeWOkLLUNXSizbO7VA8t+GmuMhOYfm3s
mi/w88KBoHnxSxeaafnBX5Oy7FouBBd1v7g0PWzbOcxtbD8XFLeWkG5kguyEh8D6+xOqMn88p5EM
oWObYFI3aQQnTJMw0IF2VonkdbO7r/EFSGdLHHcXsYGzpmmV0lTc/9c4Kwq+W0M9JkY+4YA2jVW4
6SQrt6Loc9qF1U1Ao0AUIIN0/JkQgoUsUFBC7NomsQmOQSHjT3GWmDdBj61DRAb4/CdRpDwsXDm3
8sCzCzD082PR1h8peSsrH9Eea5/oG2ZvuGfrn5gu1veiWxZgQraUDxaLizjwvY7zbxLntvVevtCe
dwNn2S14asWmTYYVUaK3v16us7/d3pOlzSVEljsoVpNSWfMYMGkcHNRncHyZ9XxgoX3tMRUYmIZj
CTDCihY43Hhkoyhe5kI5X6NW0hLVgij1yl8ZVH4I3J0XyT1CEI0CcXMD3azbxS/EX0NsBhRuOIeL
uMQj1OSn0i3PSYnZFG8TKhltbkkchRehJF/qVOa/BLN0uBHtXw0mT2IMkkav/0QsfRzWU0uOW13l
AeR5y7RTX6j/mh579qg7i4vB6rEzQ9OO9Vmgy9zbRUrQcUrpdpqO1/Xs0IBfGl+B6u89bBk12Kj3
z6gJ4LlDlcqTK/u0QtfiMaaJwDgh8HjudDndTuToYeSSnwel42zQoHhoBaUAUJgZZuB5rrzLuf3K
FLaRz4jo5MibKYMAge+QLgxgHRqXehaMqV70gsZu1jJiwyGE4h3nOlciSjpMtkL3RbbDfPZu7AZs
Ixs1XcjEOmeL2NKv+aMnOwH4xsXXDY3zXFy0UXq1W3+MJ9FIsrOTm6TNiZVyrep2WDFU/zDlCOep
iAXToZg/EMgY0YQTGudTDZ67fzfLMd03TQIR2p2G0JcQmLFVBiK2/LgMmqNUCqs8svJbKzJ8qpJ/
4fasC1YdWGDeA/FpuD5HJgppvhL1B40mdrVDBCHwpz5x5IQwmzHkMOP5ay7z0Y7VJdbH9ANtaOko
eOF09lSJ8DCEQ1YnvziTCJROfc8avhV2468aXmRuBCaWNr9VzCXQ3e+ggmu/T1CnnI52sayGH7SC
0/AdHTp3AvwGQ7A49GsfvifxChiLgAwDDJmvbXeL++X/dYNTSRotRDsCfXcQ7H1flpPCbnXORtpI
PgyNcJc/E8VJnzdJYof37cEVt13pVPsSHWCH7S4if27rVF1VYH+dQ0zZklHbblSxFOKN9FBWPXgH
/l8XgfQoYh6F+CLXlBQKZQ3EX91gHeOgMt5aks4GWCB7z6a0GWwUyE2rFog+tl8ejGM0L02Xx6jx
AJ1+1zZ2g6u0K6ScGLS4Y/nBk2H6LK1FkO45VTMkEJoQbFGUIX6QM4ujZFbLplPqVXohCkRmE6WD
82HtmUx1h2hJbGkWcqxid6UAyN+AEudEE1Y59lf4YhWN4gYbP9krHK8IxlWF+8h+/UAfebZoA6oP
kWVFt83qfNLlvyg7nECntQRThiz/riYJ71TdIRwp3L0mQTRqhPY8Jj3xzcdprJVNsbKGqbsiKYRh
wl4tI9XSlmgYY3Bn8Skm7Kb2HDmsscvyveCY8QGei3TptzmatEOX4r4Kim2tksTWJn9Ox0NEe/oh
MjTy0HhKxT2NPDFZEdiwBuDTNjI3k7fErx8aN6DO2KCMZ3YgrSWNQOA7UT1Cuc05S+Kz4Dzzfpg1
T7w51sB+CqKF9fuXUWoFpYUNcUutVjmG5Lj514/C59DFgFjjLvMIWYTfOa6Vh6cVpH0Qwvyu37Pd
LNRDu5irKJNxp1TYC82ekU0gHS73XbrlK4Dn6yWG4uh6LjPvqQH6sA4WUzILkTYAQ4h9082mO/w+
mBv8m3Tz8I6CHvbnpwUhX7KJ9Z9EVTCPk7Yqz4CUxYzy6GIaEOm46THbrobvo4DREmWGJ9FBBtDy
B4Zmahq5laPRqNHWzVWClDMhbNCBIv8K+mOKYwHHm1gUG/US5iezC5sgKvZUsaGhMKF/+ucfjVyQ
OKRLZzBG35mOSBArSc3BAuIKw3B6ie2MHyWwcvCxqXUi/rw+2DUetj9FqweaE15fMAiAtJHDBnnw
dNzDZJ0nKH55a/cYK1bWZt3iTyvKdtXDn0NvIsINLdgGXZcYhOqvDnzb096HdS18b3FOw3lQy8R8
XzSe4yCDU5kjanYXX7s4/4P9n7NZ3IfdqNNwJBB92dLBjT61WwWdPRYyJTnlfOG5l9UnPJpOMDyM
+wSnwpNVxvYbydq3/MaJLkntf3FdUzb165tFm+9gbf5gD05Pyme9IW689Z1XwEbo2LGM29TXs+zC
0j3T6/jI09nW2tR7NFkvPRTo027fRYvmOtk4wCbmdN5HLuzZC7wwbP9KuShOFGTj6Lvo4R4EsJl4
45Nz8oayH0L39XpsJgLZyGntRL3X0atesdBRWH1dd+JA3/jeDDxlHard62YVshC57zf2wDBxnR2Q
qgyKXTgba9So6kJyVjswV15Id1hiekT6Hcr9M7XiyrUwXG+1s6HLUZOe6XoI+yuK/xfRtAt/lshH
h3M3J//Ffw15b8mom0JT3ISi8Q5t8eVP8+UCUTQkbGmy9ogSV/z+Ll1+C8HFK0IBsmIGsU5n51ny
MAXSJUVxJC3U0cycsMx7c0PBhzEHS8vjnA6mHeTVP268MJ5clhnGImQDS7+MzVpaW6NVwf4xhKzX
oszvBfbBHfEm0XIyRW4/A/OTiP246V8wLisKxBF+gmsW0w+/T5zwedIXypP65lkdjjRWjRyn6hQb
PpK2z/kEujB6x4v6Y7T/b873WjZ9LtQ61P7lAH2IKcTIfqsi67GJB1f1CqaBCebTDWlZploa16nu
2PJqzXOexsOS09gGdAs2nj5IBaWrpU0ocwc3EHxRtnifPHPIzTyo13sTuf7lMu5dP4tCWrMsBoxN
MDMipU1LJE2nhn0BBMA408JBOnyFo98iFP95t6m+Jl4/gbl65WEyJxhZxLfM1l4zuBnYE5kFDReR
NJEjO/PpvzSACTNo2rtytiNVRSn8uqviWHT6PdacqgEG1e25gyQQ0j2TtLubU8+Q3mwDRrIuf93f
sYKTKnqZymkecBx7wfpUnEM3ZJ/tSdcWSB6JMRm+p2jAcbZTXtg1JoteqXVunDjOJF7+KqR4Ppy+
Wu+3FYJJ81Fv6HyqbJ6GfAkS0r/oiB1rP4VoPt7YSlV9gBVU1Kr02zeCQiagZpAMv9Wzl0GvW17A
yCGvre+YIDzlCxKfK2rZ0yL8PtX6/j0DAq4k8X0hzNdeAxk6ihmscWLJIQzsysi2RqC7RDxpy7Es
/tO1HevAikxyOOQPmYP47yPjUVam9Rz8eQkUiDKskqidco6UXbZzFJKk7w5XUzMdLOArOMKdx6AM
a8QuF1DL8C2B7hKeC/gMPQTz3cbXScTs5z+iF0/ekiTXYfAaPoGPQIB58OSfHMpKoP09dSq3HFVL
HEJd1FQ+xr0/ThF1vJxEt3OexECH/Z/JMTrio9/V2lP1bmug938TjIDTcZOvFS6nKcm6Vpj2e+HG
QwaIiOSUEDTAtIZIBXVN6e7mktxmDsl8MC3bM5ZFeXLOzFeCuVsDeOZDaE2FrU4iTovOFkJO1r6M
szZha9hX+MXvBtm8L6IHWERHJScsfrasHe1lEeIu5nyCy6XpVS+71POS2wtdK2INH4BY9hcgbP3R
16OBhQ7rI/qdT+MwxgmoEon3nZvfYZATkLB6T6kWvqnJH5f5By6gFxa2lb6NSNGIl+yRkHM0QNh+
TzLZMBjVJyVXq9hhAFYFSRwrWqd9bSloJ897TBsH1Pz5bjIRBsHL+/J604Vizy6xS8NKxutwhrBG
YKLxlHlit1YCiQEovjQ7WhxCpP1nvNFbYHNzo9UfL+7bm/SF4/awt/CHi7HNjTX00pR/XZI+EWE3
VbXt1LvvGEdDKep0WXoP7pGaD40l/4eN+uNWDmsgZFBHJ4tCGJtR39Qv5cv6PLtpxyp72ke0jTCE
6HmpGUXCxCt+lfZNmGH5ugSlN4OV+La2lv8M13ABGuXSnlcNW31NRGD6Pe+q4gj+eshaNK+dzwyz
2at5SA2+2BRkjSqOZMb1QRBTJcG0eRialpYak7snFyTdLa0Jss5MxgZW0MF69sbcZcWmgvjVNMaI
jLZgJxPSzXKLA04NP92uksI+0JS5x7xCqc6j415LO3asmcA/+/KOpytsLjyz7UuG1DVxxoKSzo1i
bzHLanVW23tmH93To77HCVIES7xJLPYWpKUPe+hl05vNINzxb1blmDW5FFS9KqPnbFD35bW8L+6g
JlwUooebj+ThOKiTIB+YIdWOrOZzIuRxoD3nf8XpKIB4bkzzM4+mtd3amc5O3WVMGMNutVzx6W+I
0Lur9nty4CmXNZuyPNnwsOQS7AcLWA7mbkXGxTh74Q4j7bliKBj779h7dWCQP1LPaVJBhG4JMQZU
hAVXx1OB1DibsbNDp6fNYBsAA4ZL5IjcObc9m2J8dyJ51t5tMIZhQfOaOz/6xuYXLgURckV5Fnxn
+WXipfsuXR8jg51FMwaXG+SSycyL+cuhiSxYo/wb8dFdFPV4DZDFGl5iImjRCFGWtSC9TZLhoACG
Zd9w2KgHubSHFw3+H3JaxSdmnKcALYa0iv0VJN+uszPDIHN8MG0fKk6ufa4kRpFrIAT8/aPZYFfb
e+YCp4WG/daK2ZcMWV5aFR2fJVroJoLDcr+4wtgBryEUTKrzu3vA7kzt668SiJVDChFq+mmTvLn9
4+mAKIKnqgQ0ivCrt1auKrlf3WnFpQwtzjUTS1eNSp1vQaLZ84PQXFjaAIkV/Tl6zgJj+u6Ak0Bt
E/EPPdqa9Xf3blo8NCmLFWyk9GQ6bXOnH69A41WE6/caapKd2x73V4k5WGwxgHm57AVDBO0dQXJi
x59g77u+vYN6X2aAHlAdiuVX1dieZ2FSCtZJhN1zWPSpui9VYJzoUlv1AJBZgT87h4etU93hpLZz
EinHVfNWB4G+8+x4bmry+qJzALzwWT8c+4i/OGfG2zF0o6it5tRks7eqZLoAfqKcPZpN5xE81QT0
lIV24JtgPnu/WiGSCyMmzX2NfscybZozs55QniiNxG813FpHiSLM3Am9mMt3vMiB7vG+NeStc9KH
SXSjiHbTYiAEhWbx5Q7jpdJ3SwGlBAsuvyizse9T0PY/lMcwGnH9Ed/rEC4oGR6XCaJKKVBOle8c
9yxIw3fQbwjNN7WGeRzx/O+H75ut6pkBG+z3aoOh+Nw11wchn5WN0FEd+chIA4BgRe4n5Io/lhRo
1u7Vm70qkEuRNfhNvUjDpoDR9zv5FSXP4FDSClzcVDFxgiYjkq1Kh2iNtH8oJhb2SBC6FyFb9/Qe
GGqMHDM1VX5Ge519+hYP9AMv2jF2ZvQp4FkEnHuA6Uj2c/SF/oY0E96bRWFvrjWMG+wddPEUt2fg
J896BiKb6K5VwfOZd3S5ftLTHcjiRRj5utTdZTQtRwHkkbfUi/7VNjnM9fddOf+cugu6YU4spZs4
7lesF4xeRHhCoe02XJCMR+z0hReOng7aFnvTWAqnpmbd1vZRuIehgerbAyMVBiHzyJ8NZGXVNGsI
kVABsoarKoLCFmHs5cpO7onXhV4QoAApUgmflv7xJsYBdX4YGxMbteuwkllkurLLhWk/cJ9d4YfC
W8cfqqfZRTe+kti9pkeFkRF42+dHCQdFu69ZkNy9ftyXbjuKHjs1WBgqdVVBlRIGA3bersF1Gcmw
A8iB9p/Dst9fRxsXGnk4t+P26nol3cNW5glVHTB2WNRORb1xHHwmoY+VxgIRNiAFGP5XzevTQj+p
PXln99c/bfBTyz4Vop2fgDhxJdA30YeAuPc9qS6LNsQWRF4euRST8nbKSVA3XfQmI2PiZP0UQhSK
i1LGV7rpWWWEifBDsaD0LTGX6y56GT/7v5FDrE+RPe9HvTWIvFMq2bJ6tcHfO/x2JijHVsXkblBV
Ren2XpLTdCAuhpDW/UVH8wKnuK+R0CfSeuIwCHoMzPxiRajb6Fn0OK+R+9quBuY11e75y5PKzne+
upOU3XF6/s0PVMim2l/me8CWF8o2UT29n3lukz83M4omzu7JMq0vvWriqRcyDW4/jBUdG2YKLLq1
seuciFeiuRISwIn56Kt2XmFg1Zx8E8Vh2rjoFkaikavsHxFDy6GGV1Vt+wApY68vQxaj4JjEnwvD
iByvWeRt4ateWBN7D6gHjzui6wauQ6e41WR6InQZHFJa+M0mYeHeMCVF/rYL5lrzjRQfYWoDtQhJ
pAZv5JTDT6fw2XYIY0pYbd3nMLv/946+xcHQHCTBcTktz/HZTzihH6FDbK6xlDdA1Je58QMImcsi
eMf8IFQNFRPcNjfoC6wnunidf5wqHUuMjn5jzjeOB5iNicdpRuGTnEqeOsLagtVgMwurnocarwnS
t2ip34shnDRMMFeoenn4PAJ7xoSlh0TjUBhIJ3MTojjIxcYJHOZ4zhzfrbLMFq/emFg7AiYK8eph
g27FU2IAEMoXNt1jm8L47cXMgyNSY3xqlFSg9/pW5XuRVvc0pAwcNoYc9k8nMeyABhrvDr3NA4FF
EWWNXrA4tEkejqQCgY7uD0iSagMtgbLr4TL4vD4LiINDrD1a9J0/u8jXWKRtEUrrq7hl1O6dZFNa
nh7tO9fVIYGV9oleKY+xETVrNuR+ElfuwWmo5ZjGDUWdN548ihW4CUYgzV1US5jmAwI19Uxi70UX
KOxWlm+uvBrvOeywbchbP+Fxm7n5qzi+YdX+thoyDqZsSTeFHXEokMli9paXhT/N6dux+3CPYYzU
N2g1y6Kw5jNA1JpYZRQG93wDAwLR8Tm5W5p+nBgm3GPaueuZq4vL8N/DTNZ5ijaCcaqFBsyklm9N
Zj9DCjqiLHVWDqLy2KMCCAtTS1s6Je+mXRAPn/Tc5ObZ4FgRzYSFfH2P7VpeBNnV7eSqjOr5W3QV
rNyJQ4MLNSnE2jXzmRaqlqlnhiB6UCabpyYQ1QxeQoqnKPWsXAslVwbmO1Lm60kJc0MXgxTlZDNX
arX0yKhCsx5OyTRp5SGkqTGRols+/LPaocg06DBCcHqxWKOkn/Srn1cnotsRMWqIyCaCcA29QSQ9
ALaRzlRyJzWApQJhCfeYB33qg6G01NZGk8te6/BU1OfPm2NYuDVS44ogwcy8rRUUnRjPf8ZHy87u
rdQYyYdcpPZiaKqeV+I8NkQbC3g14p28sY3NmkzKGA7OzgmiFuQdi4WyjH2OBt/hr1m5BDbWk7s3
qEjyNHVts5IERa+b1THXXYfjE3RorDMemIJuUnYeGiQ8mW/tN9oUE9bkOuEaOofcjZU8j/LC0B68
C45B5UumIGPddeBQFvji0RVJ9prJXls1vnJSwmMM3Ve/oEdPceXH2jndy3UC2gbEcq3kVKCOxka8
TK6l1FQw5BTOsFFdnNbYWMCyN54m4bRxnDk2nQluaGVCPA/ZU2zJ5dWJHX+IWOfVpITTvGqH2uP8
4rwYjVA5G6EqZmotvsBv3yH5Ay9Egx+1y0bDil4PRiLmJmg9Tf2VRXcmm836XQBcTnLMDMbJb9tm
LE2m9FxWKWCTbeBZ2b/BIOq8acAhxKmUa6Z8akpMVeeLHI6hByr5/645WosemMzz4/rHFzyzZddX
ELmYnfLCVaRS8nCWTUYxpkNfWTbehbUtQyYisxb4n/JCMZD4QKeK8t9L/QhixQKk4EXBsJEDgpqK
jPw+syK6DqEvlXqe9gBg9Kf5M1WHYC6bs/9+uCYky/c9mqpd0MZZej1pXtueHBM799pJcxt4LjLf
ar1NlhXNDfUokDfZ6Azibpb18YxHwy7rZ00brQ3hW9t+qppOwyQLsM43AraD0uVDX4snm3oWX7hq
+wdcTpHaZiFNCzVKuiasL09taCkbSGoSA/s1WzosxtNZMKK9/3i/rSusAlAhXp8HssqMXRMok3IR
5OAEsgw5n+anAreglePR/2glkyv10HevNGWBlN35sURkQBY9q1SozyvK/DMUTgSflwiHtBl120FW
hPTfLEE0A6z9nnvjfvGrx/BCWdHD2kC+FLBW7AXF+55Q8QBA3ymvsp+z9rNyNZPa74zz6Skin5SE
FLth3oSQvLZ+hXu+Ab33CRFa3as4rBSiscOq2zFWc1HMZwSV1uX+B32Pm9PtU/NYIBBZMf1JdMvG
F1wx9+x6CFeSS6hRqcBw/cZ0vnWhGdblh52VomH0JV8YS2Nan6iMO7ISzPt9PxW15rXQ4tV+BQb9
x5/92iD5Q0y8o7xVODUULqFrFkYvzcncrejDOaUGqZJrwCsNn9YCkU0ttlIg6TPUmp/czmHtGQCc
cBZQAFFhRiVZgQHceb9KL9JyHDq3LE0Upd2BZEEXcr57kItoH5sq/z0MTFk4zoxxevY3FUDiH5fY
14oQfKUo+TwzFcP1eFJQbkkxAVpx9m8HIZnl/2xvBn4jpPgnxBBeqpI0r338/DUM6km3XXuTmnGy
NwWo9qR/xVckdjYVP/FcYXvYeZu2vtTS+bAGkK5AwkXdlxxct231Nb3yFnMJ9cuTmVEqGYkw6akV
jUWGwUDXHvS+uF7J3HDPn/wwMsk3j85klT9bRQ2xdD4zli4aKg4GFi5NdpOdAfgoJa1VSLIurn1E
BGgc5bSisga82xB45sdGPgBkh/1PnOuocSPkfqFE7D3Ge/knd9K1qxQ7mM+skOwZSEcQk3/p9emm
GOy3yKCKXzirnCdmRd/RZ1tArndh2QvNHIVso0r4zLn6Uljna6GBft0l/IHPuyyKnD9vyciXjSho
EBHHp+f/ey+5JcKxHdsuN8y0dHT/5MYsI2iCG9zOkC5W3p7PpxoXpv961w0oK1gV5dBFbVb9VsOl
CHQZW56IgjcFUtiUj9jNK4xFKPAigm/bmbsIywz/pXr9PEcVlN33Rp5zDol+bDtV3P7Bd7RSb9zi
YI5kXo7WM+SkeEFny5ELtk0WlVYspENTW3Un/xJ9TDrE/A0+MsOwRCxoBJdjsEoiMy53ag9e2s3V
7fUYZW+CxMjeDA6QSk4ScMmdicPktBfV9nv6IBvNy8CTmH2Js86AkVfPe2PstUBADGMauW09yajl
7/55kRPet2fdjzvHOALITrBttgEzsw+Fke77+NSOIM9khB8zR7q7N4BRjWYTYqIJdT9exdJ9YAkf
QFiFoluerhLkMnlrpxOjkOrENiiWOXn3faINqjGuwxNscd+apsg1IrNuQ/CQfZFA5K++icmziStm
VCsAUg/j6V1h1y7fe0H/XKzqtWL3RLPJ6m7TiFFbwaMTfi7G6EFpxtsk2f5c56osoWg7kR2BcoZx
/olz3FCnhl+fNU9HkHTEumFQ0mvlkSk+pwWooMql2Ge6oql34yWsUJgQi4BJRt5ALOvTNJCBUb5U
xEi1pCl/Qg8ui8zHWybKGIogav3ElsUJLJ30ER8+egh+0pPVM0CR63XmZbqjqvZ/uYpdILvEDxam
O2JIDnwk97EUjqpyT9ke06R6+IVi+1KzDKl/OkQlaDZRk5CdKhS6AMERErIFcn8gZ7uDGEQGI4eA
WzQre3iCGgTs5h8rZnIChqVQAFWYG1BO8qZSR2y+MA5hFF6eGs3z2LdOxt+8bvKYF358GLTfBhS+
rDyb5pxDtsuafBoeNMh10d/rOgtf1JodHKH3IqpLkF1juGWPbID3Gqt4DgnD10gYlQghVSYSDPpJ
966hI1MKy0ULrZbnBXqzZj3e1/PJgLvbOLGIa+s054GpBMPvkREh3bfNUruJ8PiOBz519nMnOj1f
maE7teiaylWgmADnfG+RCD7YsP/8I/UVe+cctKFdk7ZWzAh0kBiRysY8WptPw1M+heNEVo/rfgOf
8OUA7qVFCNxC0bZ75Gu1NREYZ+h3qxeYpE8l6NiT+0dXovJw1sJxe3Ln5tTpQlo8FpXHg6vh09Li
Kf0iUgQG+2Qig1KWKymAWNTXNx4QAzwP4umklQrwXYCeIGIkGA3HrtqTizpEPXTCDdLOSPUYWGYp
FlDMuvFHCLyAkG8lOZPXaATe4DKWR87pT8ddKtZx0Obv7rGLBKLaK4TjyLQOfBZvcCmtNTruWotE
xmXUnf7hULDdQGaQuZfqh5MN1FYVqtVHx7bvKnWj4EmmwYqc/YV+mxY6A8gZH2UN/o5SUnbZIKR1
D8udxrq4diuKt1I3w/gRN1ZiiQ6EjKSli5BRG+uoC8SzYaM1MncNrIEvGg6hp7Srf3c9xEHqhW1m
/IlLKhaMB6nuo8u243zDOjiePwj/izfdJlfGUNL+mzEO1v8b7UJFqWvNEO1gTr34Q5YUx1+fWKXT
99gga5WFJlcXO2fGBwZkeiu6w8NNSca1HmHeMNLBTcAhIvejFDwtzjxZprEe1rQ62G/Pmv84MG9F
mdpTKNn7kZeOQNbQ6Y4k8wPIs/zIm6NNXEZyupuJKQlYGRLe7X+Vgi0lMd8DBVBmL2VL1n3O1Hsv
EbKTLth/ke5r8D1WesIaICebdqrIA9uQc5WFDDjBtnwD29b8//qLFXWBusbCZ6wKGE4ysH2EteEv
P99mCLbQLf4O2d84LS3eNl3hQDxqSUv3xx9AJD4AzAP9Evua9k3qSvk+pOtfk3uFAo02kapdmqqI
z3cXltIasVVkl/1YLfWhKfSOPj/eqAGd+urgPmuzyHOYuZDYk/KpOqNzNSR4Z/JsayhXmiv0JsZL
Il3SM02EbANFzUZtGytHO25ZXF2+k9DthtMwpYGzbR3KSPtaK16RWi7KZDbdXMMQgYEcNisPR1G6
jDStZ9mMEQzZxBjbqAQBXsnDBWzQnBk2SkGcfdP3WwtjHsSk0eCMTkZwan2lK1gHWgIWC07W0uHl
uK63JIfAl9qK16QNP/xl5bNfoswsT633K1E0llKiJ+PHuINdmHfDq50rCHVH2Q+6soXnBOlaBdke
8ZN+AVR1sk7e9eGZ5byQC6d5bWe6lLYUb6HWVmSmnzHGKMl0usyagsXWxiXb7HWU0HydnV3kEdlO
yxCbX9c7IXtXQ3xEo3gEgN59rwJg/mlW8IyTt3fnVJE4eTAD7pQhUDMw1HCRR6jysajs0MbD3GDt
XJbAYLF+J2muqeZ3QsplToB1VbBVSbrQOmHnwviJJF+Ls82JYuKOW/hJwsUoBWU442O6Q0Vtxfkd
M6JvyIytFCVecu2/G7d/7JOLlgR5tnTNKyVq8HNDDYYAXlA9tjXW0qhSJv+w/8QI8tKUoZSKjmvQ
ZTZQj2KZJumMvKG5VWa9g7ka8IhdhYpViLoiP6a2u7+yDA3pSbnGUFbt9yDmlmxmXCfYsfoTb9bN
l9IKxLNwo5G9q9SLQyKgi1j5alXKZ325P7BaJHR0Ctq2GEwkBXBTXl35fX1Uv9v2gcacH9gjwXdd
FfAEAlvooEOHuLVRm2HeViuV9TvgRntUB9lEOkHNevOXFoYP3m1H+y0OCzM78aa79IIHhrxOtNxt
9agLNjywe4HJ2a0aL7TKr+u65ztV0tfMoFgYqSebBnJRwyQiWdWO7Cdk3E0ps3uL2jvr0M2E6DfQ
zWnYN53TXYesrbiDrJK6zFz/YzR44RQmUjy0KlwI9Z3tcm/G+rlrWIJab2qRfLOPMYrkfZsLlA7R
MwHZYKKOjrOBtXYlvqRyPsxR+7e5ger22iM5YzpRxhgwgNAOr3EkGy/XHU2nS594qPwUTztSY2/Q
KlCyFFoqjxPm0AOT/30cqEPkcpm2y8jqwoAAdPZwo5QKWuayvh7LGFgM35k8zFvIIUFWWneFvQ7I
dJ2kE5fJ8yL/+h0Ugx27SXDjEOTQVIyEwOwfmoeeS55qMgnC/q+YNqO2yydmA8tn6cgHrNJd+k84
eC7Dq40ukNWDppP8owc/Kr7D27QEzoJAHoP2vtU9RNuNEcGaNUTTlgoR8Vn4HnsvPb7K4thzyD93
pT4sYoIgyqyxt8+4cR0SI/QLXyFBlL8I3TLUaOdKom05aLrTyxO6qFgtyM4Nonz3l9eLD8qr8wRw
UzebNMGVFrRP37qylHK/SjjMkjc4Fn4QCXaELsI1KksXhzQmABvtOA+WnBYlnqjjZSiWaSLP+dVz
OF8Ph8ecPXyZGqSeKj59rYb1k4EEJuMaafK1yUrz20fdNHRwcg963gg+1M4OzSKPQiNhP06POzrh
25YgVC1OjRJ40IHE9Ek++UFhSKcDKh4tj/iaJUs5NYS4gwHOyDw0USGRiNJGS7iRn4lRVKymh5oY
d2favdBh970WMGMM2le/4y3yQTc9knrC0ykj/a3eGykP8cZBxezbXFvUoGjq4YiaGUBz6qFVe+oU
v5/n9NdjyfzSSqaMbrzkuUazg6cbJt41jQz1bsYNDDTQNHYVyK3RRx/z34KZ7riTMyUpRZvFdLcj
yQdk2Fb2oTo9ewhxLZit3bD0gDyCgCJOStgQkZi2/OVoj6daXehhfeBWuAbp8cC+A7Ga91zNjcYS
vn59gVfEJB2+57bD9LE6lmu9SOHqK9Njkc8FSV4Jih8AL46V9i/kW5wijPN6CT5liOVSLwNQr81r
hAhKLxQDQTQPF07Yt54GUuFg4V03HaqGc66WmWDwokphfemgddg+rRvollsg0aH9SgCjlJhTmi+6
rXMxJSLLFD4etqR2KEifomHhRwcU1dSQ/rfGE2+sfG9CP8FaLPIiNoFA5mgG134NpxAwBm8rYHZI
Cdt5NMK+PDWD8o0pk/bcYzVLZo/iXRFX7joAJnorhPoUWJUcmeka7fnHNhFcfTShxvVzXJ1djwDA
1NbLATpx/+Iwhq54AN455zoIuHWhK4qCZ9i/JPE5Q5y2lQwah5aQ8ZXShIT45OvjxmGkqXKgaDPa
nloZB7GBh0BBtsVvNOfwCQgEpIoPf/u5S5EQTaov5qJ2/8ob/XwpZu0eMgdI11GW5Ivxb/SdqRB9
tX8uFVkBPbk9uapkQbAMrCB1JTv+OBHSm7pilQQ9LEpUSp+RjngtRNr2oP3Xq7QW/GL8Xt1ZS+uz
ZXD7oD/LpS/6Y8dtJQsGLiujSm/dTgMbwo59Iz7JE42HgIS1Z8rLvfRop+BvMV9qnmwfQRc9nlP0
gZPDgcDza2j6PZwPdo8ewSxg6vvJNIemPkQ0+mkeDxcBASpLnX37RyobwpTz9NbusSXrzdEbwz+n
uvOM0qTMMuZ0aDTeru9hw2dmLk2bCjFnMhI1gT6gcsTnUv3WqbiYM3E0gEPU+TL9HX9zuPljGYbR
toDW7BoBmhYxdvirnebfbPM4LkmU1eb2ketJxWzuFG3KdiywgFU51oGyZRWMhjqWqW+8Qt+IwcPy
rKjlUyx1I+/TS8hOtYAFf0rFFUAO5VYA4kUZveL++R1qn3MamwBGGDn5Cn1teusb2Zz7/OEUrJo2
KfTTJgQ9fQ634Idp67AYjvb0l49maCUsTzfPK4qbh6y/NA8N8d9HoKUSwZDl4Lbhidk89BHy/5vL
R0kXyUQnvj77+seEbcY3BFoil3bg01CgDypYixR05NoioJ2ct52Cyx5XNdh3RdYUu8UFSGnEy9P3
bUh8pkUmm0yqIPzJ0LAWpZMT+El64qTiwRgSP0OC8yCPwgy6GBBtU+i4KLgpbIufvEjltdKrDeGO
3IYaEMrppvx146PEcM0H8BNL0vX4FKr627hyEbZWm8WIoL6kn+onKvhZRu7+77rLP+ORB80ODdYO
BtQeOWbchJJfagPej6GRO9+IdAcNpdINBBfwzp9F8kTAMEH0bzwafLLm8NcXEQ0wBFDOICwaCoKo
SlmrD0lxBcZUKskmEkjK3yPPovhdGoei5s2BUw8pbD+jfppiuKdY8eYtG8y6NPy294hQWGY7v13Z
RusEPi0Mhud8abDLcPTwTEuUjBjlv2jNOgAYgqhkxG6aogYQzSTGh3w0mko77eD3ZXk4DdxzfJNX
EQ1+itkrI/3aDWh7MXjBw5V6gKsuJdTHEGkrx4P3oY3do/9XHtphqsS17+3Z2fRp9oMEKd0EHFPu
/L52bf3TIzaJG80OWJK/oGJbXSR/86a5bRCKoZiVXLbReW3yI77in13gDJeDBFBEmVyj70CJy/O9
PV9AozeRpu5lHUCzNqcR35klt55/lkxC8e38WsArcKvVk1ctZTe44GB4y73HhDrFPKXeQQhpXY28
Meh7IuNIrzQeDvSO73qYVV+moalZZDjEFDvnxkaa0JO9Sm8i7RYGwMxbOkagXuLhZEl++LkIFo3o
NOiCe4O+o7mCUZLJzjyMuCuMdDszuseJBCjtb0PbpawUn/ALGpjycHY+eS52h6jJOG10fVwAqIpF
eIwFsrUTW2XtpJSiRW1f8p3IZDD5MTNKR0tK3iWlV/13MYe/0Sz3FtNz63KMPCUnVcyajSbRLGWn
Efjcn6gRFkEg0ddn14GutDqWRlYLwA1S+ou4tM/lagmYd2flya2bHhIPzxpKDSuyxoe64BUjr4k4
4GXl+aPYRAysW4nG1279jCs6jein+Tdbi9YR93mdAUE4xIHAE9meA44VtRhxEWMkN61cNRd50npf
h/oeLH1FXg58QIIbIeW4codBs80iXA3ZXV7YgDzc2mquWfnDRRDAiVDoWpvTtbu7bYJ6Zx0/68lX
QhOBklPyjOd5Eg5FS8Us7bJrOHISiP9ruONeyvj0cATQeibEjlAzT+vTUDT2b3Vje1Z7SaQYZze9
qTfQbPJ9exHeNkOeJt6R8GAiOsRpjwhJ/Cb1cXUAiYNfUT/vP8dF+y86e01F5v4Hrux13fRlzjPg
nqrFCqcstQ3dIbU37bVFnT1RovGJKpi/EiO6rbZO3vIQ91QBnhsSm0+/USuggHRghmUO93kQ90cI
aGHmUtTt7uuEQO4nVT0EN8jUPfhBzmRKOJZGk88lB6at1uGDdualdYJ3JIAf412m2c6wqfGwFSso
1m3Wly8gFQam94eezFP7FYvorh8s07lp0fNf/MOrizDuwZmct1O3dQPoAF0GKCM/7GLmeNVdTwb7
uPFMK84MJOlqG7avUwWKv8KPOA/xGb9O4B7WSTh1HX8Am4GraWG1+ZPY0pYW7sUh2jGOG71lU/xL
T+mS2mUVWveUoT5W/ts6eoEwXPgqPKQ1c1CSSYfJo1dw7WDp6Xz9WmySvNMTTCPbnJmXPRheXnex
b91oQIiqM/3aQr7gZtpRmodoV4H8tdq57n2gfTSWXWGelVP6vgy+7SIwPURotAgPCyQCeWKGGmFd
TwBN6BoeKMB7YPftO6Yqln2/pUIfmKXC59Kn8if1azk1o1/+N+kXcm+YHtcv6v3aPcB/jx9Grnzj
UruqDWPtGnhXedVjIu/ZxicGhV5XBYUpgIpcw69NqXhRN/gMat5nFyB9zEVK/LeOLH+eEAPy+aoH
qd44MxdOALRBt6XM0VX9pr64ULniPbf5iMcCywOxBpVBll6xoS+LK7PzPww/1U5onK7EE+ub6nuG
t8U3OLjBb7sf0miaW432B9YME5rgdYwMg8omsE5WXGAdiX/txam7klXRDY2Oryzs4nHUTRqdViCJ
/zREOKSFcdNU5olCWsOOIpbfX/M319ewFvPJcLoiGsiAu8xUOB6zMvgMSwZCBLqNh/eRBzSGldQ/
QCzYQyHytb7TzHFNtAFcoakCSPdCOzZvlYlTisTkZfT6G6kVqRMSMIKm4P1+Y9hmND0Vv3Yn+QSy
3g671C3zW0MGzCQahNBaFMkRuCu4AEXH25d1864MgaqpjrTJbYcWNoGTB6Myuos25yoYYWusSqP+
DREdAAg2xAp91rhruIdjjao5nfO5GrTYDDJTMILT1p1hL7TF8m720R7ZaWzXqrqi6Krqx6bniaRl
LjYozXtAz/ZD7nJuRMFvDBr9CkiI7ONTMbBnD9xNJd/jEFu8MXdPl3FTsvIB7bnMUrTxbXrHrl2h
MbJqWnyPJqd9GTnYuPtpNBwzdnhUkVubteUpqlvogek83nIuT1Iq5jMXCN06ScOeeEZcOtbqKfBq
EHox0wb+FlvtH6q8G48utpQ5IRCRYjJGPKT29EKGEXheMALGkDBJKyy21uUCfeO8wmueXaJGXmRa
JoXpY9FyZ1H7MJcJ36dxxHmMDQCsCe3JLwRdKbWjSrVvAM6bGjAfyRDUY/9a32MV6Mh8kevkNC/c
ChkFn14vwUcBhVbXZKdHpSJVhFw65JUux6E9wmdmwZNXx5DmXAom93BQXnEZYRr7wQ2kPnN3ajRz
PzW/dS1vnx/4C/zUdhufiGfE/zsNDEbf7b4bwnPzZyj9zF6WdvGqdXgYbN0fXocCLE5bJBv6gtRV
AcSBhSSZO9Egl0/rn4oFkmvXP9kUU0yqfUJWo1I1YXmeVfKoa1q2GwApQ0vdSJUQUG8yf9gXnZMN
xsWltekh0qjn6YvoN76MUcBUeSrtj+ZEk52QrUjgZk4WyAvySZIGRa36a4blKfXwXEtc8ik17tSl
Gk1i1TXxJlaf6Asbpz3kUABI+lTXWmuPkm1yqIhU6xtGJpaNko296M6ijrxTY9XP1zHguWGUslRM
Mvm8M5NiJtNpT2abJ74ltoJLCNbgyx5UeE22uNfBqGhdKmLv39OJdsoKW9/1E8LAMW7FMAJuFyR0
9bd/sUBtg2wc575+6+XwLi/V31QWReTXBM0AJk6UrpljMkZNxbMWc+ibUhX6EmUsKh+NhlVlXubl
FsDeYR8z367uMetWpIK3/Oa+C51jEsKikJqLKjwz9sdz95u1gH/+ZVM8hauNWkHWS3ASOOgyrz46
Fa0XFpsrkyZLgQjitSePWuvLdjj9gteZlR/QeRrRbswY/DAUB3UQoUylbFz7S9TxrS14fkc8LLbJ
EEAbfSzUPPt7xBi5PAhYyu3Evj4RKJQad3YdLOxSRym9Gk9OFSo2jnI79H5sx8MhvM0UEZFNXoZK
AFcKmWkl8gGtwOTxnErmEkx/EUHxa2yey8sew2GWZ1+v9pJ6rmxkxsWc0nsa8VNFd3Vibftl5gc4
QX15aJU842nQmEVeA8D/9d9uR8Pj5JFGseVTIQcbCTIZP8ulyISjXw4GrcxGvGus9jshFC0qlNxd
ai3m8xh0OjcGLERgEGPLodiAyDPJLitVjUyIyP97J5VtTjsFuKc0cp3R1NzxZvssr3IPtw+BYdP7
vbc2Gu2aZjwBpJAKVaN66dMW8ES6CLil7b3K2i0tM63uhn3l4nDSkZ9UMEqHNOcE1OEE70WkAM0i
qnn8V5SqmciivMziFVRNJMlCjeoKpAHve0ogmUd7a/fMI6kbqNgxFl3cYV6/e59a+1VttFs/SV+E
rZPumm1uxxWj63UcjST6w9/PLET4cfPZvx4FJGlGFMGhwXz9lrLh5mMxHSKoTTAVQ6wV9Gdrt7AP
vHAE31ZyHKGpt8QsQKrk9jJlExqPPYqOw0BAaEwY305vYzSLlGnBIv+1ehciRVoGwYlZrZt++PrX
7NoiQy/wamPU4u9e4Z+/AJp2x/dXzsv32DCfjFlPwrU6WyaK6Q270hd7m3e9Epb5beuK7Rprs7Vm
euCqtarL+yziDR9cKDwDvO8fZp9IVTLJ8dH1ivYthWPJCTGKpguCB9574bLPRt6TuF7OwZpFXvDv
dN8CO+iRBkfuYo6un0xzHALylbIWnpxQ/g3d4wH4s4QOPvkSDfncdqwCooTQhRw5TXukM91I32hw
NS8hfR+Wpv1I0eh1y9GvloXlkVxwZuqxkqb3AtOlIN9noVHn7Tz2TNzavmcgPfEZ3ahWCjcNix1k
ZWOfuZhvZyQoqRZ3tS2XfQYLMBDraJBriLT/gMCm7GUz1vbWzFyL/x11i4HFHWXpimFelpnKwewe
BlTyM3PxvMg8fvIOOKyVmejJXg4wjGAhlvH8q+b9NcLslbYxK6P17OLlrLvpLaPoWY9HEyvBGKp8
efKcui/MWn+J71djySeOvki7ooM3T0NLBgH8dB9xc+fBE/cY99p6Se7ku2wikeEgk/ZnaWVDFvSz
zzdJjcGXxqq4B1XCQZ4/crjUY9D0M2D5iow7bZJ8RlXMoO9olLwhxxlt5woUjm4UJf8kMNoQZl+H
gn78fzKCtZNgM6GKOdQKYCOu2AZWGq/50sJ2C3OY9BVJrudH63rJs3iA3ulHBTyj6NxsHLmZPsUJ
/QXmXdWxc0XGdF/L3EIRFyCTDcHY31+0SRPI+CpE255zLf62SsjQ/mXWo1RC6nX+VJIanUJAYpWW
tliogP6f1X86rhCcXcmnAwtTZHmOHiUZjCJPuhl2AXnytPbdDbdQBvNVfR6eexvca6jnJtehtfuh
Y1Rf3PqL5EEQkIzKlWummCHuF3XF5nFvnNC8CfUDVCFV9atWqyftrLSHPZWd5EJZKlM5z0lGP26e
xtNPgLFSCN5adC4A1lIkvms8Ql1z4DFBg+ursQD0L4FwyTZDDvTorgNynOGXudzZxv2cdwTS0+sR
7KsArhMZvFXP+jrEDZ7NS4qeCgsn1i70e9Fz36ZOZrsAytxM3/qgpBrU50AEqJzjM1JhKwHYfYGC
U77sbuCJZ6HXYA1JUrKqPbztoMsWeIFTqaSwZKBkr26PiRJN/8+jp7GVTn8ULxBN7nzD3DoHkrMp
949XAU3fv1yZRhzSK5Oad++MtKd1yUhgR7BKd35Ihb4I1Ud3gqOFtO/FRnfxnTPKQ3RiN4PrG5Db
Ie2W4jfWqWgzc6U63DAYbz5WhyQUcYyn4iRt/V1Ws4sDECKP02NPLcWXJQyJzSbt1oUyfV1e7c6K
NFyr/H3RQ7J3rv89mwGs4nvu3fxePzyz7cet5H6xNbjuuYiXvB0Q4TUDS8bfUK6/Egt8qhSDCDdK
jfFevs46IcHLWJ89aNT8ZaiBm3A2kHWqoOkNChlsKgi/u5dOQlJd7G9El/sFAA+pzKWhwDyFgbfk
Awcg89gHYjA3aGb9Qwe2kij8FClYKK/g5STjyJBj34AvZX0dC1W+FEH6Yx6GxzXkaPLJ5nQFK0pC
OitMpVSEu0+CiRp69hjcSR3WQjNO/kI1+ozg0KxEylSOgTdL3mlbDWWHSRELuEyBPxzRM3SxNUBd
I9auPc9gBpvTVg3GxVlxIPCZFqNp0fUixSo/NRFrbsrxhWB+2Xy1g5oMikN1kY06i0EjIEIJLzuE
PohOWVxB/X5zk08qfMAOGE/Vn+HLphJI5qRlmB+z+04YpSwfbXZxqX4Iu7wjgfqP1l9B2CLHa8c4
3iZnZiYjrlPvr4J+An5i4nhH/GG3lT27yrp7+0Ev0N1NeLAwxw+/Pk1u5kyP0fiUZXhgJPNUewuI
MUIoMBQuBMX3m19+Dy31oYtV1woLwAX9vxQRdkR8uDOuNZU39N4ij2/fRPUCm/zLCuqJf6Q3lv5H
zxuMCyhxYQyBZN+YhfBquWTR5zamZ7vHoI8pXOWmabCi1od1zw5NG9w+Eb0oaYRSYWp06nmEZCHK
+zJTJ/tkTg0zysj7BMYW57py124Q+lrw36flxHVzjxFOYyXfnYfi1pNPqlWucZVfEm4db3UlcUe8
5EO8a9uVgnfXS2aXcZZiK/6mpUYcnYi7w4Sd1q78dqctnc+IxKvtweluFmUjx0oDpogWA5svvMK1
90dZFU3wAc1Yivw23s6aSEgvC7TwiuwX7T1496nhpCqNmrbAfqerel9qNuGG/lFlPlebVQHqDiCM
6OuSoNcqfXwfs0n4AdpwUCULwlsBCLaCjffPV/AJTGh8rCIveIBXBZ/ktmDqMh4UiZICXKQovpgJ
KxInnSQJg8WrKnD9z48jTqb9rNCnM2Cxaky3HXFtoQynaXt7N+oxvvQIMqInM/OiNpQ0fwQjTPL6
ChjkddB4ouv2S3VCs9+R6wHP2daKica7DmmWCVMrdflQKzWrAFxZsHQmCKfh9s7otJTz8h8qhh4a
kDCn99b5tj8010DvPphDKa94AR/975Uhrl/dYEvHplaCsKqd+KpQ5k+UW7zCFOSdsH4nVzCSZ7yz
vp9WpgM+Zs/LI1NgTR7OTqj4s4ff3rCdgFi6B4G06aENhLe3O6ZZGOsHZMjpzGE7XGzerLLLAlFu
OJMrVG0EKaRwVYt1Dj3WTgAUoBktbPlxlf+Zt5MvTodTS/b4HxzycpxjI9ZAcuqC/XAKQm//Ju8g
U0TpznoMt8w7eZMEf/BwZ2Z5+FMe8eORJE5LlwjL4H9zUU7ydQDIF9DKdUm7XY8c7mntT6QjwDgP
I8rFBzsTzFfsuu7NAE4teQ71B/FpUZ2eEWUmE/Lm3wNVEltSA8inuxkjMSDongVrDch7kzgDRhbH
fnYA1LqRidnc+Vvcjo1sJWuG9+g2DDsrtVfLyLAct0XHU/BX33VuxN+iyunv8qS3yDZOSi7XZoTY
w9UJGWpgCM+OxSXXLg5fh9uiL9MJpmrjJZQ0bjcEf9JRwTd5BqE7YkDSbOrVG/etd1K+N9cgkmaI
B6sXm/zSj9xW8ZI67esQgw5HgpgDRMV7+BWGfyhaex5T+ZX9AN7DN4TQ+61jiojq1DmXPahGax5T
jFeC4JWxQQak24rXqLnWZMLXbx2UhTQG3vL031bJRAJIvZuKzTSgTmmKG0nm+8M2zbbFKXEo+SXm
Zmy2aX0GQx64JfpdwXrJ0FMbkgCZ/s9OO+qrqZUyu47/wJjWsu+49tjkbyO2YDFbirbVD7ylff1V
ZxNqbYIrsMbJJOTRpwIrRrpiKmeqLywLHKc0tT0SXPE55Ox/1vCGTotJ3TNi4F14D9WukGbp2OU2
efeNjUwBOdTDeWBD3GHJQlg//ZcH1Dd98E/IP5BXlaqAAmguzoHm9Loa8yI+hXjFF3/MJ0t14ODr
nItN+S+u7CULsUafiwE37OfjnitAAke3u+C9655O2Sv9Bola1+hskDE5PD99wrhCPjFGKoWmmupJ
TmXORaCAB5EWtW8djLGOHCy2K1JovJOrS5DUb24H3z7FP1yzQiWJmFzWqJluoXttW628Q9x4CdTt
KXJe3Ab1q+b3V0rVFKCiTd+3+8L9RHAq0Ld19UjUHsty3ht7+Vg1EzDRwthJmmG6HwtJi2lY01Vc
HQoI0up7ZRVnduDZTIAsr7vxFfycxBPwSXWoKh34gjOnOLnQYA/YhyuqOnm74PyzvkYZ07ZqNsr4
RgfOM/QKbtkGUk+m0tAmNQa5/DXatVZpZYSr1eFwUe2xsbJSwX34EaukCT5Rz5h2s4yoE/NvLcaE
MOg3KQXQJEcipL6ozPp1sT2lnfE2Hyn72KfwBqkgo8deQTfGUsOArW17qGh17MbkHyM1VtbQ9K7y
S9b2ci+vA509avSb/7OKp1xgS5OlJGvg2tou1K5pse+NHUJQ+wPoVZQ1uAPnsbuL8h0tfwDaN+mJ
a1QmlcctkF0PJuGaOG8XH86a7p8KJTkBkGp8+5a5Sg5REYddc+eXyaDT3dt2agp8cNryD5Aa91K4
H3UUfETxHQoRgcJ1A4v8mqrf05EoORokPqxCotSyCOgnpE0DtvbARnOQzzRO+QQUA7VTfI5bXBzA
XANdog97AjqCAD3rSz4+Pm5D2qB2hvJHA+MyY65DbEx/D4VrSkYwhJTUHfOBFceZXIBiPInmbwDo
Xawq4FoLIqZrHDmEEWuJymCXu+Z2gXRj7GQPWP9+k5watuoh1QDlFXMn0eZqCEn08Tx9VpiRpsXM
CnGN9lppbuKS0LQ33p2UtQ4UglRBPZeVgkEXZ9GscHM61zth16GeU8Qg2+BHg43+Y/47ce82GYwL
NOfleQ05lnY5wFsnluvLnfOBZ0nLg6XKBoM5gKMzjtAFFAGt2vqhzjwYINAAbIGpSPCXOXhxxVts
eVM/qP/9FvBYMDohbpxnT1EvG5r0/oUxAh/7TfNjnw5frEbj2pZElblcP9oS71IZLj5Jeq4dyLtr
TLPYzoIKSGnIL9MKtoLhD1wacRrtidNAMi3zCH8pLAGcHNUHdXrFsbsxCDINNQ61XVDK1SHEYtSU
SWvaVFRe2gVZSCePt0z4nHBE179W6/uyI/gub5s/5jv3PG1aWk51dEaW5bMyRjlAxP7QBpscKgDO
69pDnoRA/LDmpAtewvM63aSFaXtK8nQL7XbnPs3SvDkaluBGr4VGZ64ePe1Emf15RP3StDgJ+5pA
5TTv3wjQCmvI25aL+AgelHGmsosclyBoi6F/hR+8TPZdEy1sq9c7zaJGsDe1lP1s8nLx2+fwh2yn
GV8bOjdGWPzP5c2BvRbky6muFqZ+XsyflLKUjGBqbrnNrs+8IXtkR4EzKQPDpxLswiO7GxMUZqLT
r/WrCnB5lm2tvbvaRH5vFhrwebIqkHV3JqIiKMrnlMwDY4gZbc/YAATEXaerTneuOC+zE1dJLCnv
8pg31/Yyj6It/OxXGHYgGU48K+641cIO+O37/N+d7rKAMQ4StJ60lxjm7vde7y5G72tsfdEhZP4x
SIYUhnmYPRMJIY7/DFAhjUQ3NNMZsZbB/nxRi0hI+HfH472HKiwUACzb3F0kG8iIxjWiYC3/Mqve
vpt2Xn4C5H3RpkzeDfdEqQbomOtYanLuu9nR/YazQkMZCVwWlKXr838HxntSw/9HcEC4L6DqVJIB
+11HChhx/IMM7KDk+vZIYpEpPAYxPSP1TpnQ8sCzcZk4s48s4TQvDlPb0+l1hHc/Akw5k4b0Xzd7
ox0O4GsKttOMwf+UtW3AyOpgc/cdyuei8fwjMQWLQ6kKXPcapZnYYsNmUekPhE+CXmZagm3OYaTW
vHaxsFlB6pny/JTyuNlB8tWPrjhHSHv7SWh0AnTpMDy9xWj3TSbgT6jFBz2tnXu8iV3AlradCgLu
hkZI2j+4zwTF/iKsv6ByPYxNiK1e9Uw+9J2q9Ggj+neBPcJ9L5olZA9eEjOlVyUKPLDWmhZT/RP+
X6AQkabcT93PJpVkDKoDIN4v8ERXxiH63W9jAHN01Ua0yqNruQ2vNQiHKo/kK/OjQ/S9R9A9Jjd/
9tZGjYPewER+QhiwlaGxgUZTbViXpQadW3eMtokD0p0GZ0hFXUygc4DxygBZJdINfKs9xkzYmcOE
1cl7Ytc/D9x+uRCwQiu81GAOHk0F0aJKfhTnPCyq3lH/k+UGJZCH+228JVOICXK05UmjCcvmRiXZ
kBB6EsttKgx2ZFMUk7SUp6KEFunX3/EPbFB+SrIOmQv6bTWgFceRlS7IbAy4TlOF3//EdJzratzE
K2XDSZtfQjpn6GfVUWnO8xv0gYvWcDp3BdejAOwDE8sCzXC1mjmSrGLXx2iZygI8LQqTBj9v6mI7
A11m+SeQDkYbGjkixiTjftoZJz48Ay2m6z9FY0mH4AzEOIAPLyd9XDxo+opqOdFXb9vkTIGxKzj5
U4fdP4OmnXp/N2lULuzOVWvalGAqR1DHlsOFXT7wG2rn3nSYM50FDKGoY6mKX7nB5z1sBtJYUQQ6
HRvsc6axSsuIh/df1cWXKIircLP4YPCqB8p8+RIIO7M886fqbzQNRlmVkmFhH/76v+9/WUEFMpxa
jt5+F3ax/uMsLfKUitt9gWozRiVfK+nMiLFeKORS7MXcDfAmPEem/j6h/yQpBHm9K4UC+iPw7r5n
bkpETGmN2l2Nv/+nIVOLRedOUlvFcG45PLQcFVWKJpTEfxkdns7qw6pO9Zu39Y1kHOcjPc4PKW2Q
eV0D8eg5lZRvxoURWXH5R74MBq+ACzwvjOggGLlL50z082jC4h1hXKyvSC3LqqSF2oAsnX7C0Aq3
qMoiz/G+dtng5p2ZruOhRIMGmkUd4aQOwK5wi4PJF9Up5cRIVF9co5gzScCwkNcer0FDHrlxw2FZ
6gdmg07VjBSzGB8y+Nywiy034Z4PIdCYcy4BKYXrZJnR1exg+79qtIvuaLS8NX6mn0d2RmvUQYNs
hMB2Xem9dcd8qtAs0Mpa+rd1jXaz58z/FKArJ8sYJUQL21V0J/8ftRvcGhUc8mtyKyT9VBZucTmj
+qgkZx7b8oBiMI5ALfgJ/y/DnGI3NQLsTbBGfrs615JVzvQYtTDZPU/seE13NGe5Xk71PxQUzmdb
6KZ44oU5djjObbs/RZ9pkCfJZtbx1oEoByUhLAwIUo8OPWDmvb1L3cAGxYrO0RPb4TnSZK/G742M
bxzig3Z7lNCcHoOIVT/yhRZoo/tC9Fw5uxDGUBcNYHeJumIlH475+/5gmNs6mcRbGLG4fQcZ1Irn
M2Mm2CoNQHup5AzT8ox9EiHAOT8WCJ5E7Dv77KaJPfgaZ21gkREyzyqLz15fxzFBAoZ8hEihDXJm
t+HhN9SBciyP9yw4rmKkrMD98WUZEnvgQanjpqSWvrRgGNPUQEampBhHZinarZ6UZo9m3qNNR/jv
6Z9GVU02BpujlGEMxpqC3hcFvm7D58KIZ87WY0Fj72iLk+3vRSGuLZMx05CqjxlxDs3xdrLsq2yB
8jUNbpacXwHFryd4pEDLugWcxHvlGkLq18QXB/PrEpkEasGfIChDCstx8VUGLAwKdGOlQFMb6bBD
iF9aklHJvkI2bBp1RnvZW4XwNFJBc4QxDO2/iMFR7KOn5cA+3fcKigZjZkVpInSLRk7jlUZLY9HW
QBj5F5t/OADCvZltXjpLEQ/l1+A3s2dPSvxvu5Kh19i/6YW5wh6UZnYGXWekSBlJJemXHIQP6u54
baFo9juKzXyAQ6hyqhqnOLfh35fNrWy6wtIK/NlECYNY9qObebzv1r+32izPm5dToOMQvFL8dOBh
dWbykO6w5YsEXWD7ClUcfy0GhcxycVb5vYyo9TJB/q/cO5Lui5ZTj7hmCawYvRUGIOqP7/exaMnX
SEGsWQfK/jajT0spG0RmrQSkcCoRf3olMd9ocskjIZ4OeTxcz6g4qL7Qg6otFovBtUBtGssDtYxR
L6o3zpxetYTyMr006SUGJqIYD7NzDSUOoLPRGya/YFeEnaTgocw2HfP8n02nwhmTcyiTmbOLTwli
ONCIVx1k0kbWi8CrxxqcHmFuVyAQlcHS21N641HhztmocZOqqmwFcVO0wdKTAoiRqiXxO/PtlCGa
OKbEoCJfPdz8jnl59FcOKTOQMEIkGICuC62Txui8RZ5aNjhodB5EADFnK8HUuUlsBXittgYmTeF0
/y643CkhNysGkJ14p4GThyl7Smxj5MKhxCw4KiX+8QG4JAV6TLFy4OTama4ojKsbHcC8hFQ7CiE1
tV0aMVDUNzRALdbJRb5b61lxGI7wObqD3lU9bWQofHNJIzaMTym3WjH+5eNqrQ3kF2QXTVhX4OYD
wxQw1h6CYgTz3FU2JpsjU+UH4Q0Hs9IbjmCqfbb92u3/YKYXIxVD/GdsVkZ8AUe5fG979jb8YDmu
ulLW0JZKnoCVpKpMI+bPubQ60ualgIbWG7JRMwiUDP+gh4YVkyWsd57YvEOQcMyWlEm6272q7K89
j3GRt5YsDHNK1hpK53c1uAezenbFuXwQpI9QIKa5sNHiNVNDHdFTBfwfsLwdvxNW3CH/rbGGM24r
1e+Co3IdL/xObCRaNEyjwgyXJpz4At1WHm7iDviT0L2YHN+l3mVCGAi4harkFYOzddmLYIjsTPLG
MYhWPuGziaiFGHC1UcTtJg/UPOuXgRQ0E80cVziWfcGEwkItg+7zt8TwQnozeeLglpPy/+H0MSqr
XUnwQS0u/hFmhKlwmxpMl5SeYhAIEYyEMqbxwnT/MHRkJOF1DjOUwazTcKXvSvlt9ysrUhLF/foL
TLHm0sD7OfZOyEu+wwhVwAgyxjYVjK8rZ594jY7sAc3Z7Tj+VRazyJTaJoFpAaOjBfbvV31bRbCY
s1Q4e728thiq2potTkuwoMB2etu35i8Fkc054/eskTnNJp+VStJ4vZSIYhluDuNH449AbM8+KS6o
IZl8nPZYPVC6wuKG7XWdgpNekbYAP7zoOvA8/+dARAdkSUwaobhU3p/fzIwlRqysY857KD3TU8hW
hRKAgHq7cvSjA9JO5Kzs/PvjQaxpPUKjQCfxx8jVl6XbsIlRlnPpE+xRZiRscnoXxw+K4QKYGoWj
aOHnbYFapFq3QiMKKPlhMzyYFd0/yLvczKKPbm1doHqFg8BZI5pjXJCikIOEbq1vQR4x+gGC/iEy
0o0Mq3DKnwEtslAtwf6arkSftfiw8++jQ66QPIzArDZ9HsVzGPjMNn6rLnfZd0LHJIV050RfvXuL
TCXKWaTPvxTdpxZNP5noJh/o2GCVZpOJcJOeh49NBQv/VS7kaAyIZivf2uH/GuTpNjex3BejIJUP
zOUUR5ISeprLmmUC5rdkbnI4Og1oX46e7hCX4+RMcDBUDUkXa3jeQ93t9QeeIIfukBSfns2c5gVN
5Haakty0h0sNVTWtLsQx5lzkzONnkkiaiLYco2QOwteVyAEn0iKKLj3b7BQ+4zB/zHruArNAagzg
K1/37L8Lw4FurnMQ3yxiJqq8E70vg0rOsLwSlJtdmnzCSzGjaQRWd3Ke2mEBMQtkmK7hYGBJMglA
SufhJdxKQf+7CFCtdCv/QPTbgVBg96wEgFCcAgVQs9Ipe+l2RQM/ytOVTuVjliTQHpTkC614cB8w
FTvjMF0yyQJ2+CmRsysscVOfSafq1nH1M5XQV8ERbB7Jkvt/90vs68gR1hvhy66bTAM0gtTv7w/2
kF8HNKwwXQx8WV+MxDHq2fAe/fYXzYFvsj6xl5tXsUi7IW/ceQBZYRN9eQNW6SwVLzK74js2tG1S
DZ5rgrPXnIfex+ihAyFPmLnYpkQFJNVinAT2d2NZP9W7OkXBJBTnCdNK+LTLL4fK/MlDzWX5GlHm
PaSEgANpO8J3spklOuV9FSUuWVOsSEGai7FfJGhBxjWssglHOwWf9DJavXz9K+1HA2ik/i0POObz
hku/xQcSmRhRQzDluhMn+SmIvydAWRqjKEqsHYVg+MQ6/U5W684Gp2Qq8AJg6v260M5l5OEhHjcB
FmWrOocgwMLh2j4SsDfI3lragoK06kVGkeyRBiwsl2631bg0mBfeD8cBM0evjdPYyZ+DNQkd3nYw
HUjUzZ/W7fH5aSArC+4VOdOZXAjbd78cAog6+R/LAMTWg/JUjpQshUxDJK1BGfYltxvct4fMW10v
vEBeE/r5aSX8+O7iCyPaPd1yp8tieo7HzcA+N0QHrGi1urYkKje9Lfn8HN3n9AA65JgcCf8vnSu+
T/vrL2Crx2faD2Jjk3cqm37cJj74BME2/DhQfQKIqAdawYEZS0sbbmEUym0u5ZGPsIwlxg18KiR0
OB3yNdUkN4SoFR79WviMAnm2YzMpaOtjIp2CxOqCk+61Z1IrSLc0fEzDsy6LFGauUKStdl2W059J
M6Eagu+zHRM2sNj1CRwpAWAnQWsLDXpF2T5yBRaKWevIhymJCZUiHECFkMoXjeLvP7fYEA8DHtcp
A/etRAdj60EuwjuwT2Vp9pmivnPB0b4kW/QX0m6RV2OFbJOufrZg/yLqIaq1wog2avPJwBoe4UtU
pDOEQuxtdvzdX+t6giby4GZe162gCJigcmZ1QIfgZSncQyox5jacmkAWuLuVD3cW4pdKM59n+nrh
/KOZwP+Kto1lqiSjbyuh7cCQHhXY0RDzroQy5WyIMsAvTxaihAVXXzk3K1kyCDINgEPb8SRr16Jv
/n1qh5l/Jn3fc+DHlm9CR5sxmDImHSk1qluwy/QcyUKJ80yoS8zuChwvr+Lug+qpWKTUu92Kw3wr
3CvxJQd6rduQ7MnPXA2/VMy9e0bzZcDPhMP2tjVr0iFStcAqLAHY48hZqTOsn2QWj4m1NA9dcSh8
FYPBQz6mn9CQiZgsmAtvIPAU40F9SapPYhtFtn0ihPRBy4/wzwtfgNbf0ZxzbHEVCnX1pmaqacdN
YLtcXlnYab7/kse4xu9iZuLiN99zfHoNcKn3WithJ3NvNbv69anIDquPu0xLZHiM63ElrBYtc183
TYrnH90BQHm3vfQ5HMKI9tvZwmSyhA+iJxcRvVuqYnUNXYLNmZJUTy3w6NE9R1MxK13dhaEUs6mj
vewUb2nk8tAi+v8pMOXxnxbOtdAFqgU6or2myfKrytxwLtmOqa6UsELvAxFn8hsPJWSGRh0c1h/r
jcqcJtxG3sGaLSQtXv/WJoaE8yUaD45Jbhi/ZbopxyQgijcHV2pYoYHBRVntokqbi1WeK7j65zUR
Yfc7JuLp8lB9RFJeGTCMbWJJNYiQlv3jMh0wHFQckdTpL0QoX7+uJ//XKGQTZL0I+jIQAzXWjo/W
WkY5p4xqLz1wytqpbRt/t5YZFxezv5eKLhzqTMF08JpWvndWu4ZvVjc4GzUNxtmV7wd7P2vSXXhy
GaRgp5werHwawUDQbwoFitHMvzh/l9/Hyv7Zz/NhmlqqvV/4P6k8M9ch4Bq3TbdeGo5sho3yXTcq
3jVx6MjWrM7vkLmNHsYm+Lj46QpRvhaXkQsPXqfEnkY1qea+DaN5dhBrQ65c1V77YCbGWLsggZKl
tP2uCV+apL2kls4lURhBibRJFqsc7ui1EafidrMFVV2GZe1t00dNnVujG+X2xyvLkhuIWoVwaTM6
xHhjqYC5jJGh2xqSJybPri1hNhhnNIyDNvpzDout1AcnF0H0bBGvtrKQ+xB3Y40z9uowZwwhr/Qp
j+qleWe8MX6DUhpPkDh5O5gHl23kNWTA2gspEZ8GGK64eowaZFCntwumqXl3OsDA9Nxv87hN9bwi
i6VILC8zYa/Z3Vllp1F2L2vV1BBB3jbqhGEGviroCOfJYAn0xIQWgCeeV9oI8A6rG/l4WxLfxRIE
mi1f9r7bIuyrTPqb/hjl+RU3h/D1tLg9y2SFPGwwA+1qPaSOjohq6vfHKD7vBg998Yb1jJ1ivo3p
yRQksmynwGdM/ab+SCL4iPpJUuTEarFg7ty0MSW2GnLQ68m42rY7ZCnZ3BQi6vpnVHYsYqpF9/vD
MzaZxBhHZWQ7kwNuijnIE/4UH8GdSzh7GtKAXn2/qSjSygqEsdxfseidFuV14hn4r8OnMJWtlCd/
zvATaQBMSFrIEM7x3HGVdKrkUkJBOY12wv2fqu0XYrZxklJpF3CAS6X/jMpqDKa57bofCse6KbGj
2nq0ST4Jb1r7Xl3V5kNiKnSYDu/RVQ8YrpsGCH9k/5pwAKnrfyt+76JaEXVGsvOQP/QxyCeQthAH
N6bMuQcyu4JvJPkMUBnBrwTA8jdCg+TaBgHc11YEmUSc7mNsEbqVu0SsUyI0z5GJK43ZgCyuor9e
7QehdfyYLGctXcXkaoilMtSngZt1jcd8KG8H/Xww9Be7LTZp9QvT+bB+Slg3kfVo+V+Sn7DBRHUw
obQWX4su2S7yHNIEea+2scQYOumu7DeU1MuceXX4HNUbslCTEzElG4piTNJr24g4+SQDK/vmixuT
wtM5cewCt7MA3IKJ+ThweDZEKbYmgAOs7yTnfD+IdIYzF356ra6nuMUHQUcb0NNSPx/M9XcLR3Py
ctrNqshGAxllqwVbCQHF/d2mR4v4zFPOYTWNxMhtP0UNjsLEovxR+kK7iVbL5AjspMNFHpbHkC1O
nFS9hg5fK4FoZoiwra1vampkOXS94L1bqQI54xQA9CJRa+d0GmTvqDTwZCoQhJUBIQ/2LA6zJHY9
HpSzS1YPWHxRW4moIsZsrjLQNeoXadpfKYaynGhy4pucgPtb4zhf7YRNDqWh/2e+6Ee/1yomkeLN
IKvg+d/cN1lbpoBCYqjbJoRBbU4tLFKUAdUab20vVAcNbvRngLjz2mmUNgnVoiL6J0z88BVVYClz
ePcJ27YwaieEhp+MMxFNjO2/JJit60po4F6B0/IYB5u1vHKIy1OJZGI3YHa0CHKZpQP8iiSz98rk
8L658pgCtlmrXlkKufqyEG4MyIzr/XXSu2tYPacYFcb8WfgiYOQKLsqa8fMvR/gNnvHOvcNvHG/Z
2TGGsonqiIfCdZ2U9JIQqd+Qsh1Iyr6wkK+bbXtv2VgaGUk/x2brYHkX+cd0eFp9zkcGFUC6Tpb+
iEnuiM/rjU5UJOE5+X1hR20ucJIkWnxHB0K6VO2iOfyPQIGrHV17Xi+vhh9sIRcYyJ6tpXV7DEBZ
5iwtkugS+aqPF4pRV8POPs+g5x4Vmw6+lCw+V/omK8q9YhCbG+r/rPtPKlKiznNtGQtIydc3cfYf
YSu0vYYl0seUiJ8jMucVVTZK09/0Fgmc9xJWgkSm2lNlWJkdHgfH7srtKvqsGx4YBiojWLNxEp8F
D9blYh4M4AgalJyxpCA34EAPI0wquPJBaJyiXGUf0vIfsN1423wuqnof6bQ0nSVx2JqX9KG/qtuI
aRp2W4qH1C1o52zy8kLyJbETOqJoLtFU8XB7wnDWAJDffwYJh0yXn/HK+6JBoCHoDLNzT75MOMoD
r9eLOeFKxnEgO+hwlGSRlERUpPDTOyokbPfvfwxcQ7xpMqkhT97uzIu20Ps6Iih9vh5lcsPddpml
SfejF7KnUI2eWd0kMi7lN/j8mjU5kWwe/F4SEBGJlwJVmUQFXm8JCylue9j2n3hxC/1rJCaFZs/Q
UMMwDGK8r8wwq/bXdmdHFkw87k8bU9N/exl0Wzxyqr6sogK9jejFbarCbClFwet7kJaCnVz0/YMx
vGU12KW7B5x/o4eDbBCM1WefXX/7etv7TPGmtfY4d1c2Hiaz+v8wYd05xVaPuI11QzE7vbR0ljxy
rTkBk2OYl9CNYCOHGzjwMe5NJWvloiu1NfPyaRs5wusCPJ49CPmGFI4RQnxdX90D8eIyNpvGTQer
0bnM4tHLTWlf/X44E2wJMoMaYXi0cK97wX+/lIt5DafX8JloZS+KolgZPqIj6OxcoKXtTQ7zGxvs
NVxfcD/tDT802+jc7f0styp3Yh/H9sL5ofV1842N6vEmCUC0reARKH061IitG8NigF+OgAXAuFo0
NTHSv/UHdUxf9Z33Ur3jBVXuv/tUMcD2MhgA07t/TeVgWxq4u0/wToR19Z8vrwvI/fcAGOqnusD1
ujrV+jma1JRwwNmKkdrcMjEcbdWt9VEKhdD+IJNn7J11IOUPNleDAYxXkaN+YwSJDN3kfO+Kxgqy
5gYokv5awiTr4TR/8Y4/9zhy7Y40Cr2SJ8pXyw8tw6IzVRK84CEo/gRWxKHyZYRPRVT/tFbj3OlW
LqmWuICQ7g3oEBfXaBDIoowy6HqVuyeTIRit5jPjHJnRywTqrrstCrHwTT6lrhCD6WnoEiGo872X
++2Bbd7jO2HtacBBOTkpLYmaCg6IihHXLyFyBVsmLZP8tuubfDDbSohMMruDfkhuCunliJOl1kjn
Yt4ccSRYwmDste5fCZyOq58daQy106ODggNxg5pojZZbqEdbllKda7pGkkw8wk6fFq6JPOZ0NfyX
Dqt2oS1as0IpJ7WmQeb6qztKkZMtS0pzdj/SMddyU3FO44Dq0lW89g/aUF6hS1Y9X9+AP/S8fkOv
tdjxoS8DgOLtDIcfEeQ1CfVCnw/SFVBGrMTRrppLHjtxDiY4G8aaESx9LuqSquq2KnFiMaAbxK9A
XMOXuOQ8K8DEmhl/r33SyhXnDZ9fwp/1ugNDOOb+uVHze1jVR+BuLK4/8WAXQQxLsxF1nY2ZJW2O
e+h4srcUG5QFQUziaVBaUXsKHVgB4WEm/idJtUroCCUAeBWr998dsBHw7GJ0j4qdr/K6vpPMC0U4
LjE125jCZT+7f8+HzOE9Cnb1Y3IB1TVFUelLlh+V7vn70BxdLgIZguLXEdUd1VBSp9/tjr14IU23
ZGedQa1DVCeUl6N23xORaOwlS/+KMeeP1ETd24JxFSREsrR15cJVe8U3I0JlhA/7R0lbPxYXvdNE
We9VvL8SOxuFOEZBBi6hWC0v42rp0HUsYvf9BtoX2watkSWa+wg6CyS2VCjnGXuF7owGyxKy5UTd
1ZG0v1xvBMxu3PPYZD/yjk882YAST+ZnO8N7oSRHJ+FrlsWgmFpS4bx7ETuUWqsjJPkM1CKfKe6u
nO5cU7HIaxX/PCUU+V/L3EM8GqMN5yVKqibo5KBBUZxohfgddhC9vDWLum8icueBwuiSfKIl9peg
kYE42XH66yn1WuJm73BH3cAZ2TxOMtXmmqGO8OkezyVkkyWuOlz9kkUxTkVHXGbE4K6whcT4FUZB
s8Bkd0UxHeG76pvb+4frpnfdE590KC+Y0AAeer/5w/bS77Vgva/qKqGXua/bI2PnYLonNun09frL
ltaoryOQ8lWWrW8Bv5+Gbdz9q/urHHO3tj45Hi+7IL4STTonqj4rRWIUlw25j3ApKZOtP1Gd8zUj
B+neNWtnIxJm/0jWJgugmNRQ8uSRXW/kj/qaPLXcpoHD8eOwXSgYsJE+4hj7bCVi4i9gde25JQPF
T9oG/ptAP0l6nuZQZfPVW19dhUFm1SIGXH8GLUNLWxkhgSd9NOFmcB3QjJx65tF43ylg5wkKTfAb
z8uvd/XHoCe9ZnxHVUNbtIJr3GXuPOjeJ4Gn6jeiyEZTHgyHEeKXslNO12bCveZp1QCugYcsH0OZ
rKYmrVVvzD75GJYbTd9djvakcYi34ca4x9V2lc+p/X1TiJS84T1uLKsYDGvg3bShBLrnujgQOpHE
iw+HN+s1uuZ0fY3CihhTKW8piiK526jalS4syP3qLVK3OIu5Hl4lCNjtz/m7jseZW3T4vXEOk/Ev
1T/E4saTBj/CZyLeCj34L0GqtnU1R2SH0tcvWhBwReXF5u+ZSvM+UOn01dmtDELn5jg7DhmN/+8a
/1hNuJJ0j67rpspTBYUFa9UOav9f5fwBV2dKgdJgXJyCe831d3ql5x0TCToYhOUDHXAxmoU/8FWj
ZvRb5NGYRKCYi4BBeCt03PJcbnsY341ayn3kb7nEfC/KEGOucB+Hnbn3H+WeXHKh+npVapQYkMgN
+gOP2zamEKaAOq0/ieUy79/WqNwTUaJUd6f7/GpZCV7KUDu0kEA9R0CU4JszhwX24aMMu6BHr0lk
iL7J0NuwBzfvL1i7HMKBQ/93pvc/0+PgbkcO6n9jHBtJTmRE1OsbFQzBLP3W74WweOhCU1VbF/fm
1GH7Hgkia7B1wl0SAOYAXmX0TSU6IQrqmSG0KvN0REIYD4sSgcG6hARGBCwRP6d3BL7kGQGpX1dg
nTih/6ZXMXRQpmtDVev+xQjS5HWEXOqO4Wug0GniU6de5MjCWwLX5uaY5pXzn+NN04MiStc1zQxt
+7kucxFRoo23yXVQLE9NF/Rg/cOvrnG6/MPNxG1oMNgwQqvmvBc7bq9xhskeN9NCFudxc3H/LSke
zC1JKonxJNlyP4aHUWo+Rh/Bo4qglJ28fmiTkeEHkbJF5+QwssJKC6C6UfP6vRHYWunF2HCkWLnR
H1A8gwLqBKAlAv79LRzQnWJO0ZsJ1DuE6tKkxmaxuMcpoJ9TrimBwHa4eLQpc4D5okA0cawHTG4+
DDzG3RubeW6mXlPUkYg5aMFJxq9gFzKzyaTOgI+gNutifD6XdXQcDs1wUkY0RFUYsIr6dHfDZl7x
Rqx2isp5t/tkvhve23Qi2xZgUWBG3LoDtRoERuw5VmRsupifkjbFCYr8oy9ecTg6Z2bawidV1oha
aC/yn6azZgcs3w8CeY4RJ+mHP0fgYvfkULJkva9XtS/Ygx+CZiop2AZiCNIxmkqJQiU4miQi4eD5
7IBnS9x1DwqYWWtR/lA7zqc9N4u63OU2ZIKCQJq9MGnJE7jrUErLwC/O6GX6PwtysI9n7+5vtYaO
HnRWwOCwB6RhoEBTG+/H2irD7KWRx3aiA3CH6cgxJWQtGpBkcgjUNTLwqDsxxSNgFLyzaRFrGGMc
2Hlt30A3aD4voTaycT7DpoRM/M89/t48wsj9gRdHN4SaUWIppIytYsqPF3xNCz2gctGuQlQeZwPf
eVJ4AoFLeZXDj+2EtFOCmKNPLvYLUQLSW/mz5DmOd6ljwZ0pLBOc0WzQoZzYmZltbObuuaXEju/v
04Az+frPXsZfkzVn8HJZUD9tFf1UGFB+vIUPc14C9dQIW04zvQXIkQM84RlTNVWTy3XAHVqKX47s
XM480uwHewe5LpxdO3hCfhfPcZTkLWPlgoQaBAXZVbZvgZQdcoHp1AP/fEwJbLR6j7uheNLmkLOa
lVimNi8dMaEGMiZK2GUBDjs6/RGuevBE9od6Tj6nNv+FuyYn+g2KGWx+UkP1AwrPnTNHHdKYvfkI
MyoDMmuTEh1A6MYvHwxgDDuT3yTTfVRX0eipMmL+EsxpwDjF0owshmbUce/s/ZXI6m2m/9hgLwQg
6nNmrKlXmL4AJtGp1eV4msBPlLxhDkRs8VkZP9yTlur05cVdyJI5keEdRHlbE6P3zZxe31e0FCIB
kLlAe9xynspO7I+65N3biGryV/fxGXgF6AKmIzOQJLShhSmdblyrMUGvvnxQ9CeHgZ7LjvugWPkm
/S3/zoGDZIA0oieLygAHoqPSGP/jenVFcwj6tnmyRkWDLqqD9pjAdI9Aq8CgbVips0tQxLc533fc
K+wAb795rCUfwT/24GDWx1pbFUjjlg6TSM7qXzw+b/QaN/zVL5+afiE/Xh/CFNUfk3As4OQt7LsC
AxVH9HVKehc8TCmqMQUoVtlogIIragX4Mibpk+XbaSxMT732LZcmEys7WqU7gvdLQd1cSdEEzVXG
JUvYhQtze6PWCC6p1ZsmZaF/0lKHt2gze0Hchm9SqQ4v34bDqyUbjNdwXWNiVz4oh9iz5NG/2YM7
+GBG10DRLYPsUEw/umj4qZm2X7qhyEjm3LZbKqd0fQyv31wafTcFxCyWyW+iYR5KvsM91r3ZtEn+
xe6f/jYZNV2hBfK4hXdp4lKMq5PFNWFmYAOUZnTZb63ILvTZGJq5zRo5KbNAjrQ1VBl17ooyHZWn
0Uj9R4yJn/VU9r3aSK0UzPUhgPU7KOz/pU56Mz1JpcRATqi01sZyB0SwnFmDVjH8jVOd1khe50cs
j9QoPsKFTzxrm77kazndXlc2NHFmOo0Ru9blwawSHCOk0sa4vxyTeuWkO23JwlbnEEHn9AGpzOyb
pxle37B6P4sG6V5ySjxtK3okh2R0a57y0LFjVh9s+xBZ7v4HC8e9DDHBbbZrla4s5HmnjdODWSwM
mVrag2WuFJWs4gM1wfWCD9bUdEJQa0B9+lJhQmravv2Nc3MkLiQo0KFTcU2eG0oy7SKOWf4Hh6M4
qMFa0vIU3rrZQW3+DDVkSU63yH7fpPaXnXx9P5Ud6CICb+cBPwzsm7wcpVPLVRqvg/adig2dBKxi
ecAaYkKdJXj7yLWqZ+T4svmjEcs+9VqMH+9T8B7QWXXS9UqA3tHwsRL0lqv7dNYOpvOtJeVyyQEK
UUkDpitb9fZjJbRjUqwhF1F4U23bp3c8BeXmxridd8EHOsQockDVar80Zygq0pn1tAJQM+Vi4YD/
fkLNg+2mn6eXcEv34ofmuVYhmU6v1ol2bgB45iBIJWTfcA2IUUBjAI+8S/8uyBkPGrluEzTlwzlk
voKie5+iHkuF5/whZzXKjhmwF2PahoB2LyAdNDfUdeoTDxa+z/QXVZAc2Jw6iNB1ol4TNRZXbBu2
2gXOSv/LmAC/xe8I3UquT5anv34KFVqYKzyA+KmkPW0vx6UaGj+6It0lLYyZJSK4AJpaP1FYQmJ2
Y7PUlZNjDTpVMtzxRq03XDNerlLjygnfued9QprM/PE5bBaE3iKgUdG3oS1tO7UjDM4pqs4K55P+
57g5lneyZnBTHj8FI11BQ/GwRIPTI02s158yXLEdARUE5gUyyv+E/bF7w+5LxZLZiLe3h2WkJ3K1
/Q4u2CbgzYQzMJYbPAKcfOJc6lqabtBKshHSvPTQubcM1PkFiTIC/MdM6C8YM/faE9W4a8DvnFpP
ZxNqgEcq48uqu7kqm9hz56ZOi7JLMi7OQqyFcMuNiYmD3uRFtI060Y5YLi6x2REJLsZZdHXUKT7O
XwFYFZ7itYYNvT1EDsStQZNJOhsbvas4GGegJ5XFmFgMHBpT4F7CUGGgk2WICEs85tpfRnN0OTgv
opG7dHU21CPWeP7I3qHBQxZYRVvm9taKO8gOyjYbZP0InIW0BNQncxoxKE7cmoXq2zhKptn0v92H
fjePy/JNnkb1QRU2K861eXdQrhr5Yx7ugpDFKcgztQVBHz8y6Fn2zvw5aBZcO3DjTySIJhjGOCrs
qriCd70YM+zvZKBXpCbgv6RpqI9O/nbbemxefuu70OLjXkPPoZjGsd+F/vpiZvfuuz735GdIuAb4
1iyx61QseDPywZe3cQ7ghTK60rHf46jSg9V7+Xrn9OqxJuuXlA7gL1IwEVijGb3jIj9nbtXAuUV7
VGaSVZW1xB/610aGqVIuSLRIqNcP+0UP+UZUGOIrCJarzdikXxIK4bxflNWL+F2G+/cjTERgxeSp
wel/zU1MF0oECnnhst7mzAirx+xCMCrM3CI+w9fUsX48aY37yxetV9Dt8dR8qYKR1JLK5HNVojg0
Dh/HaSL+YLtr04t0cFwPfhdcfWhEX9lk0VaRApo7q+pk2IiNMnmP1WMVUS6MVPrn3b7yVdNC9/G0
LVL4P+1dQCAONHqk4UUPArWK2+L2B48ctd82/pmey0+3gPCzQSb6MLcHWwfW+kz6tqAyyFmzauSl
jjnV0OdH0sqbS55f4K5no+aN9AHEfv+leSUi/J1WH0Ull4cQhymXoaZyGFzt/HhwNiTpo6HXKoH/
mR0FvFIjsUp/X52syx1n34PDqGue1UmS5OfANlBxoUBrpZUCjwFU5BliW+PZlXmWfJPIsmntaIbf
VH1/dFwo78+3HyCcfzTzHMpA3iFbEWWxDUryTr4+htpILZ7OLLAyG0FQ+Wqv5T6zOXON9AmBvcCh
+XlNQsrNtAkFmS3Td5m89qPOBqBaE0/30kc/OfA8cw37QTRj7G08i1GRIlRwPp3A4CvD3cnA6oYE
Ms0TXTWzH/Vzmpj5bMbHXqWo/K2FdMrHuKvsgM32J62SfyyNiwW9k8jGNdUHBnJ1O9DcR2vBUEHU
bUh3dp0b80KAA1UhbUgOoPqOdO+Ic1wYdPAv3TWBmH4o6ix3tBbTLm2wKR2hbdG4WadTwdeCSuVw
mWeIqSeKZWL3614zqMwu9DDgkX/9pnjzZwA7PF9fgoQjsokfPsAjByeXzu/3BnD1ZHoUXD77kNKm
l6+1F9UfFLR5R0dCnk6HXkBn8RWSLwrTU/RgBe+a1+XLTaDI/PnUN9gfs7McTnTqR9NjtytrDWpX
Bw3DsHVR5IOy0Fh5hs41HXEMmILyWenNQ+sWswbXEupz5tQsVs6oQkStCbkjUdXqdQitSTXPGtwY
LJ3AAF14gkF/FmBA//H91AIco2wgH/tnVYk6aCa7MQ5gQJSyZyry0j1lJAL7CgIIgsoaG9Ax5lnu
QFYG+7MxuWsl6PZsvupgNdOLVKy+BgE5JSLUl1Kp8V+IyJnkA9t9f23B9inExbPWUrQ0sAJTslNV
Z1TwY47Z5qu44Ssciqa5aJV75ikuJVpQc3qjDPXkfejAvcOWTajRJ/YuSGTwJOQqQlN4IvBab9rU
z3DG4n/OOC+va1njjY11BVcRZQ+Nfzeyi01FAkXMtx6eMl5R82Jnpu3KHbUAwaVES7EmiAOpK5fr
PM6nczUgVstfBa5K1Vh375ghZj2sstR05pATwvdQ+F42hJYMqhTvceqZKwBVyPzspF83mutexDIO
FnRXgjgBGsFWj5VsmQv6OUi4Rph29qxMoPvRlQ0x+Ww7GY9bDm9u4nhYrBR7jcEdv3OcmehQttkw
9uUeFg0LkXHqBx56FSM8aCEoIe5BhY5IUKjxLfXNSxEVR9nRKFWeeXgPcjHy2ligcra5sFThgJK2
V0QLfd3KCF9sZtHVKZD92VEToX+0DAs3akfKFYSfiSfKU459VHwgKQ00X/UM0RTx8nqsE621NeJq
irbS2wA39odqjvHxdOzeUaOjZZosfIOOyGA9KNeP8xm2cTROxHwXaRoZhAMd7zjALemcmfMvy3h+
uJkRg8O6vHusX8GHOFhBZnTJlCRL3NFYO75oQuccxIgBGwlQhtfr7mD3JQtp17unaZIpMJ3J1HwI
szere6Zc7pQe0j0RSKYo2It8bVFeEDSgJ2obNyLXliw5g40tbxCzNDekvV2e9/Fpdtb9z/5ozlYo
T2jdwZ0kGSfGDItBl6w0toI/BmgkAU39zEqWxm6NsK3BiX+MrftLcgh3BLWAAcZ9emqnQRuyvfGi
Txg1PRZ03QBncJQaQkYkg4BZMeQE4yrHFj4oU0aTRcb0zIxESxMJNTaJL5VYb7AWI3QE+FdF0MXM
nEwb14UJHd5A4UXxzq9ml9TR5R2NGBF6ZeJkzCg0xXayjHHQ0enOd+WAi4lgWB4J6kZxPaX7wQoR
dgqV6FMrKCGAqjqYETv+SXyDF8tNLOeDZcDh59u+LVWLRKnPdd7ns6jOwKESEGA9ZPn8GBVSL4hJ
X0GN9Yx+UPq/8G6vOEATLKEyEOtLwft9wkqYMUBlw6XRyijMd1bHCQu8KJgNVEX6peJkw4QCaeHM
YkH2SAjNM4sOEA3IL6OfBfZVSSPQgKOVz2YCESohdUSo7kxnzx5wcVHimk8KNRZKPctR9wMl5vCg
VhRNZHM9iMozdw8ZonhZopjIHifhNxp2UPh6GhA8ilmOT+RSHlp/XMttoqUaw7T+Sre2SXmavvuW
3VI+jygAJTdzeh0FYEpoO+xY28fuzoNZx0yTgiR7vgiXvIWVbPsvua0mPo7QgfLFILnPmIxvg+BL
9GDr3cbmkeXrVbU1iPWbHKMfdTrQ0Tjl2KQwwUni5JR10UDKxpXuTqF6MPlOO+A6cqTO3HTPNTUT
Zn0L3e0DOwgg+u87jor+y/xuIaYIbPZsGOIyrdbMhh6OCtU+R7l/93Ayp+ojMmd+awK50aBhedjc
DDDSl+5oFiLWbUepyimpfOQKN/TnFSsVd3m3ro7nu27w8yM9tROPjeX7MjYoqT435813s2j07YpA
Uq5xpYNIlwYHzKYFBDTwh9m6Ubq+BhPLBkIabKLvhciP4yPqsohmq/wvih9SO8U8XM6GAjkz8q5y
GSFLvQJK5+EwW26k3Z9a9hW5ZSy50oKwWzMVgPyfdU3BGxWzQbnUt9MHZVB84ZapaQ07K4kkWXCf
42GWi5AMuZKXQD4MNhmmSQrY5D0C2vb+x7hBGy8z/0hkkQ886wZsOprmAYofLmrZY7iFDIpUrNVQ
CCyzjAVW/jSnnnnW6QnNm0dBUSQeK9Hp/0bpqZuwhTpyinqCVa13E5vrdZSeS7grWyx7Y5+lwnup
o8O79LozKwkoGgLcC2XpfneFdQ/ZhcN6i/0u3O1Mzpv9brJYymGQZN2J676BZtJUtFvX3WDfjWwN
LZncwvwK7hZUULCIM1kf1abs07FWbFCbUqAB+abbBOyTWBNUTS1tNAieD/Vwrh/vVLJYcP2qQFBu
SxUhXF5rin1hLH6pUwtbTdFaW8IhSorrpMdTma8o0Jw8V7YcALmwWmVXxS2QTGkVsGL8nwOBAs1X
aF+aOQ94KlfmYavurnwf4S1R/61DELXwTTHsnIvfPZY3Sv1llDinZ2nwyX2Yz/MU1v8WdsHfgSv3
/NpbzQKlqbGindkJ0FbfafIFfje3Hbt8DuGncMqB2k8XjkuBNKQbDmZzcAw5Q6Qit6LudAC4Vrd6
GHLozhJu8dObI5foYpafkpvwuhqXHRU4tqCXEbU7YA702XthQSh72sK+5Z/7dophXSZmz0nHlCzo
maUz73c7GvjSPqRGaCqYRFNnM9I14N2aRie0UDCraUkrQB4iGyHoikJsGcIYq6jF+kO1toIRe2XM
pg9XEIu6hmUONTbYgJSnhsuL3RHXTkpcxbNSc0n3M2ANCnbs+Ttmzu+ztRbDuP13q0BBJX0Fvfm3
M4K1J1tlTxCjlew0oWtWx33iQuttONjPIf2fjlYgbma5+TCyNsitvExykoZoNvceUoBipIuBBW4/
ln2Hxfz5SQSWJ47aJryLCa398ua1mpOe78Q/vztwFJ5zDI6LWPiTcfKFKNZv2XWHCJj6sUHsvCwp
u11e6QCi34RELc/+RwJHQfqpsTp8aWW46TOuTLkVId1h+Gpn25n76UaOpszCniVlxgJuqg+9NU32
ixQeBGpZWarQ1hB9xWU6dVVmmCGuGRCw5IFmAZQQEm84psSirLZ56MUSrUZQgkIHpkPMR0e7LkLo
TMJuOrC9vBZDdVU1xqyWyDRH9vUG+YaLnVe6OZI/HS+ybj6cBSKkg29lPTS9KV6XQ4MYQ5aSBlsl
A0Vk75b5Cp5zAImPOnfCgZXsfJdznQzX1bg2ZQJmeCXwNDSiDOlQty354o7VBasolDTZk3g5OWpa
Q/2oZ60pqHkaVa4pNuMoQHyzs8N3DAyxuX+L+KZN8sdoq22YK8BjfUy5SxuFEIR98w8yP9m5r7ei
pJ0fFFGyBwmjN9urrjPxSwTtLM647QayMqI0IakSQ5PR+/Gt4InGK2CUEx5ucsXKWI46dTJsG1Hn
WC63dyQbo33XotEa1Dr1QKKK02r3YDks6BowBVy21OBtaBCoCGS4pzGpFzhtmSLtm4XjXzrsb5HD
KAbXUJd0jwuFJI9hZ0MDUcmXLBiysu53ixlqGzj8EJIK1pLjSObxwPUj92cAHer9nfNgk44d79iR
daVHCG8xw0d6PgTGTa8KSnbEedNZdg5LaW7iqD+ZAokZH59CnTt3QZF/P+WOau7lyh2GvY4XWwXI
/jfLrMx8CM8cEJm8bIvOzHfHAhCGoTdzAp58M4is22J+0woxj59hhmN0JmWfgW6UfGn8cHBdHm7R
c10e3TkVTzETTlyeYsR6trKyCReejsr66ghI2FwUunl0JSYg3uTMe0IsRsn1h2mYRyHB+HV6jzE5
tP/3bD9e8SNeNM+ZxYGI3BNi9O4B3MKl0c91hnyvzuqGZKVrjdFoBGHbD6wwoAlQV6FgJOl7aS7F
niNP291OLZD8KDmhzMTkxck0KdZAun6xzgLkwKSyipnALxnMv5qNi0aYI2PJr2hgpyxR32ED3g8D
kZClFONjK5o5v6yo/4X5LSyQEKii899LyIf1Gi7yrd+Yvk+z6bXkxS2MigWVySbPO0xicGvuJgzq
s5oQgizxLpL7if9iVRBnf4xVZ65zE40eO25lAxz1YxjpKbOIn0ObzlYg6a3s7RzYKw5Z8wJJS3U+
90iH+JYPg+WgO376R+vQ/GNJT5pvF/3DtZDNxWJt4NXeHyzn/DjngFubnJwUTJ5ax/MAbDMhm6TO
BSBzbk3iZf4XkvzxmgQDm50BchOb5IDfH+PaAS05W2MKHzhZG16TzpinxoYuq5RJKYjL/krHgGN1
VIPH1loL8q9doIGoRQToEOLjRNoOy0XF8HvpTCVbNl6e0BBfbvxkplKdZQIccm7Un2FHblKyY9RG
d2QsMMzwBwJnhtPRIFJeJGpvt7SqRbRtCo+B5vPW4LceS0k8NF1Ic4avECAS5ED0V5bsovPXfiCP
kf7j5pwl0BS71irvVGBspn3iGas34ne3gfa6X3p2TtnPlbfgh4LTvc+vMv/88tDtYE/IHNSmu23K
vmH1AGnYLpH+sjc8xSYYOdFQwSme2bHkzwN+vKHWaG8Q4PzYDdf8+uAHscW50s8i7DV/K43cqyfH
04fHSfSkaK5VXgVbgpZlR/sCU9kGP2DJjJRSy1Phl3IoiRd5rLyLVE8+rQ8OuVCkXhcTrqjTGBg7
Ku7UlY63Z+VDFlSfEJ86bg5jcQdA2TMIobE571wVBCjiBf6h8FWXndX7KDqyqTt3yAOsxu4gWdtF
Z39oUSU9qVEDnnDByE7nsBBwELK1myhY8SRZ2GQNl/75Ixv6ga2nC+gtEraVrXfNxyZpPbWbeRDa
6uxjXRt+/h/W5UW4TgkLRq4EemTd7xO66ujgtmdIzzU88xnfBRDM+ebdO/1xEbpHLOOMl9y8iCvW
/KFWwoiwOQ8rdzw7OTT/N7Cd+6ZF3Ka9Gb+ozRa4IPfodxpD+5bWG/fMVUF1rbffC6cM+UBhyHM4
1AwhzcdxL4CEx6OWJYi6PX3tqgA0eNWNZ6Ko2Y6HL9CNkWNbr1GG0Tf8arDtfvH9s9CcI9xYUcGD
nIWpStGnVPhg6YdlwLA5rB8SF1S5in+77cIjbakMPxZSchrmGQxJiVRRIUo1hv+Ff6XVHypnoNXR
Mbff5GZrbWN2CsG+rQuOt8yfVC98ta9p956Phg6Z2T9KrwdsIlSn8fO/nvXRDhDq1bpkQ1y9z05n
xLeaEMFxnZOZIctbm++HT4VSWI18yCjSYNxelP0L9+oDkVJiDDkDpYYKZ11Yf4RnGZM7uqexBhnC
lGkluehfQimXgOQbbENwrTyJEvusfpaAA0gR2fVlkNkNo4TFEzM8NdjCh041lBJXtEwaiADzO+It
qyLfC/IoQStB2KvMe+uC4gl9iX5OPpvH7pRs66I+aFiOduXbTKboX85R5W8udztpv6MmksDTc2kt
SctQjF0b+9v3d2PcYJbdVkhNeAPv8jxcRZhCIpe12wDjvNXqoSh5bULXwfsBgnuphZAi+vfjHgaW
TlbMqcluh/SY37+P824tq6XiJqgQG31lqjh7GHFHsuSwZ+BQRvz7Kc59YbWXgj9MqhmR0xMphJyq
uJV8RI1W7E7DAQsvdKnoDpDSd9J8PdWmzSysV7k20pKmjAQ1p+ahe7+8RsnxSPHfswGZ5+dve/0q
0pdjyX04nTJuFrBaAaZ3/9kyENGneKIp5eA3NpxHhsy516K0hfYpfPNFh0FbwtjXOFAHON7bdbtz
6lQAtxDnHecJFn846MZ4GGtaSILPiZ0zLL5DPIR500WzZ6ILvOygYxMsOdCGYcxkq1u27Cj/CWuG
PwAnIhPy/zyLrYmcRH/dCVlEw5B/AaITmSiwyWl+o2Ywt1wqkx/6/tA39eALmi9/bNBUp1gWTajN
p59RiqNDU93VeXnRBHTOdLTChFrPKt1ZanZvSw4ofR1lJkgMEyN1sAQl2Uha7JpFCEERkEgqJBuM
Bj5V/uajjQTsE/QoRZv2zBavZxVIbGi09I/lyJDs/fBjtby4l6s1HwcR2mJscjfAMVet5CG2NPQp
DOrNR+9Gf65KUuAq1bZsnkZoZGdFAxiHImPmsGxBC95h217/t9kMSBrkUcmjwpCAT2pcfIsB6kA0
4P+JpnAZ53/uwQbNyyX29JxmUn6EnGb07hIZ5uDeoACOtwMc8L1QbEOLvRkIpk+GQwvYgEiugJdH
z6Iawr5XtUY5x9hT9n/91sO8B7cMd0PwAFZEGc2DQRQMT6GTNryVufQ0ZgOAnxM0fF8qM6uxNSo0
twIEDiPKTueijR98zvxT5r3qqBdI++AXjBXpp+k2gMrH2IH5Or5TC2VzBZZUBh+bA7itOeQCRkjC
s685ycCdJFyxj24OXKXmcqBLck5fSBcbpBZTmi4J+yHe8CWqixhnpIY5GN0RZQ/yv6UNis3jNYtF
w3t7HbxfSAawmF3BIYzO43c4NThHGbmcZ2mm882BgABmf2+MkNovG8UZTUpgbVvs6mPPr2q5L9HI
pt+7UQvzZbTZVOgy+cXJQMrfFlkHtOeIj8HTAbPqC1kf+nV5SSORjr0UIbBD7t5eja+kFzYtXVdi
aN4+PXOrg2gcUzskZwbRjvlgbTAIeei+w5BsXC8y03bn6u6ihLJC1fFETZwBEKqHuy0nKShzyi4K
cWCnFcrQYUTLgHZFLy2gl5kcjpRYIF5PNYEFrEdTDI5m15Ka2/TFyqzakp96HW+Wy/wqXVtpWfGQ
h+iTeeN5NYe/hYZ9s4L952653om9hVhoU+ULtHFZ50SLnGGi3zYUu4GXpfx9oC2d4pbKcbzA8RP7
7zRVjDfPaTvjBNf3hJ6X1M8FzO+p8JJeogd7hXyfF9xkjlOFJjkTdbSqAZnVTmtrvPVLiv4GXNay
SRltqfHwGaDlpdcfOIR3wUewxI5bbvG7UE2ub0tJEI93IPkFWXh95+neOatDfCRN9s4E0iF8EQxi
uVbEuD6KRi2XB6M5sBi2ubxKYGzFKZ95SNyxwpRdNOXNrTwZnR5h0OmCriRBz73ZtqU5hjHzXgzJ
4TkMkF3Gox8p/Tvj5mO/9HfQYewodkY09296BA1Gc1aic4A4+SHB623+Xa15GeL78l7iGPrT9Yfa
qkpREyLhi3RUvHMX/nXH31ZveOlODS8J9gR0TK8BkqMpN+4n13vdJioSqchOjOel9Dy+wl4b//YN
O3bIkvcPVxsk8tbMLijNM3SQSgkGhmI+ciOFnsdqg9GdTNL/MqDbqZHdNhMlwMZDQmD+pXU36jEr
AT8J0tDlY8Ew3UaHusl31RhSj6F2PPWBy4GJEJaKEDrZMo+FLlhC3AyLtlwIvkCqcaZbmDrb8Y0x
BaB63/T/L4DrvQ0XUXZ4WE1Mjmf/+OYuQUaTZCrIfTJ/RI4cHfmjByhgi8shcj5O79RhV70DPTz/
KceGu70jSnK3zndJyg1rbqVFswsoEpIRW1q3X2IaAsxyR/09ghNh9q2WslAKHejW0anE44ybtAIg
0sU+FAes3yI7ml/oZagAEWI1R8hBSeuuTnaai+6vSxnlivQ65xROjkgXJhACaMs/ttJyeKO5YkMB
K/y9ZZoB0+52NSfRw/nFeT9zq6JWvHVOc7rGAju8AErOuwE2eUQOx7HOjVzkyLscafuvcrFCdeDH
bQn/JkQWWON8yPR2vB/KqiGYjUSFN8LH/+d/wH2OEsB1gASuI2KjJ8ac6zmfLXjjZooJzfXpg6pg
Yfduuq8Hz97aY+Res6LhCCV0brulAI+PD5cbR2or485jnsIo5UV+YD2iqqeFmGezCZ8YDUbXFuhO
hgrwPBoZB/TeGyBlxIoIDAa6D8A+ndBFKghJLu4fWOUqQRrXycU05uH6yBha7wvP9uyTw85s9AgX
uiaRznrGioo+bePUiQUIKqWH+crA+gBHhXsRr3YG1gh+J+LmxorGsH0zG6aJGpqa6KawFcRji5eg
oN64TNcHzQ+f87Q0BgzvizYgcAtkoabRtyCufabhc+IzD6WT5le8jJTa8RJbJGyD1es8z+N/lH2g
Oba220LoLC7Rjvp6JlnW1TKUXZJVpj72rO8C/U4aTS2Py6ouMKKE3XRzZttdMgWZ3OKxoc80Updi
kGAYjUBPIpjAndCS3J/VEyRUhKkCc2/vhw6ct68QI/6wXEdusWUbE7U4cMhF9cK8I20IwKBYSpLW
6oDg77UD+jajD6UegN7lwymvT0YO9hbaRn7l9NcyJdncUM+UH8NTHHEGEnNP0/DaeUiLbpiwqDli
lBq/LB/C3NWC6/LqpeUJiOw4lMRMUecWNkdwlkkte/9laxO3RSzuPgwdNqbH6Pc4DtFpZpESh8s1
Fs9KPdYQoWUNZeR3D8BqiN2e9MPDLoeqYXFfLAL8m4LhbkbaTeUF5p4LLikWmMTgtDI50sCTZQkQ
OwzVP0jCEo6iACB/YtCVzJo5x1FiaU6xOM+kJtugXvSy9k90lciNiDDLxydbwNhjviiD0ah0Gk1N
LzA8/zDSZzRxMZ4LX9/mOZpaFRkuxjHSAWjwv4OEAEo4cgLjvUx4TYkWNnEFUNKldHpxi5VLF8KY
r5S6+kuu4h3ucRDm3kHxZHR4O6AJrN++nx2nxfZeNxKEVCAdYJo1Ox75Q0+xE8sTqJ6xbzuhfsSr
8vMkZoPCcZcyL7EkxNz6+j0LHk87NWl5SjkWoZIdIcufJ1pOAKzMfk/kTUWFb0inosJsARjk7voE
fHk/4rZOVYjXl3RL7ls3W9c3Y5SjkgsASBGQn9rHwH1VsPL4LNNsLfT0/EO1h7u0VDLTy/JYtvZ5
hiWJyFRT71J2OEln1FK2u1w6KUbZs67DSI189FUPHg7sg9jKTKo6H+PomPCDfpgRQhd7nWiQSnjt
KLPMLsEeRDR5aFn/lknZfxcROxMGlDaFOCLx3BKq1UI6QdHSBInTfjHAvJMVogrsa7XL1uTkcVyW
35BWlVjOCRHo1vhH+IwWPTD+mo1KgOjDWqMG6/LY2gkQEyOOLdvVcAj4PNRTePlUYOZXvmeXE57K
QI5/m4+avBfN2zkmjp3iSsDv+hvoS+fQiy8pxUgksKx2My+i8BMRcbIHLPt6GAEvnuEJPXlCtJBo
1b+acBtaCAFQTtNTB8oSJk1NGFB0dbvczFj+84rjXbGxNpfaqPBk8CMWqkv/tY5DrFvDRwFAU1Wq
XkzBT1l6MdsLlUYd6uh4syR7Mgti5ejCPO1AnKRPHyxo4VuphcQ08/amgpr1QTrUkgykaXMeCKGD
51MLJC2ZC3E2zZhdHC5R/3Oovpgrj8Mapj0zUcYV9Fjh22NW1OGP97xdtKRMVsGca9AyiKkkG/PP
bkQdwQd8MHLywj/I9E+euaJPfsYLE6IF+rhCMqepkFeGXGm2n0BFRuTT5mXQNbxby9fyV0VId/N1
xg69j6UCkqXdtsDYgrHcWe1lF33j+TCfWmllvCm4IJd7BRHXIQHTgc7tC7tSX7uhTLF3qZMqDMf6
BhsI7UMV3pn77y2EKGtP39vRsINySnRZ22M+QCfaFnrhjvDKK4nNjtAU6jBhAkytKelOiDQ0Pq2b
XfQNYHKYvprqwZPOTJe529MeJdisRQijzR+P0ttJi911ElQIdpj3/PBnDpBASjvvyPYOnSB+/xDO
Ahf6GS0DimzeR0OaYH9GlqL3xReYhJdU2jQaqAfjxCnRogJTLya+uXZGYDeR8dL0ZOoOx9xEs1+s
nbxQSRf3F4j+yo8sx3Vi/I87coUuR/s8HJCLY2Z7yll3/RrjrJh/rtgkWmpWMZjYaQvsfFTs3pGs
NwHCKYZmHznra8SrFgaF++0UXrEsglw02XBKTnZSjkLrcHZXC5EyEOIsA8z+Sgf79Wo0uHNwfzmu
+obIbB8f4Z4tvaKwyO7y2iGZtkcSAMsCYZoWaK9X4ch6N7AlJdKuR9TVgWD188hrSlnftXN75SWj
N6SwfuuUOSk5oF2Y4385oBEFvdT5COkpEiUWKcjbWZNj4VWxs2GqXJjU+V0wEi6XeAwKmOTGUibQ
9oY9qewU8I9CjYXx602G4+5geVTg7noyH9DM5YKswtrehsd9dTySBn11wGgq3siuVddpB0dRNAg7
rZjriNwUF/g0TE63Xi1orwQtfaEKmiwYPvG4ri5XOUs6m6vJIi2I8u71kK/ACfHgH4y0JqZ5bHTf
ThtaWUysQHVAJblytMwetd4zh3OZiTV2A+vM4mp3fVr5DEeDmCMs1hWiRrl/DAethTmA8sOiIP1m
HFHI6Ea6sqs/D+gD0ApaPfDy8ipRJMO2JONjrYgZry47SLf4ILGuXre4fl22qdmJQzzWeEZvCmgl
z7aKlf90c1vYzlh2N/jVYMrd8LB5HI6Gha1khLzt3YTRtvGMh0ztS50i52OD0o/Vg6rrU1Lknk9s
9+8sI5C6nliEU/oWv1/VJYEdfcSIjz6kUkHlXPQJo1IdzkfuUcO/+iaVvHTEX7DWFUfMZMZ4iBvG
2ZDkcdy8XJNLXlmU8S0P6FvV74CzowFY39ln9VEMCIcj/m8E9WJg7sLiOuU4pbWwmdjXwgbqeu+M
c5jwbbjbJcBXNFOww4ZeppnHdFCg1g9rLp2ZcIeq4zK1hx8KJNZEiAJj1Y9oA+3G45Eut0yNd6nl
qh07LiomgNPpF5nvkhuo8JneSwHr/HEjq/JfTNNdvmAa0m0FVeUEYoU3XzfElPdeH4PfiKiTVOlc
M5wYp/CTitfw66Uaq7DxB22bUQer0YKs9WbC44JlfPPy1DC8h3DpA8sL8aO2CSTxbVWypkiuwbYM
7EKr/T+bBz9nSJ6JnBgWurd8PTlyb22XskSfXKgPLLdMm6aVeqo//zjdhtivDEqj3vk3rgXb/d8c
0MdVKflYZT2OAnfwO08KmL41nhXwlzY6DdZ4Xq2PdjUlUAsFjCAay4m26e+IwXcFAJC3Y2WSC0Ff
hc22pfNR66gne6CWdoIkzHLFC6FdBt/QR9ObhzlFAZAOboJwdavmXK3jha4cal6HA4p1OwKts2l+
gDdO9+IXHKprkUfSNF9eRxixmHcse7P4+8z59QY7iEpPXNJ+E4E3S6yI1MGqmLGilZxJL4qvzM7w
KfnXSP5nCf/jVJi3Wny0sn8eVayp1nsPXk/FP3sMdmNCkXde8NWNGaF/cdfiLZxfhK+bv2cDTPEe
5c3BBNGWghwsujyMYFKqIcMyVD32SlBOHO/SZR+wh47bYqCzbeCVtFIXRv2/+TjqZ8NhZhJxIw/0
GmtHXhzVz2WT4NVsdYqvC0EEZDJHm4vVsJyVUHhj1+2YtX3Y8Vlv17m3hjutg3d3iyRE4J4v6FnV
y0O7+gD44zXaDahb6uidq+XXcQm8UUz71zhNtCWRI7YgNCAckJ2NhEUmQjdR6S2WIaAZAimYudFI
6aaDtTqz4x6jMexQML0iwUuolUajmmqEKkv1Dpe2/5Z6KBrLv5rBTLS+qvHVP3cOk8EWE3RLkrFt
3K168rpkg8IMBLoxc5k/MvULS9BAp7/phuc3MbqdyHgrXHwKUSUY+phknFxktBkjrv/iyLKjp6lk
Nl9PxnRAfQApvZzYfvda5PPVU/dQOvMwrUW8HdciX9WlzT0nXrhTPW4ofP7gSqi/GAbkXwRjYBcd
sklr0B0dOLAYMd3qyMKYtRNZP3Q0cga95zHvbZrcSxnjDwsa8LmQBVtKCFhgILAXvq8j2BsoH3r0
CxOXvx6VR4E3JXZVr2SbOKRnDPiLCKDzR6oThAc+OSYmNyCJKPQ27gIOG5gG1+0FWw64ypxoiGMw
7o827tynL6oR7pVA97RvSXeVe/Qr2ucjN176Ukm30LjII8GNPu2wTP+yA72ojI9sSr94e6qGL2+G
VvSq5vPoXsWZ+aAHtV08z+dYXZBf+JUu0zYlsqNDsVJFhrncIotgMXf4tMYDX5gbj0DibdFJFFgV
JzAwxcUMzjoXdwUIx0ZUy4sTQTfQAvOaSCnALF6vOJrhavkDn9AGqJdAFiRlL2s3uugiyl8Kk7Vj
v+vvPaz3ZewTF8CK+ClVX25oH5qZfwXop9sOUeoaGqqsfaEs4+9YV3q51yrsTHtWbrAyXjg6UCOt
Tw4ldybhC4CA2LaHUsX9BmM5qISAlxtZtg2vxEh0jVVnzjHR//Nikvn35yVp6IY1+hdAKY9soCDd
39C8Gliy+FhgRA2UDQBJmwTDmIDMN2VssQIeBUYG3EVFgLpcbo2tWu1srOwS3OYj0AzXrWTqPWAX
OU7DbP50o9ONFhkieXZAjocac5KQPjXjquQbsqr1XYFI0C5qE48ibVv9gPexYLSgBhdB2HjCFRE3
1IiVSy06bbRtvvN1QRM5g14dd/t2O9bNxouWabcKv4Rn5EeZHV02+NWyMyXO2NjYUCPTeptymkwX
7KD5bHh9QIn0t9UgiuQFrTADN951yClVYJqk7xq8wi4DRJsGS9i5kt0D8gYFeWvkBJ29YdECDnG8
snhd7Ogv73+HfId3WSOrU965objRMAJHjFcWNBshIwCZJlEW7sK0UN4tt424f6JVWT/xBE0MRomc
mLOAs+WLA9oa3U8ZFc2UZZMVaIiD43+cKeELHRTWTv4d2vrKIARUoZivm95i5ylKn8Swb7hKnoJR
AWkTDSu2dNLBwCPCLDYCD3baLgej2YjAD6pCPSvI8LhkjPo4PkWUlVU42qNHzORkS2tJHFeF17YQ
YST+wRiV7KvFzcRgrw5W3aHZxWp7A6Eg/J1SQjyBCmMAMbotm2v5O+QA70s8rWq74nKK0Gc2ZFU3
qeQXZKNyTRcP03CT8r7uavhF+VA5oBTdc5loqSCiLltFzVzTScs/N/u9bikrwGe7g5UhWRofGJz3
HaMvhNf6UoaU6q4kIN0ehevhcyBdr+omUNz5h2Mu8uh1c4qA4+f7qJZ6QPuyyOpxOQgUeKAtaVdj
OWVR52HnDZmfKsFFhB8NFzGy2XJwJH+xYfRK1RRuqdIOwe8FwBui38zDCEcPUq3gPgXPOmijIcco
QqvO76GXgb0LU4QU/JJ16V6Efy+whJP2LyiMCijxYFlP7K5XVPhtIYJ72/xYkaYTe62cI/67O9YC
4/CE4aN4Qb4lYdakS+udeVYMIt2hVn2g0d99T9iGHFdeFoIkoYgmyJbw3hI+QgE3sEpCWJ63hJcI
7A/7AYs1O/wB1xM/BvWrWgSdplxdC/G2DF34dHJe+FbUSBGFRirnuHScXDX0bhL+okeK7hLqpkeV
i/c/UMcW/+HgClE5XZo2x9UiBh0TntdgHroH3dXetEjV4f7BncD0KU/afXk/DsmFn2DzWWDeRlqo
dDC/joImg0o80v3gFy55yloaE+7h0SXn78crY9hUggG/jOSOxIqNxC+/E2ldpSDjNjGQWlxn5eHw
oT9FwG5XmhwR4C6QzEFZZaxiztIwu01z6mve8g+yjdHkkojgUBgGJhOvMvMCwfsJqt3nnuhc/jLz
lFXXz57oK9OINPrB3dCj560K6DqqKSBtOjLz3akceVJqG84YCmX2RpqpKta1Ul6Cj3iICrwgQxF8
K5aIExSvMN2/VJNhf0ANEh3dZw79aayiaFTaJ7+FKtnzTClMQz74pOzCkjOEQIuE/tUhlM1Uw4Bv
OJy1TTWzduOLsRE3AZTU+a0y2+pbnJeqh7SJ1rApf5n6UVpywSWS+0n1AMosj4nrYAZE0gwEZHSF
PrSkaLIaHLe7UihP4BzNxzntMAsFJ+kVGGh6s1qb6e0LazG8wwu4rU1649SFoc0ezF9oenpFMF3G
TzNCrdyBj3B8yzM74cUNdrV7nwKBlcutDQt2InjOY27HuuIbZDUfhoku6gY3Ypm3djEzg0xJDUcM
pI2NMgwFqBTPTASvpIoEDURT+iQ10KiBR6BijPqhrya5FJ+zLcqeHwkCKQAoUigR/LHH8maNNFwM
zZ0k40o9XeyRCuFcCsBcLVbzWylOERtExijUfHDh++tBvJYALlUHJV56j3EDs1Lla5I5+hZjgyRl
IGFnm/6XP6+t0LBOCQQyyEFd/fRNM1aJg7JxU2lMCozKczifsZvCMpeBzXU2C8hjqGKbUT6ZKJdH
VG5ZyA+vDq63saVms/fRywng5dNNqTdt4pjutXhqszsWuV7tSkQblywn1Nt+YsAEjqFH/I3VtynP
0ZuWBEvW7bzH+rTkFVm4g4dIXQysOtsg1ibAKlg9EIdfkaAvKT5JBVEB7NXbTJHnTGE0ZzYBtyC/
oEhOs9luHd+64MAzhZR6jnGC88+ZfINir6068SS92w+I689EZRa/TQiBCn636jY9HwYX/CogUo3b
t8h2PSkhfJIPfKI8+cyH+E+EfXob8dPEEkea1eocL9JwJdG99UMMC2dt4PPS7qjrNuF5DMbc9FNl
OTGBpqtfy2pSYCTWNNxuKzqoGC+blTaw3W1i0BFxTDByevd97GZLNPFACxW8NWItTIzKnOIzaaJ0
BnniDQDpisHR34x3aKJYHZ9RLg/IsjoXQPyOtB9AERzqsfbtTb97sSpr8ARbhMFMI/4vtgX5QDLy
fTPs0clh3QzfxkOys0DOe6BAPoXm8/1Hh7Hp0sVvqn3bv98Kshr/Np8SBJXFULKhTh0JTIO0Ku+g
GRp/1uAa1d94EB33nPZ4qN+sdVvCWQf1mU/5IwzIdmp9pLDMsd81cs50ccLPanlGJNNeQF8PQx+W
13nJgiNQ6QrtBx+zf+jEQKtAhGbgQQLveQ6Qd58Ok4np9hr46XgMFuCFkMPnM92OFoiaFo1/cxac
8GUKZISuJvJA9GIX0NWBWekif2PRG8w8BfkUAneaNPSjzDDn3yGczyC7GV00FR2AjaVZuK4DcYx3
n49vFAZOqns4fVi7kuVLTFzvhKEnis8ge7uglJY7NU+ijxtETsz6qxW/2Xfh8uBVA5lXG2lAbXuR
358FIE7Yw0JdT221oSY8eR9LxN11e37EeiCxBVjB10Qk8WqM9gdz0N5TIIelAMByagbEt3COR6d1
hKBQ1cJwjesUbYnVz7iCCZuvd9Pdul/4SqghlQeXksZTm2YJ/fWao/sCyl55dI8qfC6/If3GWAr0
Tn9t0KHCPFx3uRv//FbxspZq/6Qq//a832FniRvCp3VCvPV05Oa946BfByxpXJqLUQ1RdK0eO011
ydjwQ1iAqSyLOSAnct5hEjeiJwO0rp3CJnVDhqb4HpK2wRIaUJmujSuw9Y4l1nDddAStOgcxjfEA
+dnr7lMzTiVbZVsqjhC0r55aVNnsuLw3oxHsV0jzyTL1YNfK7HwKo/DWdmTkt1GBqXJXAdnuHJrI
uY1UTBq3Hr3gvzVjCTMnO04AW6oz+3GX837TJM3cbF9mDJ0uwTHoj2rq622WyyMoe0AfNDw7XcEV
TtXwde081b/RXcz/EBVGA47z23etR0s2+ujfFctOVtnXl3sOHJS8kBWs9OOHi+2mAqdXIdnR21b2
Ewlt+jtA/p3xi1hE2GWuH0V3r4K7u+eJrM/D6Uql9EvqHA518/CwHYZEf+1+nxWXhuhQu0l8TSIf
Alf+f3XC0DSmJ4b7Hps0HWey365sSZNQzUPdAdETK8mHj6Z3j0wqeIFgBGLa+9xss600PjoisAjx
1HigH2jExWKjUrBDDWjyHT6OCQ8RzHTjPvnHadomG6p2eLWRLAJJ5GSAEd7FRDZmZZB8mosLTwO0
QzFxNC9DgdMGY5RDua6cj0wBtuuGU62udF8kn4lGTYqUcakvztVmN+kHe2Wsca9WKc01LrOwFZ6c
k871sVjARTdMqFBZHqTLUUIaM3UOAFx6SRGfxCPL9fxM3jOTq9lHs1B3uK4fcty67ERBNupi3BL2
YF1td3PiYbQyXT2mcckQBTpNXx2G6cyr2z85CHnIQ885Lts2bPQ8TluToErqhaY1v7jKF6vs3XkH
hp88haAqD0Ow6AJ0qtZ6F/15UAKlHcwa86od4a2xMHoNCRyOOWLNCH2IqvRncyAiZyin0iuINCWa
OwHiVmbzypkZgahJuaq0mjjBjDMOOqV/WjSsc3JoB1srWGGfkvq5S81TfLmYLTdxEDY5YQlg8z14
s2PSMnRT2zTHZ4Va+IqN80kBTYaa7QuYdlF0buAORxmxfPXAInTbfpXKHpZv+SQhdLKrDJp9ZkhY
JOlDqSnTE6F5Ih1YZagX9eJIi6WgzQi/5dQhmXPyILEesXy5QLUgSdWfpNs9He8FQ3tVRARxPTFN
+BvNbfBdlexX4o3yHr124xWDPjOsFo2xCygLhsWEYH9WERlz9nMm8om2ylGL2hOLI5N2OL3GBto4
Ze29rwfFNcSPtISu68CnJymFVGTF6oH2k9Id9AkMFBdRcjdEpOit3uIIKAWODJQFNHCdCVnFEzgx
4Le1mPGmmG8s+7Z0Zu/bXAIfJJp9EWyZtJBjT36LFByCha3/EVDthD0kBKFiNjA70XZSZUEbQAFT
mNjKfBC9UcSRBqLcvWAnfjzVcBkd51pzTyauvMRx2PZtXxQEmT5DzNs2nFkGq9a26aLuDrS2+eJA
EErsiowSmvHXp0zVemcMpwxFkf1wef5jhd7BZl1mvtZczLhdrCupXIXNTxjA2xXY59GbRcBZMwZJ
YQwXcSgRPuyTC3DOEQ9d0DM4/YyZmgZQSOGuQu4A9qn8yaCcTQaUcqFZBFPmzDzSwO6o3Bc6l5Z6
OoWj2hrub5iNGiP3Qvk+SeChLNoKAI4zjERg2AgHyI+5lW89/dMdmT3/3lfBl5USgBxJs4dJcekB
YqDmEFnZOqBrOmdxLjzQIhSGPFQ71dlYxrRS9Igb0smBWtPh/TbVoA2qeRy5+rbcT2ZyNVkNmyEG
oQUshTZCdoc51YK4cWUiPttaufXmqku4QWtA0Z0O5vYYV99kXioLwYBmZAJppUaZeZHphQMZfwrY
VviLV5/vGa/6ZwgtxMMLK85+Qc2JDs6AyAxln5/uB1JNK2tIWGAzRPcGI7o2jx5Hbirj+VOcJ+yH
dw6KRl22ZIZA4ympUzsR4eHm2dn9IadTcDK1M5pHtfXvpHNHLVBHhb+xQdCKFSWky1tIw1/fLEdd
BNZY4+i7UQnkEWbRbfjdDhX8prmy+hR+spIN+sFGQKzzKoB+w5zO3RMO6F8HqgnkrmRpciH+LM+t
2a+A+N1HojA8TKqn+RJT5kt2dzrBwSpGPI+y7bag/ZVbrYIDu7Snvg8s4L9t6F9OS8tA3v6+ZUjh
RPdItX2SGSeHimYV46QLSnt48yhZJQiDkXZKSE5JUqmtfGkHruzbIi8nk4vtmkoXzEz2BzIESIV7
de9VRXqQgLcVHF40ScRIKqzzbX/QbD4DYJGZj74qo/a5TNa/6vOogANO+pQritDRfyOMdwYcijTn
B/Z4Thc4hTajDtUqUjukehGGj91jDsljEjne0dHPi5p0V3L/REQrBj3g15D4H2xx7czYDVc2+Fb8
qdoJL1xrx/KEEPlfFpfTTdtLe3CqGhaP1poqnLWdD5i2XquOedn77pF9wPtlMVYehIE7NIVREetu
Ls6jzyrk8c7S0FVHjlNDVMnPRxgFlj29KTwZCnGvzt+OO2QRX+mroE/cVZW/+O+dF/mjWuPKnyQG
gxaIrSt+9u35DroXHe3A5/mJip/mHTUTSfHOWbb6pigiezVYuy7piJvnkrmayh02llaLpAkoPHS2
NvfVS9WNV3wMoj/GlnYYeVWHnhK9sUgNOhAqVbJb45O/dbXBmI3CBskxCxUScPFXII/5ul8ElDbX
Tk2xKGojaaaqR0dfHr2N+uw0MfTAoSKjWxRhuYAhd8HtIrRJpmAhMMRVywUA6IikTVSUXJT48oIh
VkGh+FuyI5l0BD6moUDiGPkRd+m4+IRQMZ/GsjDqln9JiNALNynedWKVpr6i0VpjmwtujUs/nf6U
u/c9XBWOrjzFIrLvLoWtgd7Xi2HFPfGXeY5ku3eYQd7i0VNVTGwICPPG9AyJOaq5suMBPr7t103Q
v/kOVnK8bM7/8HCeawX8B0WxNvULsKMPydViaTRMrn49Ureew85ign45ZUf6/UjycWq//e5pB8pp
hzFaYrtUYEpXyYdIcrxi4uSo2hukN1VJIcEGALrQygWiOSRDYrjD8No0/chuZq/ca9HrNzmML6Xi
NlXAjrpTclsZb6pakZj/tfZrnMhyOLh+0dN/iUIQN6efQaoElUY7X13ZiDQoFcfloToUskkMzyaf
eP/eb9fo/zCG0VWrEJqQGKwDVmaN+XbnaWxp5YstUUAtjIyICIhMb3advDS66V2YG21q+DE3Zn9G
1Tkej0Q+sUQbSazOmTxJ3AAes65mG9y3TGf11Nw0+fMrAlxpTzUeU3tAmAYJgoCCDDH2Xw1ISyz1
i0HXz7fGa20fBxRL96YvhH+8hj72jki7z93cuxOlxyQ2X1wagn0gnJ6r70dqIjDRb1uXAQlEXceY
4aoVuGV7vWUC9c/aS1fAF79KwbHRANMIMrNkwlhZyyJ0Cl7/RFqeN5Z/dC41eIhNc/3m3/BFY9+W
fhnienlzTyG+iUMXqIU/Za0Lkl00ChcXZFqdE/6jj8H1uhOfNIhG3SC6DxiH3Cm4FdfrND7krnIk
4BnEv9ld2QzfGtP4qGHyZdf4qeyGjtR0074PFvucBTGdPxW1TD4bfgiOizfUg2HozLxt/yilSlN1
HYBLg3A1uUxcnypOfnTJtz9MC375keBKkf7Qw5flwP8f8rw7HBr2cEwcorM8M5NaFeNkR21jcEf+
OzoWfEUf+Z4Pf2jYNkeoEMaTaF4RCaRQILx3AK+v9b9qRnIQ6r2DmnYIdz+ueKB7FENG4tJtzyRg
SQqHgiZRnnbOrIH2wPgFNOj1Pr3Rq5u19/X3UUAdl1wbEPiCmMKq+quMgrKEx5jH/QuMZCJijayE
HMIkOaC96R/YyVwac6+gVylY3ZQEfjIVog08XlDyrqR391ZVgI+nKdXBkmgvd1xMCERx+pnMi6zg
nhc4lwi/wvSWSGXdRi7SQgmLUDmi/ub9/SvqihUDNOqkd1CzdGmledJSqGy8ZNAmXZaHkcv5Gg2j
0mH5bZACbinqBiEcTlrqtt4xYlv7CrTQGI9OdA/6b+6onBxVcVh6YLl/Nk+YfyCozWdAP9tVZjwi
cUoiPtbRHIU/bjR70xK8To9GO8z9kmkKIS5A7x1T4z9Oi27AtD2d0io2qr7yfB4P5x/AoiChfLw8
r+0JUxajsfSksdM/Km0GxG4kk6IxZruwVitIkEIjhDUxRcj2kigaYXR2HtRg39XUxW1ZHXrshssF
kMumfdKhK5a2DvLq5/dsno4gF6HWVcLWJ+oSPsaZ1pdnt69iKU+uDZdfQSDZRq3ad3laePzUxpNr
nQcS8GrHsRclkAVwolmbZ0QSe8tAO+0r9SyPdC4YF9kKqsk0hx2ZV7M1Vd0ns2q6vRhFWtM6J5jn
mvwCZoPg54lWn9cCs6+iORJm4pv6gTfWupJ7YHnUPvfYVBaE40zi60sN5AN4RBBhiLvMP632jSiP
mol85iuk4mXtV16Nfk0WInF4Ol9AyBHgS7t0ulRnBkaRcE6mZtnb8olexSVW9RhFujTtMg72td/5
lZpJ/vXaUmX+z0OppwXPXp0mOmiFUxMqXZkrXtJuzzAvyNE99XToqV1gBSXARazCwJv+UOCj5sfL
CdxXYrXykDGcoPm1AUzPZ/p244FnTRJbAVrQCrq3jlkR2n0RtMIG/P5Wa+xGcs67Xdk6daaMw/jm
va4IORzHqVVh53l2fHxCqYB6geMTBGAV6n0Iqg85tm3g4S0mpZkIgpwNtZ7FlIb2YtM7GBsZ800Q
6WFiC968ISRYAg3c2W5sVmmALhANwgdHcmFSr7n7QYimh2u3HAjJoy/z97kmaHyxUf6apLiKoUWR
71NFn6/Aj0JxaBmxM6XbuLvaBUIMEjWuVEMkVv6A4uau5OIiFPgJkGBUzfk17Vsb0+YDcDn2yLC9
kryt+Yx1YF9qqrhQfvnD+Ap03+lNRYCjSjnQXZOhckhI9hiv3YUtJs2jrE3roTi8wkd2kmnehFja
e2psOc6EbwKDscJPujbJj3rqlZb0Ro7FmFoQ6KpiiVTgM6E7UBFqbeyCetszhwphtWdN1y7Vhtq5
6VOh+kqHJS1DCnTyZA0osextIN8oO1Mf/hhN89nmalBRAnz5auM6DFwSv/3QCiQ4lfs9lEKZLSCS
VQOTZn4B8iBzn7T6lbJ0SSsJmehjaiXZivjJvpKUSumOMp7KHI8MQdVQjBJrRMPft5m/MxldB8Bo
lPMI2RUZl5Rxej5oXO0i9+DvBKsI8oRX7HUus2dG4qSlF7MB53blM4vWLf0ajeKiaJSsICmiEHCr
5VJ7yuaAvvfiDIWkJbJAmYm/x/3227X4RWxgRkou/oaYyDaDEU/KR7hz3ODNBfxARC0rm07EAaEb
B2A4UgfrX3mYfXLof8alln1M/aMNqEQFC4uhi5HrNWWif2z5UOr66A6X8pOS7k7HYo0WG8nbIBv/
7vh+68WewGNTnR2eAbqpm9SDYvA6IbxZRbQLEQX+tl4qr1hdX0ihzdBvFbWsqDVbJ/4KZK9tSuZ6
eUhxw7BuIlKT2IEE9+uvw5v/i7agf9WOlvRlNLdV7tfl0XfSLfYDTbrPUdbnwSBlvAwo0IHqTBOW
7RXXOhUj7Ate+9II08s1HmVHU9BMSjLIaYz/+pZv7EA1Zpxng3wow+HiD1tXVsEIe2jjkDlH+3jz
8uHywFSptqo8bpBBqBcN8oymZ9wGDqs6PtKd+I0Rq5sYJ6e0bXomX7prQg8EkyusjHc0Wau94Vlz
W8JHPh907Vxj6fkV3CD5nvOg7bVy+Rcu9mhFBI1gArzIZnNK+j2rwawfRGI5FsDKyvQp1YpuimtI
JYnJlFg8+OPr4nb2nuqJ32E8L+fzKWKFZ/i1xG1rjPkKNxA1vxjtDMDp6B2ZODi6NpspsE/k6PsO
bhrPZz327tBTjW1fEy9+ak2B7NP31AWLGwhLyFBqTbsdtcWps+0Cf8BpyYTu1Y6QF6qrTEuxVJav
d8GqKv2WatycBVzW98+cQdaCv1d0FTFNzT8aPMTpvbQaRzMDeE9mU7CE7CV7+9oRPhns5pIznAbH
Edg8/ql2S6rtn+qzxLZGt8EZcqEVeKZiCBgktjn1CY8PkAAMhIfZ6QCNIHudZVxsGGJeeVSD8kSD
0hjjU12SWcGZG9ka1llBy2ww/kImjeGOvJ7OsS7ooCOrqWhelrE7gOK683NK/UW+JAbMNoxMsZLS
hhynAqAwjs0QssPsUsnsdc3jxYhDYDvyFwU6xUdKfZRdzD+pkXPSLKiTDB2jgO4L2zXeF2Eu4lvp
1G37lU1WHis+KEwBn/+4uLzk1WVTXd8OFWcRkyxo8N1Z4PIKP7zOn3fVFdOBlKlS4rzTiBgtP2t1
1tozV4Z8gVqBkAjy77ETosdWZ2xC9pUSx6AM5WmycJClUqbxDPkA1l7G93LfmsUIPkhlGR0srRnN
SkkZxvWJndQiB6GwJmdwOOl5+mA9Ped7OLC05PTTPQaygSs9UTX+kYPewn8EvsXEB0TsUw7LwGBu
dQ/AF37shilOT7wqjV34jHDZlye8ML4dVdwI9wHlZOcnddqbA76zqGjy+idRxWt6MM+z8R826fuf
ajOcqN0IOzA3CbxTg9G0iqTwgAdzKLXdd8bGrgj0Ts4+dOlFepSqFzbnsQW4xHutQZxP/Nr3OSlj
6/Ygin9NL4KOmE5RcPC4cP22TNWHthJuC3zRfZtVrgBHAg5lIkk5vh5wkrKo7riw2lFcfdm8btQI
v3nEe1x7vY3yo1Z/ll4mXhQy5GwJ2JeaUqOGoLmvbx6EzrpQ2cVwjGuxxA8nk9d04dsRuU7EGEXn
e4e6pw8EyuJ11gZDnnK8TsrIavhS8gQaqSNuqph02TJWqtKMSsP8hewIX/SEzR7hLq+QZhs7RDp/
vnoiYe922C5HfyFsCs9pEY17ci2ctOKHIk5H1xzPACcGVt+fy3IeMQ+yMi4Wpxj7YVkabbKMujbI
qQFFJrFJwrR2PtOqTGrOG7QwyacqqQ+7rPxBD3GE7FzhwY/tYbjPLd47WIozpJRZyGnfUXmyg0lg
SoX1p7/Q37eps2eqid6/vGK9dbfBU7NlG/MODwRpu4FM4w3QSMYWR7m+b3zbklSrKGjyBq4aBzE5
CQaUuBF2/1wRUBzs2Q2T18f8FQBsWq3/NjzJNYuhyxTPv2Auaa2Bl/Pwm1IPU3TEF0DoedYmfmiQ
CviHYx1ab/EA8sUOsUh6pBBWfXgZGImkaWL1F/apdF6f01h1pVbSBFa/cn4Y8df21KkNM/DqzAMB
a1J8KoG+8vgasz/PHx7SaoHil0qkpMSGwVVoFzFBtIJs70cYwPAjFTkQPXX8knxcXVFqcj2nxyvq
Afq6y9wEcJIeOOKrzJNdtMJKgZE/U3vwsXIgaDnAz7Bhk+kiGmAwOLvPiCsVIEMDse9EjK7Eueqg
pK0Gh5ztEn7NvD0QZXY6q5p2DWDLAVXtQ8fSQxqQq6MYJhMQKnfRd/e9n3Gt/AFFe0i8HOJGip/t
+whURE5qWHNk2azC13c8nRPWRHR1c0hvAmUIYaQzuvcp7PwI36jt6GWq2rcK4uDycRGl1eXA/Wr0
DU9GqX3r5z3eyEaFu8LxB2NqUpMvdpUK3hmcAz1iqGNCSXzRdyt7kWGYmNmNkEbJDN2OYJOr2LEM
9Tc9/FJ+kcguU3k5TAlyhl6cpr+sZhSdkwbbWD8Ol2912nCwehZPTsRnriWhuIxwJVVSyuN2qQeL
S432Q1oaRqAQ+2Nx7TXa4ISXJZbc98iJJY1yK3WfUXk7Ot6ksyA1uA9ArUTRpVRM30pt941rAuLy
+VzcMISvA9LFsS3O/hcLXKmKlK1MGulHjn0rRzTpdOCzM8UEwmLmS8+K5LosJW2+gTBKk5z9hthg
Q7LUKpR+lW60A8m6oO4P+kOPJ5Q+Etm8jQs0vuJNbhq7qdSuuegTKoPJ78nuQJeLV9aMCmDDl/wL
Xq0OH0hWlvhcIpZnPbHAS5JkudKk6bQjTlD5i3KuePeujpoV4AA0Hnkz2ahmi5cT3VkkpXn/x2Pc
CB8xF+lZHv4yrv0ztVpDKr5TIJcj1h92qFUjzmR3fEsOTXvhwNoDvXyHSpNW6Mio3PYHg3XLUzsg
w6CRLgitDm74e7qVhGPnIBls+YlSvWw8CGaIhS+CH3a2pOxKjUsnGiScX+B37LAHS3eWA0eKChj/
VAueoa0hV7u/L/3vU5bhMit0HUm6BdJXGsRneAz5AUWUGf46G4wa0ELhTcvSvqI4oLNcW/avxYiJ
oIxs50iLP699bCUGLwYql7/a/EOIMVeL5getLMUA/X/fLK/J28P2PSsIrRVKIZsWKOtWKNTB3L2L
SOrjKIFn8KRvcfs1Krp3mD+is8/vK6erj3r/K2YV7hTCHQtUO4WyGs76spWQDag5025VIQXpNV8S
ImWsu9UhVR/EeRmRxGDthuJeUziNRXI9FKQNuEta2UF3AoO599KVarqYYhB8zd2a7mQhHMFg9Mi6
ZJFPXj/NJd16s6aa2hXjIC1Zfj+uhzw8ktuT5Fcc/Bny4iSLYqFK3laFStsKK1T5tQClgGj2jSGx
DGCSJL19DxNvgsQATTNNvW2hzBgL7CE3gsbrzkWk60/daskxqCucWvRnv2rPKeqL+McH+lW9vtEB
ssfl+VLeRDlAy432/1ZMk90tzmlt3DgICV+VGpqXQV2tXF2UZS+ac22+Q6hmayhsTtfusTZC0DMy
Bt84u03z2C7C39MlO17D/3PQD9GAAXcyUD96Zj49ofQrQ63SJd1oHtPwkbTcrNIovfEJgYf2AcJ1
9QCBadVNBi4JxjzjzU0xCCNHqWuRFrnAdXgktig32QvWqQ7Va8cETMh5aWgyatEXmI90N2DLG+ej
oVHivVVvMvthIabI6r1brD4Vp43WIezkEp2aes6oM3NTwor/JJoy0AuA/ja1VxTR6otuxTx6tGku
VJfBJImdi1lMJFS3Oa5Y0V5VTVHNpBiRUzc6kgXcCVljm5U0+aMwCgLwCGbVP+quCulc3qsmLVAg
POEKBknOVivR+PaU4/jVp/ljOIjKAGrOSaWpvwVTEjFBVUmC4tyHqJRodeaA03EvvAlWfua9MlVI
+vNUqcAEOsca/3VOpwHC3zkSnQx2acw3FCnFMjLMEvja/2MOBS+gElrQQZDAuTrfNJrPG16Z9XwV
oREGtAEt/IYw5QlBaU3wySKZtbpS+WpPFmpAp3nv8r1lq0BBbRCcK9CNnSlA+3Z9vNuIfV0QcD3t
8mY36D4+/jf+rD/ctOtFmNgETk/uQXUbq+ta1Q83ADQPkck1ojwhTBHKO0lsVWszSduRiMuoPzIq
mRokDe9fykt1sLUq0E4DAO6FEcn2cmdLi1kCYjPX74cLU01US8MDwGr54nFAH8SMSbOL1MXPfBbU
cK/oYL8ros3ekNalp1bBgHX7F6m23zk9MihFta8+sAAFR3kppPYeHgWvwNZby6QvbNX6z6O8pRfp
My8AqsMd1BX21sWuxcrpgD9+q+eIIE0AGPeUP85yqgtMAqBrVIZ5YNo+rc54/8fyAvpQJ5hovbfn
ZqsTgdS1wztVlILLQSHphhMC8WETErTIjsjv4alG6cwjqMaxZ40wcFFDCD+q9aq2XE2KnkNjZoL+
7OsngZ8QSsyI/GA27hddSOWzLYcaKVVbjv7HQYUqoD/IKUNGGsTPvTx6hCXLlKdmsRKuEqezVvGy
GZUpZf/XFp32tBu2U1d9Mb2IE+ZyvTclwA+RLL6U8xSBX20JQuwKaxU4rdjUrMYaHTFHppkXfLB3
cwH0A/Jn4iwPIGphiLoi+TbUkPv1vKsycjkfBcH++rCJ24oVNQ2MN0NF/ybv9qc/3ussX8IpjcgZ
auG0rQclzbannLXXAcCNxvc2hNoFgNR0jVqdOLWkyCi19J4fNp4g4nFYGxUIIDghIZmpaJLGguGz
MjCQ/vhTsjXXzLarmbRJ4FJDezwOLF8iEuv2H5OIwDf5JPmPKmWW0NhShjgyh6H+3O1bd0IOSojq
g+VQiA4Fy8LWnyh36kSy9Rme3kPYWkyE9+38XHQSZbVbhDo4wwF9IXJRdabQq90PZ4N8MZ7ldRwA
FMXNMNalu8lP4m484OLhUEYnrHitmbGXkmC1WvuVXXcmCGQsEgOiEYMY/wYqt4P4VC1ke4d2YkMR
gpy2eFubflucUyswNV2/2cUSqLXq7MKtqZ19nlOCx+nFhu9Xua4X54fp4kSQSAZrrTco2k5YTvFf
F+Wch6vbnW7IZ5AKiVa/sA9n23t8KK67PLRDGGhlnG6T4GpR+5Ux77S512ZHUR7PbvUe2X41Q16G
9YmsG0G803QLbkIXFYZ3A/nL7nvxTsJMU4arirlRK5HO0g/u1V56ROxf44odL7gbQO9Hz1uQBWMQ
hwi51bY0fWi/ObjOfsYTGtFNYr6d04YqGFQ11FOy9srPKZW/C9SZ7lAVF0GFUnCPmwvxfgV6c3fy
tYM3Cn3j7GfsSvrZFXYNumJY1hjsnFvZeDCwH6/ijMhMcHXO/MuUEqzbAYYEZUBTolMtR7+ILKwF
DYYaWY3QrYmJ/H6FMnV6ZQhKiXSBKkx0PaVE/y2ac/1e98P3o68giPfnuWdhSsjicgwk4PuRPNoR
6TtzYUxDNQdPSVi875SgF8de/PQtu+XOhw4iyahst7dF7b8c8Bg2JqQhGrahbH6AMoTFcD+F42HD
An5qzf2UGbIgfAcWT+e7W6aPJE+LE0NdVGZL+yN6A+6VjiDyOLC90cFwHEa6CtaklWbBJuo/iHUk
tO89jSD8r6aK4lu5plbZobU8IH09clHLCZmxZBWH1vcPyxfJZ8UJRIUwiB/xLy2zWw0013GG8uLb
oFI0EQoA7lFEpH489BiN8qr9aWXL+AlHpJfagt43FBCTRkc3Q5mMyvGG9/KfZ3Pw3b8ivGjVkZVx
UZ7hBLZjRZrHhazn09zDkYYfA/KOkM3LiBRHEq66cfOcbn+7Rtsk8E0vVLeHYlX7ukQAeLoqJh8l
RWqVMRPNtuBf/0VDfyLf2+4QjNOwESaR6hHuhQSULxg9ARMR0Nv4F8pDBeobeHiF0zG8h6erbyLS
EmTu28bgLPaqHKBcxPY/Ci/gd7QknS4S3GU7DS2thxwAH+DukLyHQIV4vvTxnFZ9tjjj08CVVxJb
FmE1z68FTwtrHzjZ//IPnoCXWLr95LEisyFloLbm9NHRkuNMJe8yT+GSUnFEG9VbidCi/3RNBFN9
fCeuws5g6u+yBqbl7gNOKIu9m5IM36OnLdz5/Ny0XpbSRRGP6U7dHuBiZLcnelD8ZqqmahhWCY0l
DtZWfO2yMOBifncbynSd5D3xSWj9Kz/8vHG/XerY+AFCD0+4FAlGFPRlBSGQMO0i1lj0wfyJ9Dot
5lk5aQgPUkn0qEbeJPX8gHpMIJ3qIoZXcfKojFnfX/yvtLX5+tOKjP6iQ5+I/jmQM/eOiNeUMTs/
bzffKsIWHgI1eULO5YSpazX4Ds/2yAEF1cAx7zIZYMaQXyskbMY+sjbugIkpA4oWAAUxcLVksZOO
9WHOpTs1gO8ckrY2uHprTvgPByc1XfOxaG3MYUFFjR+tygzuYPSylA4TgDW3oyxtxnx1g+9+GWXK
rGUIjuYmItsIeQIoJt1XoCQg4m3Cbs5bacgYrppjYDTIsw+N7aIjo8nRxO04as4qYXup3KhxBNtn
e71Wp5o5RGahU2DBYJ8VKRZxutxkeNk3eWBhx4baG1nXevxYP+MTODMQpBbbjwElJxh9BW/1kMjC
5S1585cIQtoWYcH4C2q9QjXdQZTnyj5ZPzM/hnM0uMcN0OKnkrk38N56E/QMfF4Akdas2Y6KOyEI
XPj6sNy04AuS29Ba5RFyMeA+9cjRsDwYHFiCSC9yd1Jqj2YwYVelvX+TxnmxXVv8dkMc6Y8KEfPa
4eoDGziPV+DsVVnT5HFzl7TyQzxkWFz7QLbzbQrPa8UOdAo273aWfXIyXhhIFJSq+MZq928AOjV4
cPajxSUDlbJY9cBS1L6OkW4ME9byJ5+/nWYpxGfD9XiiiqZoVAiZcRGeiy8ZWmyjWj/fxIqgtapE
TlW3HFNyJOlv6MU1DMd9yz9i/RcwsQktzYkNoJkS6niARhOElwph7EnzRFKJ6rtRlj+5djy7QzKh
zFsDrSLAZsjB0wqNTfcsKHbM8KIoZlECeTkThEJXdN7pIjSIUY913tQ9Op2mE9cD1JQhP35d8HOR
CDgv133dtycN1181NGf0IM+GnoJIxuKuvUjtKSooG8XxCDI9MMLs9L8nAs4GWz2yABFbUjTZ2NzL
7fvn1YMS8PImLmDQawGngSLAFQNclh+TLvTWlLBhlMHMCrm610x9yhMCTLBFm2q2jzxyGVQQ7pPe
AUqfL9qm0gg+IJ0fZMnN13enuhZBIbO5RjHmgbOFKX+tyNzvLAD31hYbDMCveihJKUOrsRqI3Irt
KpTJo1btXeSTx6bWtNgMER2XAB42Pi5hSZfC8nAcYhPksWbur1gAovONdmzN1rHOl7LGSXfHlwka
u5IHnoYBIwf1d+FbN5Krs+RY3fsw2UbIuU1AwRy2+5oMgMEepOz/A/RPs2wtdGuHPzBFQ4I8QQ+t
LDd4GwHAQa3wE3A6ce2yK58wgnW3dqAzwradXMZbPtaBe980sARl8Qcst/p89kh8Y5MJSZ/++JSG
WCvg833HVIW6oqP9vPEztbFGW3UcnsDBaFWR548plHfJx0/Ac+WTb1RZt9hwgFlL5jZFIggjzcEm
dRWWU5D+vPFnG9ryxjxHCR9367dq4yIM1lpNuzJT6+uKsWWfyDZhSxmbbOXOePeZfUEFBubXUvvj
VKxJGDfAP+bTKBdonmJ4Hs8aEJ3/Zigs8Lc7KnZR5f+DrlhDIEeUGgdD1FUWqnb51a+W91eAm4Af
JrlG8g5RUIUuywXzbKXbv+fRN9fQEFysAm/662cVcAURhikJIKoSlOEtSJPKrjmrQ4fKYZBnSI9u
KhTmKj4WEUNWXOD1DDN4QbxNc5NvMo6g5Zc5LT/XcXNdKZGZ0QXVvwcc0wfPdrQVAQGG9OigBW+V
PMpW218pgzDUKG7KeTSV2SYs6AEmdej8S7TiJSqf3FfIfXNlLY0UdcZxdqbhSoC29CKb6gky/hol
y8ym7Ej1fLQOsxfL48/JdRpAPktDiZxGsDiUAyZi7fZ9G4lTRgNHW1qWr12bPpT8aBjzThXWjy89
f6Kbmsw/MKdQMtsCLnKhx2GJtiRcVJtpkVk3MM3SBueYssinz/ugDzcv6/ly5V+zclADaJEZAKN7
uuyuZ4HDW8xpQY6AQC/VszLFAFrPMMVt1HMCyYNorN755Xe+TG1GRODINIJtbnhj0bz2Ei64Q//U
WMWWRQ/5szduQ2WBWsKaP/ET3uWb7NaUr1hQsQXYR8/TP5cuRThe24y9Iep/ovv2/BQIR996LMUN
imS8srmxv0OG0fbrDRngsJVmgyfKuHau8GkXhZ230xDM9gO9Ce9JPOyzoMBgOx2XYELnJoY8swcq
qqbyiTVncexQFehiSxklgJJO3LomEuYQcSR6r2L7j4CFUrhE3kPXkih2MWnSmouVY/2pDLJ9RkYQ
2P+ChNgCObh/Gb+ln/pTtuNUvmcnIPp55izadWQ9mHzFzPbM6RfKs6lYSzGMXvS/sqifnAUNm92A
d4VS+EDEJ/AvFOkncmxRlcp5tpBID2583DDzLAVWqcNO3OG/ujcNpZiJti5ashA4OnMJ0PGQgCO/
+wDjsCqsnd5bQ33IxuMzOhyYY4oe0Gq/aa8XAwZ0R2L0pPFzpMHXpXGp65XXj0ZotD6IK+1dcdI/
o/cfpL8iTxwZrJbZF6b/U5kXb1V4tEvoXZiMHjl/Grggalt0GWdcqtqmx6YvtDIDeufxNtSCyHq8
et/IaiRK3nyJpihlvz8ek/VQZpvACJrCk8x1LZl1jxc2wmOeiXSQ2VJkPGf3PlHrtqVGylj+xLAv
B3r37v8QnugJxLbIKJqc0ui6v9GOpGRn8lAOHLT4I3GDIbl8Cqt1k2g/Fp/p1JXq1vLfSxOT3A45
F1Dsphg083WcVW5RN05O37IrjZ6Q34KvBGGOSFjKQhGwauig8E2KNMxx3w+BWhC1fRFSHnrSyw+T
RId9+wyAKvlxtqu9iR0w18UO02scwuDMIG2ss2xrAAYanovYaSQ2ZbJfoKtnp34JIog1ahUd1QwP
V2F1ftyduYvwscrPv7Ma4yq7YQ5KEjh8cOHjQAkQrx4U1A7LSTJmnyA/56DsBkihDr5jJy+ql4fn
KVPB0Is6SbJoVf65nhOx4WkGpvIYrGaQT6ysy066BLqez/BWjUIE4HFrZzN7zIMWn7/hw2aeP45z
yvnFRJ6kVjHwlZNZfldiJLdpDkfCM1h9bBfr6FoWZ3GSbIgCPzGaGTvDalOR87EgE/3D4ZJhdYoP
RMX7+wechS/8d52+6pqKU1/d7tmqH/0MpXA2O84jvlBZGAyMCmfZfX11d+bvr59PfU4SP3D0BqrB
DnnuBTfxr56trXPNfzHV+9DPVP2ZhEA0/UDl/YYHhOPwjoH/m/CC1fICkZStkhlnwJPvMo+cJHCx
iQ05jLo2T7sLO7JAOF2cnzKmQSX6uZSXcGOXM96bmopW/izrF5GeVNgW6pr0D+n7xHarCWGidXrl
mSBbJaxoZM5uyTBXUB7WH6MEaej0yalo8jB1CVftFk0+RHyP906X4lYRuo1uR7S935ETGhIvj3gd
pFALoFttFpCNSuOHRX87mUO40fQi8zUKkFqTEtJ3GpnnDMYXtzhQMwPSB+prNWQ0x2/Z0dQuJ1Ih
vMHD+fzWg9H9XSxB+xbXzCqvhtG/6nP46FZ7kM1y3ShEbyOMyEF9OVH1MidQ2c+aL/Skf8KAze4d
MCcMhBvAar5FbpIOk1AnFNn6xhhCy1WYe+TviZgzU0uOfEX+6bzP9032+XEiuYafYeTwB3NwDb74
jrKgFEPXxNnekgUloPlzkyfrALSf8nqhwhVixTj1tm0jfsaogYKNEmu7ZHmZ4NpEC5F+V9DB9qQk
6RwPvOh7Yo2DPKJyXKruc+piwlgLjhrJeUCsOoXZzJiFiIPaIAwB8UOeJPsAaAxvxxMjhuSlzdQA
EXsT1dHn+5zZ17E2hYqrp5NnF8EW8351llcADU5A1t5f8LU+yCSOHm6JQoMqgeEogcYr33laP1KQ
Xs8Q9zrBC/tAoqNg+lCObEBtIan5eYeze5PPVpnd6GOpZzNux5MG/GyiI0vLcm6OYpJJWHYWp6ve
dUAuQ2A/lygmmSu8QWXVqigfMyAjzmSR0PL0OQVDBQ1ROtzrSrRfwMiTioe/R1eWAbg4iQqpC0Dq
lpMiQ6GB3EV1IzIKMo3XeB4stWUtdoASbROID+iZvSGCU7D8rmFdpzw4B0Wfg3tkMHBepInmNlUC
0/Yh8+f3ZVbsjNLI5ntiYIEuNDxjQ0NkRxxTQrn7lDCNbqXGuz8PDu3q9/P+OlSGOE7EKeriCGAE
mETylQ7LBqEiGMR0fLpzvQN+mimcRKmDXN7c0TtD9G+LRO9nBEI+faHNTXrY+D1kJKsDlBYHpds7
4mwjAFppgyAfIodxsqE0nsMja3IMD25BkXPi4xzw+L/ngVDWvtAAPRsAHt59q0qCMh47kO7Td7dE
AuWmAJ0DJFlvg111OumvbJvIpFom2DNVb9SsP42YpDGtPKVeBGKY67AGIjJqDigIEGHMhg6WnGY4
y2NRdvEcX5+rncP9vuQP+wc7UvdTSQyIgCtI1fELskElPYtjZ/tT/1UNVo+duZ7Ym+7p6r2CMGjC
HWdipQxp/UEtUBqHbcvaa8Yvi80uy3IkHumPyGqOmH82QUaQANH5B3jo1pvdiL41rovJ57z2nYqq
DjV0mCkj+A4apGqj1siyc01oDRWpBkXGz93Kfz57zoC4DaCtaKVaMxXl4PTL5o7Yykmxbq9G7ETx
yeO8x+6W1SuFs24Bly0f6DJ2up4DPY6iQqL/dEGLLmc1tSnKh/2PBVDGGugo5PZK5vAESFmInAhN
7rYgbCZQwouUY26OqyDfOIwWvHSaeToIlUrBNzsc4oC5SI1QMl0q9y3LMqJBErhLNtCH1vsHOkAj
WF2pW7N3nVaY6k54tPKubDri0rglYRRoviEepaIGCK4DMCjo4niD6KoR8uMx0v/v84SW6Mt2Dxrp
Bh0Y7VT+w6Z4dcS+KbpmySld+GjizXWBhQEUA4ajUYgviCxX4S/I13VVyN+m4JMV32ytKFaCVSE0
xQvWMVW4N3HbG1WKSsZb5xKnzAQbNvDx0aoulaIybluyhgTe+e33cciOEyZ1nwGB+9QRV7uWl5F5
JKCEV4vkfnpMr1JMYDvx49w2n/M+pumKRWmGgwEYmJqmvghlMmLhp6z5AxVbNhiNhApZ/SeDZ49B
FW/NxD9e9qbQRq/1zvtOYVB9sJbCAhK47Twao6IgUFLnd/pVhOqlAV/p0ExNs/onggvRfG5T8E2y
12z5neuXEDqWv8QF2i7X8RcRfcYqNm/KRYnN9ai/RgGkQ4G7BxgUlymNrlra5sKxCZRvtFjQymoZ
OGNUpcJAhg+oPtFMkFP9BA8NlYFj8BPp1xO+Nkn1CFUDh5SESq/RxS3RJkgqHfJiDQjsY8eeP30r
d043wb6r7nDi0oAtL+cxysMo9j/nZYPGL8qMEZ8QEj/bJ/MOYJkPQEJHenX9jTTcREAhvdkbToku
JfX4e4X4GueyGYhdwfXGEQLrFzom/hTF2+gITyE20TxoLytbmrMUQRcFnemEaxqDcXkWH2W9c9TR
/3/UQh5sz4C9+3YyqXb4XKNgzTjxl5EZDmmNQmtaCM+wW5tCt9Xy1hOjZ1xux7IXsmLAsYVGIkG0
ZfbdNTxkFJ0wvHMFAjEtIGBcaHOd1IVNXF5GqtD7O6QBs/BcGaONX1poStA/WHw2oAdGIQVHjlvb
ruuhD8D8IbKUJrwZLqXtYc2dAwJhakQmxEuwRpDlo0Dl+de1ycsdPnF83HJllmwkWAdtMLPiARAd
6XHNFZ43makv05oE4IUTizTmYL1IIh5Jvt3IeEWNOcAO80dVZKKZM/+pyHgvmdjQFy1JRbI2aaJg
28qm8bB/6oopaNZwSG0lB8u3ekWxuWWW+X7QNY6Z1StwUyRPBEFcI0Tm7tvWqclKIFBca73NE/CW
Wwo4jNxW0AUM4ZCw2gVric0RNF+Eh13V45fVj0P+Ew5WyzW2hVBT7t1RV+LHiqze4M7egU1JTsZQ
76wmTSj6hhsZtiSj7xRB43ll0+zOi3hwXmgzdTs8lgSUk3LyiVl1PhCMfa5Xa3d7QVmYY0u5tYXS
qn0t3edVL07Do19inMSBfiauIAD2YRbmaOB6AU/IkmP7/jy3jZ2aQYFTL6zHWuohegw0ySk1Um+7
WwmPtwaNaBZ8jqH6RSjMsaVsIZ9027GIjNFRlTFZ+E4pXpg1VXxt+T0bM1rOakF0R8ABlJDH0z4L
NCAJ01WJjMhB6NDT9GP5zFv/k56DImeECM7HpJMUCwKVBjBDUBTfwCyVMZMyNW8mlr1cDr4d1MLy
45EJtuEheDZkrzHmdUjMRuEqcd6UODK9sx2HE/i+J+LLgYP2g9zwjxQoiGiY8GB1dUpLZn+wI41K
mgf+LEQxsYuJQaUchvGaAayPqot+oBP+StOUzCnJ4bIfjWDR0h7Kr6YkPZqigLbtxWVsbExXTEeC
/yxUotLLkN2pe+EWaMOO+tAFBytXAet4IzfoeAXEfIC1vnE9quaLSC23RnGAJjeq13f1BrU/1r/W
wRyOyImyMjehPsOOOk7M+8x3ZgyQ2rZgZ9AfF+1KqZGvHxE8vfrWs5Mf63GRO+dBkYUp9DZP9XyB
5lJOf47E+zDlfaqcVjYikII0nEwXIvVvw+ztQOJWrmSTx0eAakWMNMeEcucbrtNj7iZ2Npnho70n
T1wSfpu2F9Tj64X6KQxSMiyGkXuhIJBTs/1jC4sTdGMzE2WUgc815Y0zbSqZP2kZ75ZMXg6bbfJW
2xS74Icl/d6G6IIR5129DNEFO6SBR0wHosjGm8Fef/gY8eAkifFd9AOeaET3+1Y4kPMHQVFqSadN
XYsfNpq9eBZxmJ50Lr6p61w2tjc5ECEyQ2r306vm6b8ES6JM6zZsvTAS+1aEynCCjyUeRidGqTOi
HYik01Xy5WEyT7WTf26QCyiz696QsPXPihDtJqRx2kqUMtG8ARNKaUCs3sRHdZD/fXwxQuIpWetA
VDIZQAxuB6SN8OMylj7dezDjc15wgSY2uo0YcNfDghdQIL7NarL3ITuHvgkcf+P+eVuRgAbQ2ZYe
bSp553Xb3dVvKkFpw4dwRzrnw2hzToQWFRqbfGexw8+2mHFvg/aeRv1MMGPoVjCi7+PsVCZeG9GL
m3xDDBXYB7tGPTswjU6sn+YAeNTuk6vSnwhdFW7Z/jt3RGEZTxKvikLDkbZvJZT0sRGFhUu6LoXx
REZX07xQm7QybN6SRSL21Y61wd6drreCwtpPqmjyHDZZO9SONI9nNj0eAag4yp5WSGWtk9MGQpss
kk0HtBDtinGvfHDuBeoCsmn002FtY8vK6SVJIFz3mCbNAlp6GsibcNszk3sNYOD6w0UAKXkCtSxZ
iVZOplzXKj0EbCzjvZoqC+easoz320KmWTvTndWqqsmCzHMk73++8KSS0FftQAqk7ymcwPG/zoMO
bYnD3nZ4wriJtEXRkOhIOPfqVCCXItIu27K0tjhjb09VCPh5v/nc+wyXwU58i+i+s20mHRumziQI
Ijl9uclw58zSbYOEoJrT8G+pqbIGkg02B/G7G2yD64aqlrueHsK2EJ49Kn6BP7fQNzD/TRaVoNQ2
PDoOa2z7NSzzkrA4PU3o6cKB8ZxhbnYl+Q2e771z55GWE5Ks07v2YcknzYLbsrrAG+coQpMaykwp
nqiNWeX49WoYqX/aVG08vgEWEIKs1G/8sQjq7K+3+CUKgwIQtf5HQek+/J+S3x4yqSR8FuQJYorx
avsh6NSgBmQFm+ycZ1mTVkq0bb+GDspMf3RzmpsngMl64awXeBtJ0BWyOyk40VuiZAy48ssdgARu
S1tE2pOoT33sED5CTVsQdgoKr5pLgChytF6Uxb59Ozk75uvSFRqTCGBvwVeoKNHmlI1pyxq4lWmP
EwDHlrw+oAiwOBVhB8ohGS7ZzMi9mYPcb7/1Yj4CK3aX1vvbBwzB2hXVjgVCeDSt1N+i/aO5/wXc
RAIeGJhIcwMN+JKjMyfXlalfur4KwRO0wJGzj+J4pP/qPFP8iNUCLjsMjDEvvXi+0rHcBDegeEuj
Hip8CVWdYiU5yVeLx7sTsUfurhTBvFNGhRfxQOg0TJYYvGMSjDR7aV5hz7RKM9iYOTH0i8Wrvr7K
tNw0o5Jm4ZxLVnN1mG4OeAh4hTjJrMTuXIS99EiqLh+WBfP5np4Ogulo3Dp6W00fWvdQ8zbNomc8
rm5WjZQiXdfACBaMIQV82o6R+xNEZTyfWt99vOZSewLQbF+xbKf6al0O1MYeAn+yao+LlMcFdQIP
EL8Q9z8555+QmZ3DnX//Ckvorc3nWs/1100DzVBBtI5hoDKM+1eueZgBeOmUY99++Wic8gjLRjqB
VCosdvsiDUgz/kJZsTVnwov/8U5ksnqUCTPHJRh2OD7ySjqaV3ZvOBAL24uvS16AtdnBf738H33g
989Eo52ScsKvCuPodxUK1Qbg2Uu8OpWFMvzlcGiQH8VJ8lI0d9T+NXul+BwNIamY4NYPjJVJRx27
KAccUYh7UtzmwsmKbJjwyS5/g7eigIb8SCevlHZZjjR4NDYEdm5Puvcp1vVdfb1Jt1u9PKrTUayV
LFyJ8bHgGttEA4KZxWPh1NWSxLAuHiSyuF+YWQyrMwTJIqddoWgSmBCEuVoL9TgibwPYReH+k0pD
M0wTaCl/BzQrCpUI11tMoyFJ5oAk+AKnJuq90HIbnsaZ0l467qyx1/twhET6UyuOc3mFNdXJiTE4
dApM4rK8mvNV/sbsr0PpyfoySIPY9RvD7ovBFpPmguaG7GwVhWmAuUYa0CPq9cAoHw73JuzFX9at
8ktXZLCTMNZdCFSfiEJHEmnVlBpeCBKuoAHntENeakSVn8zu0BkzSmGBVyvp7+7yJmBm8AJLQfPa
adMcir4NDzDEvfTpltAaqWxMSvF9ZrZiGkLTCUz9BMO+JMTxweu05QBn6OEn75aPQJTkx0DSbLVq
B0VB83ptM2/GEr9TLtfR2loO7HZZ7ClRO3y1F85eamzLS37eFob55BXu+oOMZHLuULoMILHvMuSY
7NTx7iF5KxHGCCsVitbgPrXnv2cpPJumHNRCTbFM0ByLEkgsuCH5oCVMJ+IG7Roug6EqwviULWjw
uAdmMgcOG5rXzj+W4b3Y4BO2wgMNXoSzRE8gPLJIu8kvmR6X3+blwJJVTMtFg/XOgnYpgeonTswn
k6fmt1g2GRnzETvdGlXKROHMikUZdPl5neecCOq3sJXlU4yRhRSdE6JLohvFjAD4GACmLr8F7dhh
g/8XyBvuYqbISnrCY6cBo0I5YgingCaNZl6VsEwTf0j7gWIxGjWSLU8qQUyTkhTxWg7EnYhvR4Ts
33tZq0PoCbahKhyJIi9oognhY4Q+72vxvrAQzGclwfF67gSmiHcMAw4I72+vd9jB3QRUePyfwxto
o9ew3hUY3D+RjGIjbIVlrNyyyPw6nqJZoqQN4QvaRyg83PhQljxjAaLM1IJYnwkgQpeOrlUgRCS4
hgiwDv6OHnvmHvlXRL3IwyNz/xfdBNdkboavQVJBfHLPTUgSXdKskdWeN6ht/eXUD4U9o5g4H15M
FnS4Aen+Dj07ymAs16s4IDdMSd84nLbdbidMqeGcrTs1mNydrPasOoNIFB0FVPBdrCRPdE9IYumY
MEhfDdmqjfmMo2FgNq+1TGzHrk46fJ2uUH2nD+/GUy36buUr0yIseLhh81ppOQff3CqAXU9gP4LN
+33mkXAGZa8+02gR4wKfwmYGjgdXHWFffc01lxj7PcmIFSSGoI5VzytEs4fbTnxOkI9SwGG5I8ug
o7UrgLRB3gq/N6skTlGcbefvwE8Ity7ZUX+6zcZIeSezLHR5TQ3Wmx2FkPm6OcFFKo7XzsrbC1O/
i0TKSVDIEpD4awwpJa0JI2dfiB3DkL4olsmleVvS5LJilo98MJaoHqzHWxMuDFrVk/zbq7XuvMdx
0rlMNRbuQw0UzBopyrKb55e56Q0Nex/4r8bKcQM6hOaclSEWoRd761xogoDzzeFw0Yp/+jcflK5j
PH9kLtzDJiib0EC5JSv75GfogiFX6V4IbE99YG6sUw61JULGpx9e105rcPQpgfTqru3bxrZsHDho
PEW4V1hGnex7Hkibl6UJSKf4DFnnOVayERvw+HTudwe95bQw7mdRs/opLhWiepCl9tN8cqoZEqzP
NA/IfJOYeE1Jn78Nok9Bp9DQNNGOz2XXFCgoz/U+GK11ujOrnksogxEFQQZvQyqsyg1FwzfN0/t7
eYWFOlfjkyW++giD6yIBY6v+FOCyDq2i4WD3w7NRunMX69OqRRgYQmQqh/ZV5nMNXEdeLDxMQdzv
Id0z3vJllo4L06lIsrxgk8+ObhRFroNZqyXFe8ddkDEtb6XeCLHnQBUHOFAZb4iZqY09uyyN0j2E
Jcz8nGZdhq0PGG0sN8G7boMCRJNnWIcCbHBUPI7oFTVBtPyaEYENCSu+xp6H8Z5RpAVwkkt72N68
sWKrn5uDob/ZFHx2XGoIYh6j5k1qr3N/vl7JVDZGV7u0GDFcmqPG1tr4KwLhzX9l+3rWRAsN2ajs
Nqng/bqOq7yIislYFuv29UgCfOqE7RLs5/v3z6kWvJvw2WRnTzk/uW0RpXAF7YC26eCRn+TA4Rrh
qVVgydCclw6dMvQsXpD1baPrI26DVukKKex7exAPeW7OXLsj4QmL1Isys9EQaS8tPxsin8RsSVhg
cpPit6zGwVcIamQi70Mddve+P2NgzNo2G9tt/ir/0b4/kqNiAeoytQogHVdSmxPxqZqyUO3AZIJe
N7bGa55aURNhjCKvsaY4roAGq2YRUCTFVZUQ2nTk6zaw8QjqNXxR+qwq1hSjiNV+6hyT5KLfYy6+
j4uBKFBcIX9o6aUvnISztN/pdrLDpQaqD3bBcNQ8XxupOb4gMMijAVxgK/BDM20cKCjpv+moCzUF
T3KgNNKTnl/t0usZpe/T8rJxXmjTkguX9GwWgKig6pHMIy7/JUqGJNukCzt+h3UFVUdYL9DmOlIV
RwxBOuF2gAbVOeJgAH2JHAwDAV2hBadgQbIsy9r5iyK9UYPyiPjPlOFvhRy7thZDrl7OgRuym9Q8
xVsrlH9fRlGzWNzto+cwgMif6uB1npQC3cmjhBh8jLXUIauHdzQFM/PFquf4lCjCz0h1tQnYfLsd
v1eTany+BQKC+CaPKBwcHcxfoP0BvGHqoIoIuOFQ8eQiKLRjn56PSEgX94wvauQdzunBtuI14QvT
4HDdZ/H5RbGquLb9aV6Cd+0XjQLA3cRqtjAyV+nWjxH7XJxdcK6PAWED+iQgUckvHuP5jeiZ7AP5
suhTKxPhKtypMJrRGpRj+v45MAMjtfeKcrDISdIf+sHFTCP/7Q+BvXXibPLHXk7IIbjiIajEN+PB
3SqIqqSyFLXOA9hN2pvW/Djgddtyub3EhXWw/lkZBF0WlBEuI7p+E9wq7utwznzUrFL3And9oVjE
cfqRELZnQYcnJAgY/wcf0UoriFxLIDdOVGjEwCAZ7BQyHtR00Kp3AtOKPi8L5ha2tNbVzqKF+nzf
eBYMWz/VOkca3r1JSwz597h4xyyaAMHgivAVpfG2ce5PFfKMm+sLauKKQjqsVhcH5aNEGviKjZsY
rqIDfe0vowS9Lp6NeYxCddQgZagLD94K+4DLE/G52khCbAgCgvmkADLD6w/vpPOHdtIdshpC/OE3
A/fESlcVN+u0O96aPHC3O7NHM1wLNQ8XZv3ruoDq/vWMGcQwyKDjT60psGQCZpc9EgB8twZ8uGrz
oFzOIz+AxraTLRuyUnokFQIqCePXa8rwyc45i6lInloG4Wo6lo+miDbioLEVbMrYIcWijCPRc2iU
UMlAgJ2pDfzwMDzjEcwKgubv8dnjkM58UFsI11PEq4GBwAc3mfJ0+bV6SwITbgOJOeR6+WatqC9J
CmWs5sDzwhoGXnhLSqNrIdzL8x69Kxld3lMUkQbke5+nxXiUKkOYYBoZETG7POnJ+/5d8eohdRTi
iUonu4iLsJyx/WLWqE8AmveWmjt3KeXReTxd73LiwO7KFGqEhZGYY8l2rxSexYs6FrFftu9X5FGp
YE9ENFZ/2YwvnddoY53N84uH34WyLTDKCnX608LAptAiBIswjtkyrtxkI/Zms/OHNc6A7JTe9eGa
dEbFR4avzuv5IReQMfRCOJXsDbskKH8dvuOo/VkYqnOFlSDyYVOkemybCXKKOnrEReOIMtb55+xT
tVyTBCwlrEDBaYWPAj8jTjB3S9eJORNagnRCEXwk9LSTwmo65kbf/fVNrNI5e/hP6dH89hPcg2DX
NZkh77OBEywCThtfOUAYwgUA9NKAcBDZOE6bTOGLwgLuS9SA4jPrB62Cji8z7IknD6NZnSCxxmPw
IajExwni2Giz9jIP9blG/qbIBZbZvbd5mbDoUE1+wsuY/4VozozEpzREiXSEHvU102ZWZVrOoWlL
MoYd/qphslcpP9/NPWkHkUYVVM8EmBSbV4QddgE206y4N7QJ458YlJbAFpYvJi4mVNeQoW6F54rX
VYKykiuAfqlo8tjbFbMLMp0d1OlHspO5KeQ+JAeWbSxXJM8pNH8o+DPjQGud0zllIWvnSgiFxmBE
iGaYXHXVg1lLvNkl6aM7IdzJOOgCTY2RG28szwkgzk3alayAiaDD1Edb3dGHBFNqhGmJ94N1ftSB
OiN65jcDxKJ2e9f/ulkA5Co7/Lm5rv93NN5NMkWz7o+LMUl0UAZjg+3e46SbZHMLlo/XhsGMv0+r
VK7aBrOgvhEkFaLv2yC9Ac1fziQxC0wUWhRGyq8FrumnUsuiaXC7m7Ex1i2vreOyB1fTP8QPvzCe
MVZbAkyE70L15vtTbU3oA6QBVLpTe7b6Fa+nqsfNrTlKA52A0RPTjqzQkcxtqq+TaisrbzEutpdt
YZPIOj5iGjpoj55O1mn7DpnxALHlDaq3umx+C03sKaAHV2kiDxuTIgQgdqD+8dbioXl9gxqaJrmC
FvhBTISjunWEUPoUpKWXg7kjGxD4Vuhe5M9mF301M8FcR+fXOf6YvlG7TtFyjb7ljirYvXq7OjOb
5lQu1CTyPUhLH4NH3c9u8ByMZjqpg9MwYUU4bQCG55s3r5fvtoydHTlEJnv7MxS3Y8RjpLR0QoBd
+P7T0/dvjrErNTcO9umb2X9avgmyDAR7bsazHU9rTLrM0pualxkwxe8GeW559eVZu8DuMU3kz++w
eWnHEi0FNuioHCLrFQjJrgiB15zyqKyBaSDeJQbkaIuAEJuTXT88ggJ9+oD5KsHEoqSvu5V7JEWP
mZF8FE/0NvHvtTPwe0GOOnrGUJUvoa+KO06hO0H1KOTFwyhKuFRouyxcGhPdyclM8WMMH7Q5YzL1
xyHFBqNScIXi4QbfN33bA80OOoOb8sbAhEI6i8hDYAy3r2kt44TDcjKHVR04RsfKdizoPZbjzDa+
8G22u2HbbAovt+e6LDU3zoqRktVLZQzEQmcUj3+k/dtKuPLLGja/z5sV6vT+VlV282TfdDD9GbNV
HRKZXDqen4q1u0KazpISlAeJ5D4dEocauP9NA11FYKoMGJUeQtj3+MOZph19i5I34Id8YILrJnDB
KZ1+8Ch+w83Iy2f0ZcPt23WBdOjFeef7MpebonAx+WStT0bT8ZHhscaAUC3NbYZDst8EsPr/iCku
6lPXieeREbDtBfhx9lUow/WWoG7SqvjOZWaIcrmcEk+piQkzVw/HMnaAoYlESy/4kuYSLLTitDA0
iqj290Jce1os7NW3p9JTBiuAZRFHjjsUBMhpREecUJdmgmrPowcDPjyoPVZQCcLSrhyRs9EIsXoo
rb3Z6afy2qisZ0hasJzzXwf6YVjDo1wEtR7l0ZrEV3LWl0emj+pVXuGkERG27i9lF8uh6/zqPQqT
wGhf1AOgyr3jWRVcEmMwBuZtpXN3fP/EY+sLibv6gwWcnaG4V1JpFRv7yolnlsml986pp+9o1PU8
Jdrf65Ra3FQtTpEbDgFT9wO780Z8OZ0S2vYqptnN+nsl+NG3sAiHmTUe96uH/H1GhxDzpJP/bgh1
FvsKjUXZifQF465dinQUEBM7qxwaUyW0+Zh355WKew7SsoBEgvkvVtk3og0kUlR4DYdDM8DlebDq
+dRV6V8/h30Qy5kEiB8wl7mlvaBAAgVbXGFJ7S5MWVAwfhaP1BNSER4aecBobUsUQNyLxiJ9BFgM
RV8jcWr+sMEKXAjFWAvvyix1p34+b9ElEgLmsqNZUl/8SaRtEpNPTq7dq0pgRLbZ23QXr0Ui7JYb
cBxRSnXv181Qu9j4A5rWbsWS8VLEVNTt5FlvzMmMF2xkNgeKM6A6cMaNfIMIEkZHGe7v7Rejinp8
l9AnzIkcDyZGqzr/+7uIJed331b3bDMzOP4NlW5uDtAGCUF/j4fHRqKhBlGWiDVixZt2lzcnRmma
oZiUAoT7AOvMFLhlMCgVLKRD6qk6C2poZtL5zyyf5ye3b/Yh9Tw+AsE7NgPAU9099zQUlORlnh69
12SA0TGCUU3DeULHecFOuBuu4j2yzYJwejLMP8wh+rOHFgr6cpqYbEe0XDQIUe1O0JwyY0oTJq1s
W8InbI62cJ7fFufrVi1/gsA7EL/n1puP7azoKM1KNzfmaBHWPJJrzeyd/t+5uoxMTHOtG97ciyS3
wKqh0/lz5iDzyytwwkqDCMP8oPTP6R6WxkzdD3LS5TWmOESePQk2kL3qBMO0l0vdx6DNIOcx1lOy
bJpUFg0A3xMp9gkDJJRoxxqi1LuIDpZbNTvgioV3ApQKOn/akhcEXF0BFYjYvF8rTOJflZBYhcnP
jydbezPHo454oxGc+WACKTRygdNb+/MSKGlTtAIyN1O6o8K2tTWGuJ634yneTwAbgHQPPNBkxjDw
z8EThQLMylO2x5GWiNfjVDw82cJn0AerIkw+CPrGeNi2sR6CTn9jYLxT+OGM9m2PbUx3CPrAEkjE
ox+nxU7UDwqjrinOfU7wnKUCZwkQLrmiPcmhp0aNHOs+S4go5MjqzEP5v6vCVvDOC9//gvJowoJr
W6Y9NJ0jCSq9yJnGg7vcgD3+V8THfyOnakn0dynJTK2TKnJwyBhNOFtqV6UZdBFXmtCbIcg3nc9h
IJ2ug+yq/62Xcp2zZTOPsYsOayZ7ntjIdz966mcKTCMou/P782npgSopcnQgCTmTEmEmv1OvwpBe
L5oPlOVf9NnFB9GjG55yPlnxYpz/Vv5y2NHDoFFxQKnFcvdm++WWoyciG7AGXSuUadhuIKyTioxt
l1vX2OerSBKyKFAfgpPgoRddGa3bVUaQOnDD2qRAFjBOc+PjPQF+u7T5Nsz8oA97674MrJTUdWnj
rpm1If4v0GpIhBXFN/83kLxECdeGcuCobrBN4WX9/MO0nibDZlf3mCm+OlynkPA8+/kFokC9DMHV
0jCo8t6cyjbJ9AFbceI4WAMZET0QfDS04MafN71rPcL3hxNXavWpdK8mYFdma5wz5+PW8sukZ6aV
GO3S8SRs22EgNRmDGpSCbQf29DAZmgq1+Wd8vslSQtIS2Ujae6VpiqBMD6+58NU2TZ6U1/IwrmBI
/afMk1++nB458lInGIhcqMpyl3rP4HeyQgLkCjj9IXLt0JLoUwxwBpBKk9NrRayXRJumbdaRQHto
cXUPYjtrCB9Txr3p+SreU+edaaMdIpjg72qNKjmMvcsuRlcx/nYrJlZhEn06XqI4vN40S6aH2oPU
A0+E5z5yeJefx6caHHe0KXbpTXDL4H/mby4a8ErKHDgmkB4cDGwI0U9WPwxqRRZiFe8Ga0w5QA1v
9G77t4BhKQToS144KvTd06rAtcBmLnwvrdDDyiYMk/rttPwqnFgalmjFI62Z1NZjFZ4mESUETUbV
/O9vr8KUZwTclXIqsxRfRaBgc2Pyj8WLKMW7aj8j/5nbQomrKXSjJGSibv8BBYs5PA9OkHzxpe+n
wLYJcC5NQdqwEczJg+HHd5m6xpb1/bZBEo6hyDQzuhWa0g3jiz3g42v9YyDRnC/6tNAOqw27mWIt
hQJNHgAOrZmBgkpKS8p109lgwWdU0Hz+2ffP/392NKFQwtWJwCoD8/OA83cRXq6zPnEYwKiR23v/
nq2AKG3gBl7DrIuFSAzXDgtXLcPni8OpVRc0dv1vVAAyLphtElHBQblGWxbfsrAv7Xji3LkHEI4l
12UonDbLEUde/sr86KHuD2w2GhRpQNohqGroZkjJfwMFx5VuxiOEjo51XJFFB7uon5CH1z20BX8K
25GLm+XL/2ld+zD/U4I4U3VGKL2FGbV6/y2anfhyAm8q1LC+hIOO3WJUE9naODow+usPJK9QRSQU
ONpNMeDk8lOUygu3ArQYof4E11+CrBGy0LzPpd3Fos/f+4zFFKw0eyZRlTzlKqIH5QPFr4X/AM5T
LkAhC8qoSuBaUd2CmS34xIcvezTsHsReP2Aelbhi8VaJ/rpMM9BsPlhIqYzsw+mH+/jyh+JLjjSj
4vZ70ar8hSDkLt9lA1UaWx55i7/dMpNIhIjKwWMtaukR9yDHi0SeKslUUAw6wDi54vSKJBZs5L32
ShYV5Y1jaDn0e9zGbwOXivI+g8kiP4pcHLyGbmgpJ+vjtrTY3t7b27T5pYINqJ7/KqfaXfvshuMy
2ai+bBvW62FkcqPlS5a0OdiJH1g9visa7R7eYUb2QGRQ79eRT2ZypsWH0qY+k5Q7qwLNDrVAvFRV
NBMdbPBHA1v12Vmeo09mZQ83rLOCuaPlP9jrN4qwy+MEFRxzY2Dl9TBsLn7pJSOmaNdmRahlD1yb
1c+Ic2bffOIsBguVunrl4K5eLdLLRTMuQyJbuPPx8EAgbDb0P11wK9txv6g8CoUuZg3v6sGcyW/A
kU/uvOfcWcQE8BMSpStg8gC3RiJr9IIhFDGn534ZibNhU1m1Q175r0IlaD2kuJ5tsyNhsatb5g1+
icVOMALkH5p8MvgmvRPgClAW2ZPpESTNwwzTLXtRxhRv2U6W6alKueei2MjrS6OWan5vYOtllal/
gI9t8/6AOz9cE2LX2bluhatd6vTqLLuAuZEE3FhhOS/LFw9XhH47vdQfWQ1WIGxykUBOOWiFdy7H
M9acDXMWMkNzGvYkVylEFU2xorabPnBiBSzvlmKQ0awBJdE3au4jqwGC6LeZsM8CpHUdvfy20Tg4
Atf/ILTdapS9nRGJmb/S7W+ryW0tvCq9LBwpw7gaKbpz/TGeL40mwG/aNtaRdm4/D2DXEFfjTnia
pHYzSnQJT1kieK89FWEIrE+szRIxLIG5OB7nDh4IftKu2AJW+kmhWt4AXaFiHEtDTSww5gJOWSKP
ZtYS5CuMinggjA1KMDcojMpDoYdMhu/lU9xQ1ndlZw9MF/w0jNFXuhn7Q+Wz7vlpu34sLbXErfFJ
AWfxXzJHJCfHQ8SymiNXaIfG7TgYDBwl5fKqXKSIe95nLR0c6IaPbZGLt1suSOV/1NbFljSiouc/
6KzP+rq2FWj5PWx/KY9cAVxqUxSWjEDoJlfXHSXhEO6SnsYLL+lIDukSquScC1FXnnM9g81bWab2
hr3sHZHLyjcQB5fA87hSVB82ISjWeBUJ/v2C5jjfEdnAnZgI/9oRCnrk9tcF7rbTpw/3cMEFcwGl
9k3Zqx4DLTSMBy1jC5j29Z/WJGxb/IFD8oyMSGDpGSFUOXURmdiFBHBnjlwqHYXNTq7EtMuW6Fmn
p77PHqSiqsgsgGXP0jKWeHEa/UyjpsFR9J5ZCKHUm0IzzbmdNiUbPpMnGJnt4xB9xQUxO5fpatoi
D03v8S2nAQSJ0Qmg7aI3GJGhNZ/fW7Rva7ohoEyarJpxGWIi0Gufik7PWCckSNsgdz08NXi8Pobr
aOg1Wx/oG3Exhf71/dvfusuIQzf9b7t9hd5zn4pBLPScg6Q9VeoGsuflSUmZmP/KYNhyhmMmn1iO
KiunEvHoyW1YMB8GglUNRYDjNagw4R7cssepc2GFm5sTP9VEzhtpwJT6HZ9Hi0Q8n3m66OHfivCa
9vlX4nbnNbHOaLrAXwBg7wXI9pe6I3wQh8IYW2npDLWypQxxkA+yQ3VXYk+jjNbN+zEn7q2Cwhrk
7QCFYv3pxGaZZz7BSpJwsuBUgJOiY8Txnt9ZBGNiUgNrDPcNK9IhNdMeUzTwYdbsVTQK6U8fcTyG
ifpMaOND/2EpnHo9hOLjOvWcckgh+SHwOMmGPlpAiCP8LZKIjhMRlDUEhuznuhKrav9qbsCIhhuW
z4heZQorAQjdZ2CXy3nHVaDQCHA5YY4js66/hdQ3niomyLRCfPNMCcTEGjfZWY5zqG0ciYKWhSDK
C8nXH0L5opXLNwhIugh/kKyvb7MnzGh5nuNUyx0o+baXkRZJO5Hp9/4Y5g8qrQNc+ArYHcLGpeBJ
CZ7myfce/ScpUx2j9ZacwJ/KXEziixer1FIIzKmO42B7DOyYN/Xsc+JC9KaORnOV6SfuQMKccqS4
cXKt0m4xVKBTjYq8/aCmPWrdENJZoBscCvO6OD9BHY9p4s04ArMenwHlavX1n90VXVCvSLA3Zo9o
TfXM6JOFD0Zmb63wkI09IYY7a9UErMshj3iRq0ewWBCpFEZpbsWn48jmo7JmK7V+6Di/llZ26uCy
5YZeZ+y5OyXbB32MmuDIuQATCiipo352HZrGAyvgAkIccVGQPKEmC652U4icd91A8YhKCUq5SEVf
+ZWhbOdoboektzH+jYpNztuxZgYueuAa8yN+CDVCwgbFA3XokK9w42NXSgYyMsSczHy2F2jKXSEd
lhEjAfRl7dsp1eeKIbTi9YjuiKS9vNDAthVb3rqqsoqHYDNktsjQa9oWEWkuietKS0siy9vDRY4J
ETClFjaUY6gJEmhB/4servC0QKyFtJtdco5RAl1pzp4RL7CI6wjg/OaRF0+PbNCv2w7GKZDbbC3Y
NSjPOjyh73p8xP8Y/40G8cE5faRMByILfN0xPUG2sF5JBplmrYb6vQUAPGWT8B/pAJFMiwE6K0TK
0tq7n3prw0SByejvWEEMBuAWJEtClYdwc9TjQAQ7Gxt/F1BKbYKSEfcJoYS9COm5yYoO+6cOSZp1
En6wJLQERUBEegXmgUmab12Yc+HMa2b38/CeiG+zF5rFj4KrWCaItO1gDSOeymWvwpdrauNW6VGn
3g2Z/Gfaf6AspYlVkcOSzp/9PMCM5l7ohM3gzhEVlRUTIyOXH7A0u3XeTKSwhJQdtO+cN1wrN3fR
/KnxY/Lq4KaY76OO4sc8D4uLG+YpmYnBi+g3P3RuLCdlLA8GsTREJdsBcfi4wmJ3IfkHKU307RyP
Oa3THsVUWkw+cySAndG2KyckMbv9PDgb0g0PfQojHWsrniFOsc89mEa4Cv3GjKePX4hfoFMS1xQy
pzM5J0C1rTzH4EEL3BPo1DU6yvDM86wuNFVfVeFJS6rL8KCcj9CcV04Zq3aissV75SH07M7Q8YcA
ZlZsB2MbyigtzijXL+VO4MmdGvo3rCwEiu9HFJ2azZrw5OixtSa7BiEkKPkY062oxLyQr1qdBSC9
lBrISFbwAQw067922pLHQywr57avXhcdbPsBsx9V5+BAC918tngqSyKV43sfBkIqdC46jSwoM0nh
RUIXzqcSTcMXS6MxiF2+48D2oX5nlyOXr8FMnBiBbflzqnLmAbynvAyrzznEEGvomwSIQUhyNsgI
TJlsET6cRkPddMaLBAyxWfqFdmEMkeZBcwcRzqiFiFkARP5wYGv2Nq4zOnFYuON0l04fi7Eki3N6
9fX/Eb00O9B62qWVqy2TBmDYqq4S2VCEbhuW8Xjk4NNWDDTROOT1ZunaGOtOHoI9CvdoJiJJx6lk
QzXqK8cxePQwl1nGafUbGM618q3i61a+aCbcUL+8oVKJd2tedmd8uzqBLlNl7RxCZkMGyev4g4wz
PFH/BHsQDAfwf6JvfdHUbLgJ+zMcCmn1JX3mgAgLsKebJ0oOPIk5d03YHEe4bLwTcp+41l/4GJPj
3iHEUlzs+yRfAp3OCPHxGb+izHlHDm/n3Hy66HOV5oFz6Q6hMhQjmkHp2mSNI2PNnHrCZ1+c67LG
I0OVxz3rGNdP0Epj+6w1LTwD0AZ739lZPwfHk1Wz0IKIyoKMUglllEjSIgiB4d2zM1+FCeFORwxQ
OrhbCfJZORDEtOljibMHjz4BQ94BnR60bZ8TRBKID/yAWEAhNWMYMfU9QZmp99EuA4UDNLGrFNzt
A/noYc6wglJDFJ9LW/egtJFtio6LW2krFfG4+pFF7ue5rhZchzbcMiOtSR3qcFzGBbweGO6BXGjn
+yQCblZR35RMUGNFJc4Krg+AQkaHS8ziYHrS0omN5ropL2ri6PE7N0tHlztAyujQRZPAszkne+En
KBK3Ue8emzkI371tNmWGNB2X4Qk3NjIVn0E29YSjUZV6TsUXRTajyTEJKiT6mFA02sTuoMNIXj3o
62Cr2iY4FDm43hicnbYTJfJrAXiD1aSa899JTC17Is224zAVn9b+t7JfUzJbV7yx55ZPeoCd4DR4
VyFF1YPGuecYGrYBH39LCLixFgmGeu58hXbDZdsbccaLsmFKXNIjojaeUh6ZGMAujV1T1toA1Cn8
+Acp56Bk+f/A2Nb2FYdXewhIerXO68xaVmcGo+GOpPX67mzcgw2DYqBzlSYa1jGNjDdfoaieaupQ
OdKf1tisdoUq79b05HbltAI2Lz+wiOzRyhuW3ujAwRyMGFi/RP3YkHeK99rnGXrk9E2zcjPWu/3C
/gwmkX32uPzaQIE7DLvz+11YHrcq+QkqRJN+8I2AEvVdemIVxLS4CwNiOer+TUFfmdT61O1M8XBl
zm6wQLTSntzcAR0M6ZnQORlvKnhuPcaSLvCzWkQe56mStGRjMKOPTbcYN4E1mQfP1FRlVG0GEUL6
wTJmZWnZxDH1b10NNkuR3tQ1cFkz63s0nX/28rtG7rd9cy5PC1yjORtY2aaerXHIwuQCZBuw3yjp
PPUE6kLwBrqx/MWB74GM/YH1omU/X7qLUB7aeILkV4e0lNJ3tvIpighiPLkU00heC6Hi4LkH57vR
n01mmtlbjM920yZAbLQoqbmyU/7yh/a4GfUuVmCRm13cDqKrJUkh6l+4sz1vTzdMYJ5/xv2FSwkR
9ZJl9V2bCxI1UEXwyHui5jSclx8n4sd5Pd5aP8K3CDRXIKB5UsaIBU5w5KY+XBznwQ9jlSqfRjiX
ifnPebF8JEGqSKtpQ7c/zFSsvfi/63FrUIB8ievjDUN1CKiH0npRooh+PjTZZ9tHfq6Y5GzcRfbL
DMjJRFKdxsAhapwDqUNniB82QGpIFQlF/g9mM0Cr80rWuMUxN0XwsbwBg6FNLACFF99lgsYPlpLs
VVBqWpmQbKLuYe8xjMr8g+DEeh+ILWoNy0/8CXmcSc5URa8KOk4KH/NYa+1ZgUow+/JJ/XqW3zcc
lnmF3LLENesDtidDE30mZZT3avMiD8Mi7dFzrg7KzVjMCxl7tpZmZW2polwXeQ9t1/S8fNC3XbDn
v7Od5r2Yqbi37PnStE7BSP5FKs8MUUC3PZ7aalPZrBTMD/8hPm0sZEAxNCoI5gHX5g4sqp4sB2XG
i+z0ateP5A9ubEPobuGDYXBrx3SirzxJZhxy+Y5b2iYTmKLHJMHJYqVbHczgZfrtZZ7lTNkgTLSP
mDykfw5cXlalvtkm7Kk21971gikXyv0uVdhhErBFez9y619LMYSHn08xe3oXHZ5V3whTqXXkN+ec
S2o/jW+VY3+BSJqt1SSKhk8dwfgJ5Tdo7xceHMS3SsDh0siSiUkd8EG6DfaqLV9S96H6iDT2RMDn
CJBC39UeQZVK1VlzhCd6zhrP+qDV/rmZj4fIPD42QixNs3zsBT/7Y5ziaUKr8/SV/KotnDzVqBg9
y2SJra34Wm9i2mERMu1Bb0X7rHnio4SHkIwMq1jWr3sDzkCbr8/xCqtLmFI7x8yQnJra8c+uRwGF
3fDjumdqK/aX1vCjcpIGo4l5PRT9eukIzpYe0gf9YTjDX3bomlC7qtc+9HAtk5zE95clepSM9lLH
tagTdgZ5YxU82I6Iz4rPhaTaWu98VMRuGDI2z98kFaq5UntT7lB7b/LbHOrYNzaSC+65DycCAOmS
gc0GIsDVohGtFSGhCsfZOLi9B4VJu2/f6rhk/0nqTnkSwqOjb2629s8gQzSlCHLzo/H69+xRUYnZ
qeBwpomScmF8A5dSm7uzOgnJnta1oO0s0rtAU7+vnxKsiozQIVdDWOYqRf6gPNU5/t9L/N2tKb3H
vYVy2upcLGy0byTuTlAyYDu/I+UVeLaeEDQH17FlRPIwzF3ZDEkz/axxVzC7o1Tqf0GNR6O37yuL
3rSBCYzPWA3cIuMvCBjCwmU6uvotfKCgu4kGxYDR4KWdtqDdse+xWac4GguH0PlRNay14ffE2spn
ycpz29m6w6BmuXZXrGKtD1nBBWc3h394cVmwTbswGBTHK1iABbhq3k91YJmhIS9OEegHQJlbUYKy
EFvTqgzb9PMjsmVnDIu7CY6RBmO9Rc7/Rn6YvtCWKzR5ThVsaGrjOsc5WMxP4V3uhVjKpBo5tyAV
Zg0JNfJ0vO8AL6Q4OssmVg3EYCCAkxMJLla3nQSSSHJobfJ5wl6NpWTBy4eI2ePzbXUim94hW+tI
bL/5EhbXpWbrAtzxQVMQwJIUa3qU6qSp1EJqg2GnqEtygCF78odj2dyqJMZ18AARl+0+znGj0hYq
q1k0YUqAnhiZTM1nGqEVeOu7oFbnNUiK5Al0VIf7FE8JVyk7BwehwIDrtf9adBDwC2zpQF2tewf/
7u1C3CE/YVsyisvW3jKlBcRtISwcMcuv5F+Kiq452Jz4dPGtKN5E9a6ZFNCYP71VryCrgfCdticc
j8awjY2AdAURUI3mAaRwpVV0ScHPefhIe2USvOwJdAMt91ZZQySkDqIQsu7OQ3yn4qSRfBkHRInY
J4fnRjMUrYbM7rpUJh29Bt3kOil1gmNtBZYXpUXb6hCUi69nYTaDwUL8wj1mM/hgTOYAGPMUBGFz
YfnrUT8Hk4eSVHLpzkEDDRV1JkSab7bepKHDhfQocQPSjTREUoznqUg4UOaaPRaRKp6DKSPoSq4z
D/CHP6unAfc6tTsaFQ8bHRoPsPy18U8GayZiDtmnjDIJPeLGKnKVx+KmiRw4inHz174bQIR8PWVw
vy6ascay5Ot94/inJyfxaNpabyC6AQ+fhQ2z8HawyQnvDWBHG02YxgyBchH/cbLHIBvuu+CoQgLt
rJcgaVC3jbG3h8fAtcLj8367uDY10JtLoI/Lc4WdgaRq5jPtYBtvNroRbAanr2zT5dHHUrMJ/WOB
2btsEe6iVklaPnHg5KalehyBHNy5q9pX8ZzOuvkT77Yl8PuCVirdsb5F0LvDUzPeqqwADqJenBYH
JCfD1b5PDnuQHLBM7/jurOaSKjnNrBVaDu8rOoKU0SjkdrWM4LufgbUPwyRUiohVLqoCW38lRlAC
GT1ek5J/zkO9yhJElvIi+4et+buby6PFtPikEWPBfVbInet10NuceRm60rMc3iYD5wrmCSKWldKq
okZ4Hg/jLMde2ryG+tnS5NQASNHTTWZGmCrL400uyOmDIM8Q06ci7MYOKORUnLX4JdrWfKTlHVYc
Ueo5IQGhniGIF+dgfjBqtF8kYa54rK+wceRPvpip62c/a3F6v2xK8tcqrb24FZgwYBnMtTxJ9+h6
iMmsswW9uQLo7L9UAW5xm4ke9H5d0m03cwzvYSQ87aWPzRTfAY8oYc953cjF2hymXQ/avgOY/U/i
qV3lmiPyFhjIx8GwMhAcFOEOFA+eKBcZRlHWqAPxd78y+0k+01X5Kh+PEUykTPRlEEvafNk73J9L
UUNkPrP611vvoMdGtD6r4qGBXHBvmuxSbFWPL5432IAoPnWZc87I80/i+l4xEpQQIE/auSe1UTaW
lerrAdoKbOeD186E+k/cVq8iAmCqx4JsORlyFszmQl5GcD+Nej0UPE+7wcJSsG42NgjA/5OLT0Uy
GvIPK5+Bx97EW+5KTbZ/kDQJ8STdYAgqjPQaFoNJevJC35oT0YlxmNRkCPSiibkQ7VK0b8L2ITrw
4XMl5OZ7aSdXhOkixbFw4FJZKOuK1CumTH9Ww0liZasd8B1yTvejo1lcOymSGJlZ0Hm4hTTUpnXF
LbAx0qAuDoXe6glL/Nn4qVmhFhiLGnXh+cuhdKHR07FCQ3LSD/eNM5CxyWtvb1kI0l/Ej4y3ChD7
qRySDimDGZiIZLK3qp1l3BPUiH78QU2U2odXdVBn8CZJYk5CClsSyCnMhnfW+DvkgRFWlazSPG0k
RCS5KeWYY5XAfr99THMtB65BjujLLaxDjUsLbS7j9LKCgBUg84dlnCN3nA08YiQKsKpW4lWugQi5
GF8dyUWx6WiL0/VgpEz0jqpmSlwt/JUzGEc6r42jIviQ9e+SrcLRgNN/kJzI2NtuqHLgb+iGtZ6H
XT9zovTK4s5366V7ss0iXS+FE4TLwlQUvvuvi9n2oZzNI0AMvreTv4cI6JGRefGAWMkeuL1fowCm
JM8M392vf9kg27Nf5omfDGPS1Nwh/gH7O8zyaANqDM5QwTm+m6g1B5kFJndZ1oOTVikHTTzLm24w
BHUm0Khgfg+HBnDFztznw0yqvipnaHcmgNA7+PXtOA3+XHREQLTfQf7Xpuqm/koZD52AHSCZCF2/
ZLvPU79nQOhBETRo2VNuy1sHwnn/G3+Qd16OM6kNd0tvQ4pS62VIAulzXGe0/ZhzNpnAcC9EQAS7
kLJpGWF4VDbQXdF2SObwz6oY5ZoK6gZrH/Ff3kMi8W3tT4GcxF74tLfjaXXMMvuzzmnNQ323a0Q9
VABrNaEaEw++13nbQAbiCzPTMYwlgIEISt0OkgMlm4LyJ9/CA9NS5AWmPrZSlZ783CyVYYEVpdLJ
dhHZ9WwgxTD/wBxHgd1IP8qK1kYHGh/N0cKHS26EGlg+zUQ2cT53kXR4rAc5xD20T+lliXB/9wxP
T/JJZQK37hdH+q0AG4so1MX53SUbnKdp6dXXPJ7E2l9mSVWYUTcPbfTmrOxJe+86qaqnfLUe3GCb
Ivg0yAy5fYGYFgx8x2t97fJiRL8/gnVnyIk3FfvWyhys+Yrryf63WihwqjVKn3ijqwUM0Pk36RCd
nY1nEU+VSRqbI3TY/KMM4iOoU/6KxoV+WleaZSzfozAXSAYtxypqAvs1KXmx/8BvgN/1MX6XLk9j
6EOVEp7AgqRAXZPI1uKkKtsFZUOwMsaD8RwdxmirINuuVK6Eiuqu5OsHXqcWjV0zcnbAEbpnwQr9
556IBkIgyKFqoEJP5I/O/9kqSwelDaQiAgKu2JppqCp5e0/hwKFWsSAz3LotY4kAE5ygDPOWds1k
C0s/Bh6J6/n3wV6/iUPdtwadzl6aalx8Qe8X+lcAvJaDGzSqGqoVfQUkfDv5Tkfy9CcKK6FH/pkQ
aPMNNM59F6qsACEUuj2RO5HZ8pcf6HJDhZPFkmdvDzgwaPRycAbTRWmVpkap9r1+jJN2VNrfw37u
Wxp9FIyHMBtQZkexe3zJx9KnB6x/oHBTZ/z+NMA1HDvy9k8hDnOie0KLgYyhXQbYXzGqY6H0+TrT
5xB57GCFCrxNeCF6ywupe/U7prnU8AlA3Wd8f3Dm9sM6K3FiaV4Smb65D7u//03aFtmsXTjXL0ZM
deQiGe+nRztw8SaRoOp+2oTPJ6U5tPMOU2G3fQ7KdBaXKMB1is7NrRb+EZb+fvYx5furZYgJqnPh
8HwYgabsM1BS4+VcC+hZal8+ffNgUzKg9O6rNmYurHkV0RBnG2nvvSkBSz0RSYJQSR7t7QXQLH5s
3gfA+V9hMvRuQuQGEQfaYKklBQIfEwAjBaRtafBpYv11YmMfrZv/st/UlB3l54a/rOPB/I1lEzwu
5YnJO2KMxib2WghvMtABzcRFHO/pxMyD+ubrpmcGbz2aWquy1tbB02nns6DclCLuzkU3rgPPz7GH
lnSHVAPhSezQnPN8ZFbkyirsaT2A5+m1KlugwqUXjBK7tPPatCP+WjQk0biC+JcHnAs3ft0FGJIU
O9NvScqp6yf8HUSTVubyA4xRhY1qD8QBxQWD9a+03aCgqC1oFOkH0DmuldZ8aL8q0Ez/ZTDYd/2/
rSacvXlNVKULeIcuEgvmNmXkPQy/MObAkY8uhEeQVdssbpWeV2xcjSPZd7iIr9IrgzdKD5LI4xLn
tZH0tBQUS1ZROd6aw/6tP5WvHnD+T0nWNCxQjpv5TdHgiQue2jr4E6gr+n9atdBQ26C4i3mYeUPR
SNZsugHunJgRLfc3tr6bGhkirLqD2BytFZtYNmG8nOjf34S37m9lZRcUZ+AGvO2v2/fmnnQN1XyT
1IkDFtON9al6V7aOcqJXDVhSCA5ZonPzDb6MG9JcrKWvt2wcY3FQOM2yVy/wn+swM/8a+bmLNiDz
6f8dWH9bn+7h2M+EjhvL2jy98udB2ctyMjhSX9PHlpp+JZdo6JRjl1mAXsIlYIzcDWc+ed698U/k
OgMb4jbN9GMre8AMfCzLFK8KjGoCjwCAV7TxfXqTi+W6F764t9w0DI7HkEbhyGQ2iUDrbBM3vGeW
tA/feaKpoLbo+91e8qpS8E57gupaRPORTcnpU2VPIDJW8oDQ4J/pqNkIU3Z2vzVTVg9sjrZ6tdId
bz4LqJynv4/5oz3rUSkgtRkxogO1Y3ZLPH2Z6Xcow8VX8rZ6HmaLoZMRsJq3GY1Ha5iBIkQpCrp2
YL6icAqiUWNTTcpFHyGiRjsyBNwj10qVRztdEihJxwbx8Qsipn30p+sPRop71M98REJudMmuZuQ8
DuuWpmBdZAHI8ntR9424n47cPRN/+i+kCrAHsPoTGKtl3LkXc/tch2nDVslp+wbN0u6c89aHn2OM
pgqAjDnBRlyIxgQBmtEqjJ/XC4cBqBnOp5YzUOtLiK3wPA5dbaIxsluZ/47OgAOi7hBymmsnwH/M
bghqhsfjVwTcoQdwTBPANfjwjHJzEV2jxJeF4V+7y/yBdefX42RoTPMPHTFDeDKl09lTpDlmggAw
oBD3kj2dxf/tKMtH3iHr7K6M7Os62XLN7KdG/2ZD27ZXK78hx+zhla0RUN/jX5Ex5IjBuQ1JFSSu
tfve4iF4I7VJ0JBkJZQtUgIkYg/SryRS21P0cCPLAzIREyG1wx+GcUylVvx3lzQ82E/6NFHumpLJ
wL0VF9wrGVRV69HUX7U8xKy0Xxu4pE+50FZVhR1vM2rTBz/v5xr+OiXshHg5qK3xPMyJA15lthn1
z5vmW3t3TEAxt81WVkhriYX6OMbiUmD3eBWmrL1mxHyPvjlWaMwMPW/0e7yH8V7ZO2IQmZ1PHzGO
KnA+iMvV7L507uSL7tKh3ddV1kHKlUXlL/aR2hfl4/RzZF8zZcc7Op74KVNTT5uaUsJOFM++BJxZ
zNOEnMkd6FMm2BcL+VraSFypCcq70yySWm9ygP1YelD1LZ/TAvvGhMeEYyX+ch4NBmRPSkGWMmuC
MWaTt3s+bSO5N9B18nrnYc5xUDhN2RtnyyqI94q4ojDNxiA2MaSO98LOwySVso8CpM/JpSteg/QF
B7uaLh8mo8TsQuEPRCVmfgnyLNuMgvIFAPvgbFpDR+oq4CXBLbSyUlmKyeEOPhb24toMv1/uOI8g
LI1OCiZq0Fv0FEy2+itRDVua5SJsW5Z2wVBJ3tIeTtbqPpzkhDri3N9uOXmk/+OReBRZfWjuoVgI
ZaVSfAJosoc+wgxRBViDgzSLJPPHxvZPRa4hVuHpje55k2Xew9W6DCd+N6Se5Pv85Yx6hsgW4Wly
g/NR/kfcLa4tg3NpMDT00Pv/Hv9eB2eqIfFnNLBy8ra8luGCgO/XQbyW7EUNIBIkSWmsGSOeFyeR
5m/DJYVrRyxqxq5V6Tc9YhvsfbUmsCj6PRFq1/pdKTUa4UBIrrhV8X2FjzWBQU+KheH7xmKps6Xm
v6TFa3QBljSas34qdNMYPewen35Qx2enHqzsLvkN423HLMBRrxSUq8egCFNFqtWuOTcvuKYNrT2z
BV8ECl9NA79N6nihwFATNkho66G/juoKPPVfyChg6ccVO8sIh2ejk3yCribz7QvIKTWeUJ2ZpxMT
8Wz3Qf8cXrU++d+VbP90RxGA7ULGzJgCTlApr/2KEJXrubkkmg6DI2vFmkDqEQBEyk7wdL/ouwLp
5nOsTMotANj0KvX4kibh0jaJMAm2jNaR6GhjcU1thdFxO475dayyLRNV9LDktTinmLj9DBODHuJC
+OhpGbFPbRN4VUMDJRDJWyV4XTkOUIDA5p6gp0aCfXnoCGxebLyGXtwZxbcvc/8tYsjZnPMCGq0l
1+hTQiU1MLjCYdtlab+gmaSzH6DBfoBuGIjQ6JcfnDC6NRjir2dAyk1EWOd2w7zgT6KHSSJqauAf
/HcPQ5UKCjCAMA4uM1g2v4qcn0wSVQGD78y84OQVZ328rNm0/M7xlqwzqKonceSmKSE9Kp8liuBu
XYZ+LCJr+tD37RpU6wYwi8uo3MAZxdV2JqhjiDxlm0KcTlzEGch5E0zp8E1+OakUnI2Lkod2ZXKH
fENL5SHxDBRxUFCwSUSFC4RZ0BpWq6MWua73Ywa7d6FkU0YB6y8bvtlY+QZqtpyj4I6CRTMsaCQP
w80bQFSTPoCQQnzBWsRNqqtipLoPk0SyZPDupIDqN+6saX6FsFARb7vBVBb7h/CTLGfJevGbGoFp
2NWN2PEJkbpc/rxwgP4HrtdXqrRXD3YWnB1buVMg/AR27BYrNcSqI8yfe56Eo4NW9r20Ko0ridgX
4vgv5AN1f/uxnsTbRHlVf1OKVJnVIWaoOLrkknC3Nz6uzFm06FFnRM4CdkxBpsDkz9dl9FQZvCXc
JS9VaEMNge9nTf4YhkPvihz/ISnEPycg0+Nh9YDDWS+rjCq3ai5pdVRmDDHPMdSgj3h/JdP71SOQ
7txbA8Sbx3bq1kMf7eFKFMYpR4tXEj7xbaO6PFYoopBpzYmyzgrJO3yM7TwZtzqnx3KSm0aT7hNX
nUwE1GGeb3UJ/Xltn1AtdYL0l9pnAhP42Yn8nWoJ3f7teb1mXjDQ1ml3gj58Y0IOtVlyZCDp4VQI
XF1079wOTClMqHDzPyEJTa46bDdAzFBgiizx4Bxk5XutjINeb11v2klh0u6ozSuo9qk5VfhOruve
aqEYq5vYYYMGWENl0ncJ5LYzmeKcsQqF/W8ChzoAOOqJusyapfZr8Hemsp6YZzygvwi5hBF2f8LD
QE7kW5KyFUJudmLJH9QHAappSmcDJgtBXa6gCMji/3yAPjJ8QJQOfbPxHBEVkEa/jIb/AyHhosUa
AIT46NKvkReQqPsd/uuC/6fcRZNGTs5N0UxPFd8gNagVhodD8PV+GoMBD/RRIo3hvgu9CBhPtMBN
MWpeNeOETo1zfQqCdXIh925xEancEvKF7Tiehw2llvdHqZ1gsl73zUIn5i5wyXkuKXryZPg+e2pr
yXdb74/ZJnRmE1tzsk7ocP4JGzonKqXH5n0dWuZ4SPayrWGnUVJDwqxugX+Ph4B5UtEvq4Zl5+m8
NGWWjaLMa7v5nEuVXTiVi2bXVQ1iSqdcCBHjv2xosuYURGLkEPrHHbzKyGrGRPw61/7gYH1MVWK/
yPM8T65zqt4x8Axg3AxJnGugl+MbxEQc/fDHKvGNf4swVAgbG9vhJi4hE/aa69BU8R7GCZ+/cy1X
0NLiPGX1m8DnY+6EEAYowZyCCXkK/AIZ6amfnjYxEXzQ4qi9KGsg89fgKpdRi+0jdIkCUtE2I+Um
/PaQUgsN1x8hQXC6gYe5bshHseQyuEtASVtv7LaX6GPijQCL3mR3Y7eodZZEFnUoQ76Koq0JP0hi
hGU3IgB8GsTcZSMC4NppIGfeFUUyt6WLpzTeslG5d+QoxwTuW2iVcv1WzBIEq1XuHFZ1jYrETghe
EcJayE11H4x/1cUywfvc2aQtKcHTnv3gp0i9jqwNvLrHhucMB/zUW+RsQmxXOksHXIsd3/P+It2c
0VwuB/lgXE4EWOp6L/0yaCTDo7rS0Z/hhirqvHJAQxgLJhEZbnH2gEDpzu7T5t1iTl9Qy31vWMYT
MhEGMymi869stQVmXt/9g47eMuCpoeGhhmrkAHVr5SbyF9nP05Z5eW6aQNN3HjQrHHgeMyMHJ9Vw
9P3Bh8iXWXyq5MQione6elFoNbEMh9Y7vXPldbVuPOc7ixjybRrRkfoIh+3iUDsYKAxOtY9M+O5w
jPVeMX3CtKqVIc2VSD5WeHJll+f0i6YajFt7LD6294+OSDR1q/UYzzl785dp50K7tC8Sp/btrmqK
9SV5UFEPILPCWwqJWibe2GEMbrd8H+bCwOgTHA4yKTynlB3oSR3SsAESnfA/rkrQo2dYkEO7ycJB
DtbpFt1XoYu1fIOQdLcCBuLQPpGhvkBmDD2NIPjPjAk+lj+2aKi3bQuKrvUFiOSjJIg8I9sh9W4u
oWJFgvz4JRvY8VAxpwmlLJ99WU1BaV9cfGa5zOZKuiDoxcoPrdmUTi1OG2vF0vRndAYceUomb+zc
lfNyEJbPnxnvPh92nPEz1DX5gp7C6Rrqk069YIG70Tk92UOZnGoSn3GQoneGis+XIM82C2PfSNRW
XOVsRBlnuAQdEnKECFwyY//lFIUKSgLktQnA10eyDkl/u46Ifq3O0sTZP0L+yO3jdG3tOkHeDUBS
QJs/PSmr7D6DF9MhiHmjW3+XP1hlg/YXxVjSMTljwfIFAB0221TnpdHbAecK9JZHJgDStUyxkXyQ
EZ1iQ8tQHV3HChTRls6xaKG6Oz9zJjZ5+0JYml5z74gUwznodvhdnRixry+q7tweA7eFnBo9fp6e
gFXLt4khfpEPaOsf8JywEsnEc8w7ELGZNz46Ii4fJ1O5dSaKBA2GcRo5eX699nVld9s7oxXsqdfi
d+Ik4kJtZC9TPSii8TMPYpsXWmFO5q6qDVpn8ktSXXRdeOnSeaqKgKbJ2v6ccRYbvoPatae9ThQ2
+8zFBpLADUHrV2WvqMx9uANpM2YQIb7yhLnQs8uJZKWDlx0ygUvEbH81Y6Lxl63QmtSjinSrs00S
D8jZqHqyfAc7NlMpK6XzxfS573Rv2lf1H1XKvBETFt5JTXghaA+gHY7JNM85bSphhlM4oNyh5GzM
peAu9UVnXwFayYKqEL9vFBqvHP3wnJXqbse8lrdJeqmYUqum9AOwOlHPPJ+66wVTRipj2mEgRjaN
e93eL1Wzzp2ZKBjfGtJRmZnBz22OV8CjIVyDuAW52Kq0Dh/h80/5fjesfbJWVAY4s2gSLDwCFsk3
TTnC1g8qw5InX1IqedFOuTgmSVbkQXUwsPJKLW1Rwf8N7CNFZqMrPjXX6sytVwutjF1uGKKYFqPP
wND+GHKZ/8Tv/sFPoepcLKuCKs2dK8HJFqKhyPQ3B3YL2FEYPDKdBpOx+224Y0w/jw2Ha8bDvxrf
RC86B/Iu+dK9nRF6VMw4F47AlejYrgpAxh4LsBcTJY4B1HsJhSAM8PFjhvL7EyOZp+iVrUhjOXyO
4N4sQUGpADQydf0vYbjuqI1J063aYJu/GyC2so4bOLUS30ln6xlGZuoRy3r4OPmypD/bIKaoXmSV
qsEBpM5PsaV6k72d5PHJ28VOzstEZAsi6GZZadsAOVny2+PIryvjjFU/ONCdFg6lfJEEFV9Q0ZyX
P6YCFJi14LNid3n8fwSHPHfThmj/e6BWujiXz1X/lLWVFJjwdXTQ/uVmR0R6Xf8AnPMt+U80jZcN
4OgTE6WsoHDkt1K2r7+zY+FZrVcfwTH5D28oSMfYpztbfvTmuVEK8WJS5x4yN9NPLXDzOA6uDF/U
gzxezjT6qtHN1PWWh3i9JGlNVzKuLmpM8E+Xr4dJZgww36LvKD047Wf7bmek3mA1wVawW+B4NV1N
f7YF4PdXRiHihC/UTvcKtbKDEUSyRKSFPkUIeZiJZ/MpYQ1ixVWh7NZnWNtFIB07cf4bVflGpHtb
IUAJ20U6fjxHcrDfYfEcwH6cSRVyxmuPnalup1niBrc46bBsFciFXYVxGN36zO380Aq3v3b5PlvS
/47uz+rhdgjQafmEl+zEHlzNsvakLdf/JttY8lHZMVNLTQWU7dwCuzqToC0I+4t4XjtauI8X+3u4
yszJNJcrtxuGEwak8qn4M/b58qeUNNE1vByDAvTG/a/U1pApQLzb0s55qFLHTw51gs2Anw8sJCmD
WEbQjeox7V2I/aAmQotTsiZK0KIsOyc4DJU8G2MBGeNskzUFz5KAs/S3ynYWY4DHav7PXQiCi3n9
COQCvQFco0inhyx6rtVojvG4I2ewh0LH7HSxPUMh9IogMe+qWimqFCgzKNzsYYbeQN1rUgQ7mjB1
3T/JT90loxvZeTi7a25s0wnHQUOkWS7l5O46mU9iPu8wXrxsJedWN75ujFk3E6aN5Tc5wUI7oheD
OnFr+6BAe+KZGoB9qAH5isIzH9wl5aDTS8Eai3SEX6H9ynmh6/Sav5gDijuAkNRgrUUPabahaqIp
DEEXxNfoWJ3Ma5n4Xqrbw7BwkCHem2hjCR1T5QZVVzz5CTRbOgAjvPE5l1GfTBlkcMI0sFIJZ5At
TI6tPU99QOks3X93uaHYoDftiySQD6Y0AQsX2Ct6D1gIV7SR7v7JUb/x6ZODK6A0qiW5YOHbC83/
Q3f98DE5Wh27RzKk83U7pHR++4Vvc8QEM1Wj5LZ2lI6V2zmzk9xWiX0KjXe6lkhvO5TIh+i2m+Or
0qY4sK9O77TTFG0+tn9MVQ6XwdVcHMgOAm8pGSb+wiNTr2VpD3fFOR2tGk5/hnYn8Y/M+RIySB0u
UiRt+MDGQ5NJvx+QDNfZTqnnQfY3WROEI0TwVPGe0eX4glBrpOpN7Lj72UlmyHMYBQgN5UW4Mdv9
85KSQgHKOWxREinAO/1/mtHnefO4ydKDRClBlj9thkLAGBeOZny6sPsIP5lrNkE64u4P+nKLUb/S
KXxfa+N8b/uKhUNpWLI5ohIqtZBOst6xcscsbQuCW2PAjI6j3WqEHCgZtk+l7ySU+8G/0L93OY4W
Cn9LxrYKUHkYzXp5brpdomvHVFzxoQrQwaH60DtIwIhvE+Q1oVZTRKUXr9vTNB0qeUxwsXlAOwYr
ki0+LBiPDheF0tTGNT0XYzJ/IhmrdJgCDSvTFbRjXzyLaQlmeXWY2OWhRQ3s1CD4wOCZczczDMik
Eu7yZ9VN6x+HQ1GF7zjiXCmu5nRLVwu9cp41r2/JMorVarQGhYiMXdqle34haxxWooEEwspT1PET
YuYqwKzw4rvfW3KL70ZdNibQMiRHZ3pAZPR0v2sjuWFcJYkrbObDtCF9tqXLDkBamyBugmKPQHlY
zuPnTiMmRtH7KiapqMtSaVelxtJ2UnmB3J1sdIyQ6vF+9iVVB+eBPD/OP/x+gFQc9jK0XfIvMPnz
3PZrDVGx4UISZxGQyS6Vbjk50WM99nvCkaqZ67pRvKMpD94M4Zzs8b54/KQSx4Vj18oqBVjWffkg
RncXUIU/6Gq3n7/AmwRecnfUFFBSkwbr+Wcc3kam5wWErDcifRy3V/yYAe4TVClmXzg3LwU9IbkK
8HpO+jQhmy7LiHm/7XCZYFeJ1GlA09/zzp0+Oz/w3aHH3boW3/tIgPxpKUb6+Vua1U4vNgJgrHKQ
gaMYSC07at0d6JTZZNnUYApxd2dSXesz3WXsFhFvxX/rD/4e64Fnfg8wiLtYj2ALoBLu/dlheK8/
wZTEHnDsHv+6HHenxpZSXVMek8GxDSPToGPxS9bzr2n/aH7dV/4e7bBQmt7s2/nnv43ulLFc+Pes
XMIG3kz518pDka/VzDfW7SAFcKBlTitk/wLRFqRLXKWrYFIutB+l2mBmW9wZj2kW3ypiuC16Eofe
S+aj+9xClOrzrYgqGdnWcIyZmeq/8MjpZm08qliy4R06Bhx8H5h8euIW8F4X9D40ooio/gHML8l9
WuZr1P++5jyUwev8uqRZKi617btS8jmRrOisxGHhezuFNxh7Tt8qNah9UcQ3e+A4xVnp7/j8AlaQ
BMQE0QsD4tdz9eEiq4SRULZDV+90PmZPqO/QOdEvSpgwLBuuoTg+e4kGrBM2fZj4Q4UOL4b9UnUr
Gs5oiq3jeNZmIIgr52FXJck40G79hdibPWQ9YuYSw8dFSfp8NyqfkZuau3sitPIks+X7aY+7EDUH
4C/CxdMo8eKmUnQq2op4OPcpRQiJSMoaPAGaqXoL6mJuYZv1r3/sasS2dofJaxZN3vNZusA8EJZA
6+ZhVrguSUiN01tXEa3S5LfWAOmOAWsbX7WdajMFZ3TzhmlqKM/gF+uxaDLSExeSxxBPfbB+5QuQ
5XfWx5EYaYosPpd4a59bBSivay7B61vUmdiP61B9SD2kOT4udfCJsrLrZH07UoSPH9Il1rFdxF8q
vwrZkbxwsa2qLfLnEl+83G1vLc5Z2n0hKlHCjf4m0dERWCQrAJFa4DDc5kicT119IzqosmUJeBOY
5jD1tuhnqZPPUwBDu8OFJoCyJsNSwRFfilTPlbk9ZK11i7m8ueSKrAPR6SUMtHOD9Jkq4NoUeGOt
/8s5EURpwVRr47PO6GsTwRVDZQs50tS7Txenmv8gog0dI10wRn+DeSPD7P2tXkUfsNQxecEVxDKT
44HsD5jzbDOtlU09aV3PtEdzPz+Q9OXC0Z1QWh2EQ22pLVHaEsidy98xAGJ+8R6oWiCMh4176Pt0
hiZm4qGITrf3yjrRwFmgB7PkpzNmPP6OddaAvBpI0KCfsN4Lrlsnebvzgrl3lQSs+xSHj3sdxcV/
38Kqxk69iJ2t9gYwEZRPSme+slqrqmWmYDmnjL/lSwmT7NQO9nacgcHhbSAeYyA5qUlU02InJHqi
gGlBVarQrTw5Y1W27XhOgS9RWbCgr7HN7xTstvI4wBNV7TW/pSUc99rD28ZXYgwaqEk4DGf1Sv71
smDNHk8d8ChM2Mym02r4F6E75gr3N2iYaNcWHtFqCM9L2mTtEuR8UF6J8WTcTXL8iVHM7Ne5mFPo
rbvsYbDO3pbcdVmtyBC8Bd/8eVveJ2bQfZlhAPkRt+GzTlXN/4tDQ915FxmhujB//4I4HaeWGZbc
jT3qYYCCWmMAwRTVHryWA6L9HkcHTzECdxN6XBZTr9RcUdKUEOh3xDsAYHa1xHNPBdG321q8vApY
yjKewXbtqujcbtyIjAl/AWTM5cfEQzlC/J0yGx8XVms+Pt953ArrVFKrICnCmIoTr7K71rjTnXGW
s87Cxz1x6jWeIajHZdmn0wNSwmZg2jc3N70dE9M+j28ln9UecP39tP2h+MndPPhvScLC/Fzz4bdy
wZ+SmLa+hAc7fKWvTPgxREqVvoN8aBxVEOguFoDqeiQjz3duIe5dTl8EPJLkvIKOYordFhC/4YjN
tgsiefCSvNyB9q4I1QGqdZnKyylTgDEO928rDSiheeCoPCiffpEYJHz54w9USvurpwUzETUZRREG
30eihV1Vvzmu8wY8/ZgqYBx7/EWoabCqaQId18aHnnXXVigmgR5VEp7FrsRnho+gC93hx8ON9NRV
0Ma6flnpWJ0xtC1DxwqT3bYUL6p9ySWcvdWsuZuEyngrzdDqVkQUELCJ+gNcJPr/i3+HRIu9dtZG
F6cfMx64CB4UUnWo+hXb651zBl0OxJJfMqwfvaemRcMf9U+ulFmZQl570OAKlTigj+hHXNRbFtsz
8Xk4tNeYSYeDbeIVWZN3xus+jYsAi4YmgtIoJzY76VePJ6aLjMi3muSZATG61nkeCrTDA52mcfNZ
NNwfScqsRTaWaWCosqJ5hIoB6Nu9NIBO4BUlVEFRyB9HcfYPyw3H9Zja/ikTan9KpZysYqz5DiXc
sEfm+FD2j9A2BZZuIre24gK8a9HKJ0hO5H68yVrSaY5T4EAteLcM3dGWpWrkT7lQBUCYLWyjSb+d
OtDeXB7oe2ref+rfbCwqkbX2Ki1AGKaOdnaarvdmgMnDnFW7B01sMk/ClW/J8dYy/TQ0EBB86kIY
zWcQ/3zgDsTlbwlWnTJkMuD4bU1FGV8ePrT12FgNE+TrntERqi6q0F6E1zBw1C1z2Y0dCPffKla+
9ij8ZuOkWR1Fwx9TLUNJo6z7EvZB6R6a6g4g+s6VIMNTalF8yJ3rwnHCw8ZV5dLQdTS35ECDhBG3
XBDWCTN9bCyfeLF/+e41RdiTI4+BN3Uwbj9ByZFTUpHoNke55XxirblgvwnmZ7Hgqj+4JV8wKv2i
/vKHZrdXVGmd79YrvyjATi6K6g2l1owyKcj/imGN50Wr9MAaBYfA0CD8yBvU62LP/FJrcpkWauil
1dZfT3JlRVzCCvZw7XCjInB6sJW8+OBlUs4WGNipyFoFuEYM2TlMTyC89Zmm0AaUFwot6eKTjWpa
gB9zEFzfgISAD/yW8/KD5YqSwBws4A+lBUKyIfBmQWITu7e4IQxegF3bovKh+xEr1mlamN8slWe0
nEYV85dcC4vk26lFlWyOC71QskHQdJ+avxODhdhVLENd++Xo44bZeO7IaQxKx2JpFmQ5cinIBR8v
JZWsvQTChFhH/HNNF90oaxQup72vTxZnzNHsfXH6ETb5z7XU9w8XI2YE9PQ6LmkH8igshgIOGGBX
orvqp/B5karvVkn+M0QAl2LV/cVxEycOGiR3+5M0FZICQOVhrNOWLgPH7ksN5Tjq6FoatCsTvaRI
6fh5FYANQHhJFLcGr69fhURcMr8XZUzvIX0aFerzXxnpHdEQ2CnixQ7XBSWQlz6mxNXquQK/VoL+
1VBjR9LuLNGp2AqjiFu/4grDWzwCqYoUbh3HoIITC6qAtVX9p7gJKMvjt4L/oms7513D9SzXuMDY
PzUm1z0j5MHtZVg75wiER8JbMKX3rQCVRntXRIbWXv3dqvjAkAs+frMLThqb9WrMOYxnEQE9OvAI
nP/pvNXWsnGctNheSlvvTbhJbf7YuPiy2Ltj/yy3m94rwwD7E1Itc2arvMAouN0f06sElNs3iLRV
8wl8fBLG2l6NgtmHZ5WG2Lbn+dFkdwie7maylTEAfHaQ6ka4H022qlCJaaw7YOSX7wTxUFpU9bfe
DmT3MkIaeEKn6G3xuLXnON02dBXWQ+QapM1a/6erDm6kx3ts0uxG7XufzVz7ADhSBRl3xI6JraHn
Xv+nwZC5bf173mumpg6kRV+iZA+i62G+NGz5NrA5CTW2MHwI0X5i+AlVOyJgaXJl9uVc/JfRw5Wy
Uub9b/PSeYUfU9O6BLRmj3jOr35idfHDeKAhaSGNlU/1VD2Y0uPM4JkMLu2+sdjLUJq8qImDlcF8
Jtral3oEVIsd7BYomZsrxY/ofRJkLw0Fm/yhhYH0DwTX8J0U3mcZu6ugg/3Z+GHdZsMkBGH/tW8z
/868C5Alsg01WLYsVl+7ihRdyqF5lSbdLrdIIKjOU7gVr9Nc0HuL+uQTkgw468RWWDkTFqthNG/8
m+kAqALWYD45bSTy7elu2mjqvYp1Nvy6Ul3LSGPiGKXc2D0KWZzDcyZVtPdO2c2Hv8cTNVXyZ6ni
MQka+sFTa9zxbqEWmy69ueDvQeFnvIdwEpQ2yCjf7x+1zgWA7zQgVsJ/pbNWLXPpuF7cwVxNMvlU
DxWc5fQO7xU5AZiy+YpGeXY/Dpa/EhXPzwpb1S+W/txZDpHJnUePOCtaSR9ZLDyZJp/YqAnzZaWg
8P2vtwPqc4mLxGgM7XhfHA29px2GqhsMMxWKKVcH7jf9KWVGjV7MuNkJLS1Bb7+K4rE83iurvpj4
PIXU0B4WZGh6n5nqjtwg3haeRY2rOob7xhvm0/yDGie5rru/qCVvxcXQj0Eb5ICuUdAH1Cp2yZCf
OUkERrEIjebhMzHxsxnma4K/kpIhF9kTSitckNy4NavDGs22YpXUYf4a68j1F/b8B/E56fVrCwtx
FB6e5jq0wsbBhDdHmFtNn3xIHuJpBTbb77NWa1gYTEnlSkl+4jabX7JKmXVChqbBeKcHPoEQoAuM
6K1CFzBgntTQzDWbB8/e20iJFVJkDa5GHLYCN96kSmSTn5QXJRIp7FpBCnADp8gMpV28k2N+gyII
04sC8oosyPfRRwLAYN3tlce9joLSQ3KLJNLPi1J69P4leUrxdXGnAwhdDLBghQ52ve6RDfd1SnuU
oYTRDZX3LRMpReWlE5PcHHbzUJIn/d7r1vAPkCt0jeytXr/Bzd+i+/O8gBOaTmIABHeO4BzJ6cSn
BOlL5F0XXCglbQl2+j00k4YXsZZFj1tD2QNLX7zmf98VNY4f1RdfKyCnnTzoLoMV5KHnSmVQHzTP
KFoBNMD7FdSRd93TUIAQ2nG+W9PVzirqP88bk+FRjxshazcc+5OnDvsf70lLTmqeNVBqVUCwdQQp
nreN2iBfkch6H0BXeCPJHc2dQH9rOBYChNY0kjlYacf9zi3Yb/HFRoD+Hy6XtoKDWx151Jr+p3bG
w3LF4x+MPD9sBY8G6qaBVUq+Tp6YFhgxj1tuxtfVezRc6zsXwJm9tmECD6EyAlrVrS1eEIAZ+5jW
+LGC04S4nboiZwzWmR8kcyl6Z2jHnAeCKcveK02Q3dRPm+Iu7ycgsuqFPYvwZnZRcfiLvxIv4Z+c
04Ulk3UqTkmkdjlLZuJUbIXXoJDQfTD8RldrdHoIY0vZ+GC8OEvFw/KNfqdJ6u9QXI+AAH7DoTKO
a+V7FHheY5urANVAiXvR+GkSGZFgpIUbO8wf/E1Y8sDzpvSKrwzpZQEfitC13orPr7LUNgeigkZ5
XTLLqMTJt490EOn3XFCBONFkktmv25gHTSoWXWrNkOyvRazTEi+KcrtoTczPVEYDqyzIsL+NBW+Y
MV7dRkCy3HdrOtA5iVzx+kEH/DBS5R93o5l38+9i9xI1NVpblf8XVbaYIKFOrvfI+11sZH4NSEd+
WijyM9ErKTwHUFUeAUFRsiJO9Zke2/v6CD6hUCR5e2eZ/ctlESOpekwZe+hYzr4onC7PmLjIE+Dn
5yFIElqwFDHz7gRcrweMlfszAnmRqWlOuws/K+gohZ+m/ocWvRgoIS9gYtQrEKnec10pJVY0RNb8
Ik4sGWHFPRjNkjk5VW1Ans34DGEOPBkPoRca3kRjVnVm6yRVZTYicTQIrJKLj1CI+tdf/2HXWPtN
u/G1LfaSXGQDJYv0Gx7HlpO4QaZYe3CzhHthvcq+4LC1YD8zi+/PDDMfZ5Pj2GhXUStIHzaEIOR2
zHMn/VE+ODE5A92BIbQiKWx6SZ7Agwb24G5FQLHlgTcVPIsbWaTXmXbuDvcjWMoo/32Y6PoKhwIK
kCNwkfp8/X726BK83fq+x21QwezYPRX7XhjtCvEgsThwQCARioB6dqhLtzSQDKTpJanT8v6qwzK8
9/lSYYhj8veSgmyvW0bL9n+rrvHuTFjeKBB2xHDVlL3YyQIO9pFGh/3I/Ly8f1Y0NyZ223rCQHHL
YmR/CLvqVjoRCmF+p6Cc6aapesSBf0Gn1IV+0mk7Nwi1PdaZfwKaqpyBe6ugyY9uTRCTeEnrQiRZ
P6brPBfqcGhaIELlR/uYZ4oVyEUSovvHa27nVSfbHHee5FL5Wqk1odFfKmRuJGRSTLwOByXRr/nE
t2ZO1aV4ptwu2UIJdj8G5IVkNlR9/iJhabY4ZgzT2K6elp3JWSGrvIXldNcr+LPYF3lUGlXToPji
X0UGo5gHFyoZopcy0Th8FJW0qdSauUxUEOWsRbIvZWkdw7hzv3Mlp9rviHD19eCZnfQTykpSvoGz
nZkENVbdWWDBmUIHMwHuF/lt4TocCBm59YRCeqiViFNAfKIuHJzKOcm38N+YKk4MP0Ro78iZi7tG
WyDePj5tKkhCyYErwt95k3EpDvadHgkwY/LWvvAjkRqiIKPznYYeJuL1MH0vp+4uQr1SAyeTfVUX
2xQ0gtW5OYMpo0C+BrhKj4PjU7WxJ8WOgdzqhKuyp+8+KBO/7mdZop9rSnNrbSGlyNDCBZO6jd33
KUSmLf87rTygGvFNTaWI3mOa2azhHBy8WjvLSATLW66ShCUaM4Yc8XB2MNv3SvbdknDZuFXqfbsa
ChWuDOIMhytZR23n027ImnMeIWqV08VJ+bcPZsz23CGKDQHOwj4cy1S3PqiyyMcuoU9W05tgGkSk
BFRSqXf0malM8dz3u9Cu4kK0zPGN7vWVCIGbXFk31sxCrb0IlUB6onQj2ko/hWzhvco/HA9E2lA5
HJ7prLNeX5Q9vqHCXDnX6lbCPCed6yk/2mLaFIhGx8pC4gCWpIpBWGGwYxlltQT74jd8ytiwql24
J+/gKk0UXgkbxJMcw5Ql4yZaJgwSDwm+duH7dOFSfVCwDOdth27Z8reWyJzwa/UsHJYwHItt5NTp
2E4DSKc13GoI11zE5hDDubHqdVvgxhsGypwM7AbRR9PGNd4cGyBOQHzE3ruDKgTg95RrDph1G5Bg
DtgFDY4cpIDeLV+hlvJ1+/Cs4jHJEEbwffEthnkLSwa95QaCzfkqU3VmQckdN38/a/8y4gYIV04U
e/UuJJtJ+Bg7AqPRQ7UP/M28tEK9YfQegUwBREBrttIQ78F8EO9C8a+cX5hONFDyw4RGvuuCikNi
NbHkfrdlbyCbWWHLyOU20pqr+SMXluzZrf595ywf0pG5R8Gh8IsbqmAsWCd1zQV9Cv5l/wjm70rV
PHYMY4dbqik1uUsl7xq2RuyItJ8M5gT160esdT1yxjMMs4C9ONpInMyNXjRKu58bRx4YB40KDNcw
B63PcSUxTscIKm/QwkmE9/KcURzPWXyOJ2lYsahFwm+Gxr5VWMOq4ZG2Cp0KuwI/cYAnm8hYYTGA
FTW5+TiLNZ/TrBvTKZ1IEcMYS9gWmjdXj5NliIX7OkEX7HMBsiCV9F9fFazVXWwva2LmZbC0GSAd
/FmYhYkRIBXLlQk+e70+nMW/WteJsjm9Rza0kkmMllQW7ul+O0ysT5sKe8VUTR4XVZhGnF9+jpsF
raNCg3V8UILIz9ktz7Colq/OZDwiyADvT1T89Sm9Yqx9FmeMLd/uQStSlcxxCYW8jnTvLH7S+L0z
by6YVk/P1zqdQ4ihxEuGHoJiH8trSgWYmgG4VV3L850/OHlZXOCAw444tPI76NIPQHxA9Wz89uuh
9pOk+pqWab72JJ4hA1LSUrBEGeiZ6/x+KJPThJX6iM6ezDuxAsZVOk+RI1B4852YW60hmo346y1v
hDVjz7H+GW9ivsPiO/0b41z50qRG3zGGNhp3gt4rOveWlrJlRlHt2DdCG7AUNaM1MZxRFTM1IUOd
/cS4BuJjZuFqRXWvh0ERMwxhV48g6s+GyRcRP+lmUg19kMR8X4SnzUIPn+iHh4FdrjmDPFIosim0
kW44s/w6A+qyTBSbYYwbF1VLoXdKD4xIC6Myp0lT7/Y1ix639bLu5DNKtwnL1CZMzEK5E4xUJCVo
KM0260hFw1JWHaMyvTzzIJWyK4deGRSMVO+UyZ699bPedNmtQ91OYYCsuvo2cni7/+e040oeQuEy
LTWJzRuWMD1uFbycQOaY8pai4t+fp0oUe9d8RhMS4ogp1gPleWk+IYyrp/aQ9qExNN+OCZ0AVsQ5
RDCYxrdildlN+0N2yFJEhxo+xm4Nryj12OaeBnkaw6sW2q1ffE9hVwC8Dbx35yWBmGGtH3bjwGiE
0NZwMN+Z++Z0q6QtEHxp4YLGHNGlkqcaVhiYiBRlG0qRtr2Uxg7NTSZOLYtlYkQq1bvwGKFzuTmX
ktqk5M8hc+uIq0m/wyA8mVqlxQJymbuMPcIRtphgG/drmOEljsyHF1G+H0juffMZ+G0m/Li8uIKG
wDcnnLdMGmo1wT3AYcOKd9pjp/TrzSJu90mQ+lanHxGuIdlZ7XV4/Ofea8DVeSDmE731QeuIt/nG
OvBgWpMUiA4m1K/q3lpNhsNJ29JCp+J4GY1RVAgfGXBwp4Bs0M1E0hXFD2gTkkVvTQRJ22TMtJMm
qJPv1eUUjIlMy2kfqHmRmtKrjt44bTJToaizH9e8JZ1M5gA7xjqdvD5docLuDIYMH9MITM6uq9vI
8xcfdlilLqBwXue73xlAcT8/5nbAHMaf/063YSrGOOYm6yMx3zhCw12wP9UeqdsqfEB9HYjJ1ln4
DNc0CXr6PhCyUY2mIqjpoN0LG/DOsKwk60t1piynMsl2KmMTtfk7OTT3GbqNbpzxsfpdk57dWpMU
NfOeAiu0jvM+taJm0fU7F1dFRd8pEVUOSfzgxp5UIrMs6j1jB8dw8Kx4yH3wofqTC2zjigrFdH5/
EUX24mT2hceT1fbI2OPr5J4GVUJEKMVhMIT92Ku4pOKAqfvLT5FUEERsmOkkMF2EU61cpOwrs4i0
0CqkvxGaDot5V4wQh1XfNC1eKrCTisVgq/GfGGzx+ZOTHYbIhsmIOL7JziAch+1O4AXGoK1Ui6k1
tsWfCSzSFtY8R9ZHLoxewO8sNDsr/HnR9kFOEnZg/dCqNMxzAvVq/fcdPUpK7CkYvy2SHG5op8C3
m1nbYv/UCDduoyi/4JAuzBrdAEZNp6TuF1ttuDnfYTgsZijsy28Ctd/dClwR/TWyvrrTtToabhsj
q0pS2+43ZJzEP7SDMeNc1j+2vxeIQ0JGi5L3qUse2WtpFHWxNXDNmYNvXNvV6Uol4c0FiofALkC9
GIt1TGT69cI5geTYS72X2ayzVPolMah+6T8uDdVps/cNN0ZQWJEmUOhn5+Tf224+W8tlIN0bHLEr
QsAI2uI3IbckQZ0A4VQbB41EiiGZdoimyhxUvCerB1iiXgVlO4JLR1ID0B43xptEfFOC3cTC5U+j
wNMwrtG2r0FjL36vS/rdKI7paL7n31hCRqXhxecpGFlRNGX6PByGAmS6UF1g4i/rUhslkgjEtmrv
c9lZ4Sw8mMuCu01ksvM5LyqaPtJjeiSQSj5aZMuWEBcydy1LC3eoLTpgO6gIrEHQW2U6MRo5SvKm
3nq7VYXNty/Eh9EoUuf57lF0szopaAFEbNUxnepG7iNjXqnU+RZaY3Opjv0g0d+u21YJ0+gvr94d
xiWAmUzgZub0Uj6GsVcSVLVFprwfACd5+sSmAPoYekkrU3feUOX/f/wL7HMpXFbegYABCFyvpcou
97nrVAdMeZ5xh4i/VrNKQatvE5KGw8vLQx0Ah3tYdDm7WAMPYCQXtF3yDpxALr80mLIZtkjb57He
LqVxYMQp1BT1M9g74EL/6wgMG0fxXWQ7VWolGzkrGCgpULTDkJhdG3Z1ZEmUkfIS92lgN7OSQXnY
w3kcddBIVLmpNeeQciYTThfgUff/+eumRCWwrt33MJO/qu3TQHcmKpTzFzcrA7Gx8DWKZHr8B1cb
vmE+Y+2EKEztPYTdAHLWjU2hgH/5so+SPlsthbRrR4ZnH9O3hOTPZ7KznzzOPspIGM+Nb1SKjP5z
ngzJNnzCMeUP9jf1HpKAphggxndMA90jXVQEE3qfkrbMR8kBiPfsa6/onfozU7mEja8qwNMyYtvI
BXmybFG2UQltCpJVpmSahAtGH4IPCNCZupwlBJ640pt2xf0/uWSfEnMD2DX3dXYTrHXT43gDVx3S
/bvy2HOH5OOZHTjezXbNb3dw3ryODbCS6ix8VjEJEN3KjyG1cWG7J+2B8zlwjE5hw4Dmweb6co6I
Q4BicokK2jv/ebnDAus67b+RDQANM8+QqmI1lZ/4/4iAIGhSsuj421tUqeJpl2bWwmyQP9BOXxh9
LBaDEwDFdfk/CbDZT8sS7CM/N4ksVyXVcvrcoXf28mNPaL1otGyXgTdygWhHSZyDtGMuJkhvgGQH
wa5I4t8/BjYor8a94MBgt2bCpwCLIXUz3uj5CnHBa3YW+2qfwf/LskE03UyqIUGdIROoZrluPTWn
nfCPIMbMmldy4CSaOJNavxpzYUdU+sRNd5ogCW9TMaf8CJnTMFtRkFzJ0ZfeU6gFcqkXf23/aFyp
w0iq5flfyTzZsg5xvMHilua5td1j7aazOS2S47BVxMSR6g2DQiEaDj2P02Ph6t9nWj9KYJqv8ydd
Ra06YpH1E7yB2Mkeqs5zx/lOJO0ZAccsEG8JHQG4ourmNuxnYZXy6SiZu1lbJANcA+whosOnEhPB
oKzCiQ5paX8ws4NhKNMwc9PD1Z8Zrvj6obYolPGKbOuw2PUy3pSOonzYsTIWWeiGjmNfUCkIDzLj
K7U/UbwWV4K4lMlsSrB8udtaoztYhSECRloQs9Rf1M7q6SP0ybjb0a7yEXPNRBI6An+qgUSzFql2
iX713BCXqH7t9IxJb52by73mZVYoRA+mrN5NvSsRfJWo206mzWu8ErLj1Oy8ypRmmT0jr+WHkPLc
U+4Y87Qui2ClrkkE324GRonwZEBypiIa+EpmkwR3hf3ohCJXVjNV6YWLySQMpg8ThWXKOwxPt6mt
1IRmBI/0DUOCmvWwnKYfmfU+xrYjpCQNL4YQFNK1xgagWJOd1z/58f3oqlCyD1/8dEM5hyMhRMzU
rD+ZVx8vXj1g9tl8zrUeOkiAHX1PnJWhPmq4Rmwhcn0UB3XViVNQ0V5mV/q/ZnIc4EKrX3nIaDMU
6TnJRVIn/xumT/drNparjkSGYefwaN9jKkq4sG3YUudOJ+zYEPbQoVhp1ONOqKCJwc/poSUN2vJZ
XPdmLCnwl9sFNFv06n0LNYH9JAQNRLWU4D7yaRaPpKFdh/4XDTj+rHP6c6MsElc6SWYo+2h+ezG/
8GHqysqHlhMKX238E1UCrCT4S1KCTOE6t+MkLxvem8umJub5TVC2xb5CRrcBTEuSM9rH+jk4qD+O
9+CJcq+hOx/SXIM98mU25JsZt+Qeu+uFI8txzA3A3O+rceqh4K3GwF0FttGxHo8myf+Fhfh1s2kf
hxj09e7O4DWLlBuVcP6Np4t6x37HoHTK4ThakziNl1t0qoPikQJXaODzW6/JxlOPtFT8cNyolp5E
cyoWq4MKJUBTUmpDcXGpSemsp0umQF80FIcvMQ5n/G53vjKhgUQelZ7M/fLf1AKq47fi8tCnxguf
hSRSn9Iac5BbI0pCqVeT53Hz3gZqldbjJoZ9gCQzV5Yu0FGyGJb17VLZrCvxxC//6Ffsogj2XExN
eYZS13EA1Nz0xzlvmEU8kTQyeLTdcVlOlqXWj53bq7KoctgqiPOSIhItCv19Yh27M5USLa8KkwOv
TR6tJitJvSUZ3arv4Lo5TIXaY2sPkZ5lovLE8a9hU3fR4Jy82gh6Hatht/5DGXPSznkzJU0EX7Ij
On7BaFI+8fjJyDRcfxPswolRXD6yAMh8l4dUkrouDYtGPAzSncqqnyRMhrGKA0AdDcDagn69josu
lvPAom0q+f93jEZehLLQyd3+PZmLL+nGYIdGUiyy8K9hutIZ+j4aCh1pnqVc7IS1rev5TfYA/s1a
izcmShIuIBC/CUnkZCJ8Ydz7L0ca3f0e1dbvh+hAjjVEzd1zwJK3CSOA5mqnRFbGrxrDTi/h83+T
J4erwYbUPNQunhxpKuc1JnyzdVmBkz852ZvE5xzh54sdqSTcV+B53MviRsOPO1g24d/jv2MW7tb5
GT19JqgLy41dZ1XmwsdZ3ZHlNvxVddBbHqprnanKM66rjmb+urhIRxr+SJXI5bzzwYFm7/AkqFD8
IPuHQw+JRTaaRdFHfAuLOJkyaGK3d3jjkTGGkUxMLXSGcB2raTBqCa72GFbE11Bd5e+co+yLIbut
N4+mnE7RhwAQ1sh+k1/kLInyde9To069KIMpGHKU4NoBJZJrwZDhYzCj2C1ixUyTCz8Kik3SwT71
jiIEl93EIPj/FC9zfCFY5C2JrFzfEI1a/rwz2iEBfQFMoSU7FbOuxoZU9BzfeAtmyV2AbRP0DFqq
26W53wHu+57konXHTgrPLeTbsCZvEbkrgHzQNd2yocDSoSVBq58yLLWi5VP0/26bdtshQEnsIop8
UNPfmTNvSU0YcBkTsoBxQ7Xt/TTeJ/SetK7g8BUcxMG2/J5F6csW5BcY+0Rv8ydh1vOZAZF8dryg
GYTVdPwND7eEWDzZt8OtWe0MWy0DqngAqIjOJdRWnFxeiyWdWowY/Jjqzj88uJ+wfQ2JNbn2MYO1
zrZ/ceVj2syVf3unIL4bQcpOPFEIyfblbMjnJ+m6LRuu4h/A29IarZDnOQ+UH/+ZR+oHFR+tSiNj
Sx9WmVzQr1/T/VPEUCK1+NhB8uR/TOunsg9fiZbpN5LhOXsblRdNKaYnpkoPRXUyGoDmXaFtMKFh
i6hvYiW8xd/HFdy4GBlMXH+9mEc8jru7LTmMkmeZ4wMewTqMqipQWuqAHPRDX2/YNTuHMYsIfbbC
0jGd2ND+9eKCqj/deTi4ZKUh28LbO7/dlF7FIly1ovK+kY0B6SEpib4OSDB4LVGKYGRybbgNhhb0
ygYyTi5/GSu7bDcZ/V1/lfkZnD2SpihUogAZvhZnQzAEcu/zcFJZsSJnFAPMImCkIBh6GI702Rxa
O9n/R+Xl0H+4HyZ5BwV1TzAnK8wGWCTOB3f7IzQdHd0ukuKJ3d+uDbSmfkBKQaJjT1U+B0FOMi3p
/Q3Q92KvDiAHMX1CzvEY3hU+FiNQnbjUT7aojwDXBBJIejWoTKfbKcLbOAtMv2yG3ca8tdopYnEI
HmgJ73QwWAWVxQH4vDfAsP4sGA8E5wlBSfF8p7JiIq/a9wq5l3r65YmR3xmZ7JSODa0N66qq8frP
Gkgxlh8tZnqFxH4Et6c+f4RPxFFqDLJS6HTJAEvfmPZHOxAsmkJJxj/rbuCgnzy4yNb/HcgFhqg6
skFSnb13BB8yW8iAfbTc3BlzkDuHuTjWxctDA4MTrUyOtootCRx0ZFSwZkJyosXSNGxzU4yw+3Ut
efh/UBIybzBDaTBH+rUlMZwjiGrQ+lb2771N7pj/4DAwUUcPCFa3WVPvEXb2R94Iq7d1aDj7qWyt
iLWOMCAaK9c6HlNBKLV+Eplx3uy++UvjJTT1jIk9ZDfdAh3Zx+Fntgd+OUbKzk7xF9d2qyoVo3qt
0ptLIpYDJ2OLdngVQ0o8XKF37cnQKQRSrA1HFBNhMWDO4xrZy5a77PB766YMvIkVfvSXjMFpxZby
STBOKRU3YD2DcDTFQ3kI6U/XRBinn503zHGnVnujIVmjeiubFfwOPbVLbhnuI7Lc1AKEcH31cMpY
vPVFeoyx2YD+PEVLcuSsLb2QoHGp1UShAk6KRhkEUxJWzts8gsHug/iyRufoCEyhSPHMuudO3+UY
IuAN/evHILsl5o5NrpF4dI+ECSFzrr+37+PIGGIqzkJT1nR7TcH7wC5l1DGApcbtUvzOT8/T4Cn6
YHfBnVWzrfOU0HLYrw93NXGAtGJNCQxHMnURQaKelMEiGl4jrq3MsSrHwbiuqKUkKDFuLkgsyPq8
iFTRDQDmO4uGqGMSv4Njg9/bUm1ICXYF4z7BoMg/V2u45NmaPVcvUpaeicO+GMRhnyQayo9WxE5V
G+0RgSSTSjcF/WmAEUVhCGXjB8CtPBpoM3/wgL2eZcxsCpTVgZjP74VbldlUjrl7n+YyCkpfcXx2
brfo2RWBTsSuVw+w3Gp9dIZo0ZRhFvJD5tYFU2MB2kWlfvNF92PhKMSz1svZUaGRwA5YRzM7pE4k
V/oUXsRIHpkP0weHabRx+UzrwJpoVsGlGs5kGxMhQvEUag6lUlGNgrosiEWIK6NFpuwft7ODF0Cs
wDW+uVg6082tQKHiaStkf7XPaFfDelNHCoPIqUDimKV+3G7q1y+dzes15sfdWmd/8rwOvc+QHLBv
BCzIC+PFSoHeGeXvuztEONywcxSmo6nsceHgMgEh6N/KEdzGMfh251fiBKxV1DDPODgQPBcTgA+w
V21amz2HGeHX8WJVabelAvFQatLxx/LHZxKB3J1rWgH2+dnukA8nhbnLDPseu0bUZEvA1aR3sOSR
7mUWuFBxO5co2ks3giTCjF5kyGtkWHInD3Ykup671IAd6KTpjzc9oiWbS5W6OjqdwbUoOdJ6kbZk
go9EXLAmVeM+FOv1Vv7KYpaDbVVov+d0taS+jYGtPH3EXopnwX7/fZxBvJZAOV/N1vLO3cwayWIx
O79ZEYlWLw0qFq7zXa2eguULJBJx30Uk/w62JAA/Z1XNkrCJczZYrqHzpHSQncyIkjC6fkDXek89
0Gi7Aj5fCiB59i7uFKZde+3Lj3ckXUlVv/e2m3D2Yu0ALLlg9mx0RM+RqB1801pv+EFPkQG55jL8
lNa/dN4oWRDkgcYOfGPXfnsbYKwKMsEevWTcKIzGK/zp0XREFEPZYSVQ1bJO135zSKJXTT7y8M8N
+io+wv1zlGyu9+Dbm7PHsz+bEkozB2usM1rP057AISKD+oJtyAfxYvNOQUgCrv21XwyAwNZIqcSi
loiLgj/qqdmjOaMnwzhiwKZVtIblZ2nsb02hxzjzJOabEQifjhi4149DGKvRr7uTmGD+ck4j7vQZ
yWeDzmCEjRH6gSAl7mc07njSzs54zKwGChxFMw9cNyxFx1wqYAP+GWUptuHOL5Z1VrcECryrssGG
CWIBKvLifB85lOZEjtjQDrll6YBmOSrzTcBbAQ40vCgAD+8j+aP/eER9rjWp0CmPywusKGdug3vI
hB9wqzCw2x4IH3JUqOuoNQ//RZEfkRbeV3C0GzqZZvw5BAa7uXt3ovwnDlU5c9BRmYk4smlHrr6T
L7Vc1JOe49jWxuo8qNhAKXRjh/86TkKlpnz9txvoN6G3UH7SCuHWlz3rRi1iJrAIJHFXqTzbTWrn
323H3kDRiMDFsFv7O1Eozf01rf/dIAZNc0wk6uAUtFA6NvK+8Ia6t7YMIMJQ3OFaacSbGP0g7T65
rVXEBG4vNIcE3TAU97xgZ7EiXVLtqeUVXGPUF02WHpI9su2e6i6uuukiCYDEb165MGXuga24KEQ+
7T5PJasF3I7rgZtZB3OmH08Bknp72zN5b8KIkcIKkKljRG5cV9mySoNcch3uqPWJBrnkFzFU83Cv
zJ1ra45e1cs+lTKTNiaLwi+gyY5eFKm8B2rbQqr4P7cjT0b0MV62nF4q543JI7IYVKhkaVKFb3UN
j5IeDjxZHJIG0gZP4ZkvlM+nzzd9AqLLtbj5AcRg52BeX9x/9hUrSY+erVeTnKZOTwnUrINniZJC
hc7WOcdpfNqTMd3g4+pITyTNvs1eXz9FzsOuhzQ2ymEOTRYcJ5zxUY9vAEqRpCLgt+Ci8fLj1By2
TzASmTqRqPAaxwJ9+FATO99EGJh/jZHuOb35nnYilSVfjqVIEU4ZNd+CdMf3y9ABvu2KvulbWZh7
bFSys/3pRqMJYo+FxPvnAhz9mHVCPx62n7IOZGLEfZdP1HoHj4ITUyHjyx082g7mnZbtlOWp3M/4
QuwyIuirNRcYKAJlJRl7QPrbAKJ7w6qxfB+lS0GYdIFRCfRSFpxLsuCgJvdJNh0D3qAQZybK1sVZ
kwdSTSVlcTuVtmgDcsHehLuShtAEm07Mlxx81Iao/Hl16/YUhPdXAN9xqIcbMWFd0d1die40rtuA
4lMV5+N784rbzwHKVuEkAuAuiLa1SZyVSZHbKyXnnUsrX82AzOW4uUp8zAP/yYMx7/Mg0+pbiLlE
rDbJ0VQTw2hvedrwx0biofVoshb2cElzPYct+uEwWA4xKuWSBEEA663+v6k5EXZ9GIVfFt8l1qr+
kqwlcwR72IL4/zuCx6XG8dp0qdhOMWBEmxPaKfbXJqGdlfs1nwhPPVEkmLoGooqzNrl1+/iXVgZN
ax08PPlOyvXDNSYxlNx9CTOI9kRjEKKv5pBhmbWpbW3sM3yylZvCU+cX731LMHyoiP9qXL2lHNVs
hJFdr3AADAy+JG6zfKl7uBfeAQbGdOtegmbE0KAeqefjHvOiOKybVFz1OWpn730psgRmWq0S/b4E
kZPMeP+dXEQrysDVbTxMz5Q3EGClUGXoQ7tFOQjzdjq3cVj6hk8jiveL67WLzXI6ddw3HfGAS5QY
4tBqQJHkZOkiy0M8R91phVJ+J07TZkP3rdCETxMkLV5IMwkmXVWxPr0EpwU3DdDddiUAzYfbuBKt
hBarVrS18kDt4hASwZWP18laVvEp1y02ES2mCLTrEDSpYjhgWqMxjtoO2e6IoxWkWZwJpIla1R7X
a2awTpGrXn/OYVYu6H2Aan1NUAVW0kXvVc8RH9tZXOq+o2K1xVI6Ed88MhRWgNDnzZV0lJ4VZIkE
lYGuBRAzyVnBGoACGOYE7E9VkrL0lKgFAyS2OY9BH97367fKmvjlGnlLRij8814/IZ0DcaJZxk4O
z8NUshWaiJyQSgA1YPs/Ry+jATAJrimgJE6qIuCXyYbgD74GMKyO645aRexumdoz6SKr+hSRw/Ue
rf8cGD/bU0h9hzE76GeAfWJQaYO2p64kHN4nDVtB2XPMkS2NHaS+7+3hJX6iPedQi97y5m4+wSO1
5cPlNGyPj85yGEPu6H4j8VWWxxdOgsq04t6Z0LUhpQp27/Xtiut/vZrXS4k0MOpz/XCoZRVxs9LL
9pATQ1c1gyNXNkeDl8PbTOS6NZRdbz/QwWF/umXj06SuTLAyTI+4CjfqreXtA63tTQBTU6O/DKcA
hj5K4KqEUwKVuNmIDDmLlZISzVFcPNpNzA9HuuP3SwmNxn6bd2KK/Q8rm6yjJov4Ynd6A6XCD/CL
5dm+6t81H2uZCMlA8vmhIzt3jVKsUxq/YX+e+jafoDEys+ukPokY60qlSZPcxdm0Q3XWKIe0rDlY
dydWgthf5TnNf/9OtkUzMptRuHs1XkwiIMHw9VDvNL1RoEd+iKcz0jiiyD6ql4TAAhoNPYNAiDI6
MHy2FU0m7/+/TY554UpOF3UJhfgHjfqiwMhzZEgSiJwOhZklIhtR0bK24xRf7OlygrzTqJvQY3ST
sIyHTp1Kfd9OmBMuPm1WM/JtWQvMz6y4fdxQGtEcRMOgafCMNZhLUdRYMZEcFZnhClm4zskzPwzB
bi1pmBHv0+xkwortbzy79JgFbfzuTKQa1L/o1iVoCdaI85Uo4gAIJokm+FhqvAYQi3Hk5e/0Cd+A
YDNKOGtFwzwhu9vzSh4LmtL9X1GKo/H2M7+JEdIvMAANBl8LgxVHyJm86oB2qfDQbB4SzDfQefAF
y6BsTr6paZPljtUigBdgufEEl+NrMSFh8vDiAX6vHgwqPkIPRkKSdCZfOrkMcDVG/D4d7g33Moee
oWWNPR77TOb3Sldf5vuhu1JYIcFjYtBNosgMBVSDa1ZvhZzU/Wd4jqPp4rh18cOIHCxRslDNuUzB
ph8NAWqVhwW9Kt72s6RY4FNa2/zq8XC0RmxhcLSk/LDX4VHiKHojy/kOPVURgRsKtKe1k06VahF0
nwPPmGbFbQOc0/KDHDefBB9p5/krWcoY/6N7HxXchnuo+Rsg0GbImewP/4KyrFAJvq2PSApaIsB8
09VzOmoEgQN9263euKs2xmhvs0P1cLzw3utcSJC5JMqQ3Y9NBrNCPPmeqdtzAIEMXeX9bbBrQ4uK
A3CKD+Vs/+Wg/GpsLqkzguZSGh8YSBm7MPJuBhy1StiHziFB6vZmH1SoP0mUwxTMFfyJcxD7AZwL
0JlzDhwd101OOeANVqvSSqz3rwRXKIaIBzrl8iyufX5aGhKhhAaFbKFvT2MgmyacdpvMJZi2ip+Q
73R+QGhOymsbSZCITl1+T4vpKT8p4JIt6Gai5iCI+J2YJerKNJ1z7nfWRJGpbR/hQSTUTrdBIXlo
oFVMpZ0tHk9RM+IUl+Wx3oeieGGhjLogCz3ziALzHEX3zJsiFbNQd5kF86o+Dq5ULyuoSE7wikG+
khAkQ0R3Pp/WBR1BggAXm7OiKe2AYQZH4++iUsFYAHNCBrp+nG+ipxQLYDf5wSCEm3TjnPxjcn+0
uIlvIkMAk9/k+TZ+z+A1KE4phiGpsPbyuQS9PeDKE/EItz79HRqIzAzOp0auvZQ4g3ndPnvWL7RD
NvY6ncLx3zLEAzd+Dvfls/brSJmTwuoELzHQ3yP5QuteeFx6IpkbYc94XLyMr2M8IbQA3q7A9Omf
H8ZCf0BWNwEmLJS65/0ZS/aZkojpOFYiSah+pSrilFXDppfOX4AoC+WCjOA+CsH7CeapRqq79HIY
zocYE3ShX3CrERzRssR0NW5UUZCsFkCbnjsnmkC/wvBS1SyEUKKJBmnzjuTwpBTExadmrk1Rx5kI
w7Q+eikn8mcF3t25fBFb8jmJpfxxQUDB1Le7y4c3x+Pa02k8h70uAtwHjNNYa/VElUObEQFmbtVt
Qd3FOp5DL8EWtAPeSc5+zp0QTz2VzMI1kAJ6kTClvwnWTkrkz0TvtkEfGM38BwFEILrxt5YVNfKf
wD0oJQ4SSZsKhESHifhQ1n3/14bx/Dy6qsedLLEtIYD+U2v/T5EGVUCWAdOkQ3pkOBSb+x3GXH9m
xS4yF5qSv/2jYS4wt9BOJz6MBf/R04sKEC23Z71fgfsIoGQZ/ebaCyyd3zgfpIO0oKRfoIqhYcBJ
5pK6I36un5xvccg8F4dEX1iVqb2cpCXJwoxiYyiYWHLKZHpQPzUmv1qBZQUuWL2XEgkpfy+jfHu0
08Tp4DQBQGPRgSq+aPtG7bLn3/VYRCh3urMofbF0bSb3F5+nV0oF6MXvMavPS5tRpmY9RWAfoR6E
qzYXPnT5Ezvihca0bcQP7o7NulyJ8giimZK/9K/9UB39X0mAo8kj5oUGttjaEhTYUBi0KndeqtRK
XstU+F2KTaTnFChe2AA5ScPXQU8z6dkv7rvOuuGxozWDr/qsKjrdp/1FYz10Mn7K2Zh5gBzRq1zv
XkKMT5TXf8DN7iqM1Hg5ZkwcUF2I30pHlAFj6bN83lPH83hsrKCI+yoPn1e2+TE4Syz43vNM9CkB
Nis2WIGxHmSicJL8pIet1lBBk6v8Dl9DSGnqb4hZUYiTY2RbtTDWSTOpI3lBWVroR2rSPmnzMp+O
GUiFHDyJ4Tmzk5Yt30cBgI1ja08p5C4jo0HnfAhsEMJR1ieSVRY92LLCvh7qld99d6i5CeFjzKFD
UifLrTKtlPyw1EghGI/6AT55BFGK6ic5sJJFGWoLasZ1DqtL7NJRzv/hvneHv+rJf3gUtFJtyKdh
mLZhFJqGgQvHF8CpUw6TPwQ5FGTGU5JyS025NZ/o9T9z8q6cSIuqzKgds0W/f7fFKHUIQUKn2w97
kSZlyWKCR6BHG3+Ulr1gj02/8McYJnN5P4Yod5yDZJYoW0KP5STsW0qkItpsg5H4Chl6SXxC9ana
asyb9QGJo16TYr5ZUQdSKdB7ynHOkyr9N7hoD94h2InKkS44htG4YnI6g8pNWLRznbpRP3Pxt4lA
KrQpttcSPLyW3i6KYVrpEwotgePN9u47wxnwb28Ja/RAk7Ccn4Kp3xvDtkGIujVRdu8+W772eDrQ
smAiV9+dgOUn04XElonaTIZEQ0Jm7/e4P/0rOA4kmKkAnn3m938SsaiZplnOKbjjXqhqm2bvaCwx
xB/PO7XU/0D9IigYzlIhBUi/j3e9cur8j5nSHxWSMHc6YLIWQySKKMrjHJ66kHWv17fDoibtflpn
y25DDEbVhULL/3jbUUzwncgoOOzIgqfHj1bK5cxBJD4er589Rdw06Pncmpfq83LOaWzRKoUqVY3I
1tspM9/ihK4yQpixteJvcqlb1GRrE8NGBKx9tHkouDZXUOGDc6Rtu1FeECdPFjHqJQDO6Q91sDFv
7He/be3pb/Kv0D2eEmJGotFrZQqNt60ECEVvJ9rmFTkzE3QpToXVsz+iMi49TVVohIHrVtE09Yx/
EWF/VaHvROaPHjh5s5baRSkW6vpFohcevI7vyQdmlJHDrABIG62qyjhDhI48VK4Kb2zHckm8Oqop
OYFo0BkeN3y399Ayukgqiys0VCIW2InQvLsQ9Pb7byBYSvDsOWX+kQNg3RhPArDZAkhJiAh+/vS0
H8OWeIkW19Sdl/DHNJO3yW0R+UanThbZUheUshnNv+yZdGRS5MQO/TrXpq3jQ09hMJ4GTeBjyQwU
zE2+M8GHEg42DBQ5HbWKJ6TYAVP87BsLNuE9aJk1CQe1BGPbTByYUmpT9VxZrkQMe8pqcmP4KfjM
HWt6IyPs8MTKNbjej7TC7nbx4bvOtETuPCEFu+M9cvyxas90VUZud7t4pl+3KGV+Mlx1EOlTm5ie
X/2TzPVuvOlrXPcSs/YDzCVRJHf78Wv+YhSnPLHnN3UrDOSwsW4kfHVbNiOIE8y2whIn5LIniJ1b
kkgvVc+OHfUC0yIE9eJcpBdOUoE9aIXKy8X9ufi3hTIEjpru98LPL1Tk4QDJMrr6f/t7Ep+gPKJ1
L9NqONr/Uzu4mSeoOYbqDfjhblbdQy0D2IPX0IvLGcmGoiMPB8thPhfaA56TuYJxKzI44w5Ve8rT
Dz60GQlWHKsbIN7uh7zW2a7WencvNt35eitBY35dnQAdp67pdLbGJwS2KzGrRsDO/hC4UMNONHdH
7SJkkySvPlLQUbilUkSue01N41UPLIDn0yW4BI31VtRQInXfttCLezbSmxD35Rl5hqGaDqBYj1VD
n9fQMgK/DMN4Go8loTxldknHff4H58sInDM3Pki9rar9UdO1fdEkZ+rHi4H5XmWGjMxvQq+E0W7T
9AhiM1dIGllkAm4fFPajsK+yUD56+W+6RAAhS7An/1FQED4/rFnrgGZ1Nygl2wf2w8pl6EARd59w
//5FxWO7L1mA9dYbWhtZJx/poWaGfyrXuyYcGOcewmZA4gdcXWLgmL2NeJs6gliLtANJ4rV3ZTON
VF/nvdwH8Q6s1FpfoyjDEFNx5a9bwnJiz4Sc7c9oLOS7YMiE5SVzddUgFI6M2G9WmYZYlp39sk3l
RIl4B267i3GCu34jsfV9AkfKzYp7GcwCyYVXR1Pz1grYS9PeBulZ8IhD/vpfioroAoeN+n58vRtu
pcVZrTia4lJlG2z1co8Nbl/mwyniVOtb0Xbhsa1FAkf1u86ZfpSoJxl0kU9voG8jgaLAwHKndnlw
mIeRE+xzSX9EzvCVHzmfawYrH6+xsf4QZi3JGx3w6xo+Oev4aY191I4Wo/2jHG2vYjX1cq5X0+G9
pwHeyiaBEzn2Plgv/XJ0nhhz0tAGKMFPrKBtmb3QFIBKMV3t3YyUCrZK78KviWvTYRdhyRRxHVW9
iqU+wYxA6zURNTXTGAodFp5gVU3aL0mBRqxslo+3ZyXL123+9RvMrqoRJNu+/zbdnniYW63kRtct
H1oBw0sHlSVavSSzoaoAwvYDZG7DBHKYPVcpSHlzOy2FUNRl9wYEb34Yhrwi8cCLXSjArf7aZPMC
fUu0vT5qtG2uDuuJizO+raJn4mwsKIhc6lOnaXZSlvmzqZ5lxEliR+jRLQDHYRQBtdMK88X21Zye
S43RXa3nEKZzezto4WtzvkJOaT4Tel/GWmlTWyZoSBBCSGjv7DKzjknRnRsFFQkLIpim7bLoQJpa
4MGsYjj+EYSd2aa7SZpCGXTs2I6AmJtVKi+38ikTviQtKuzGsciwgOqO/BDOH/TcH6rGCQA55XgS
txTV5e61aOI+f2iYT8562q/R4NQG+9c9KuDNRvrAgWwwBmOoDsaEUaKUDUFFaSZE9VPzvszWVVi/
/DeOAQ7cc4nFn/xyl++5rmI6kwvX4t0rqMtzqOwdJhn8QFUSVmyHMQvGZEK8EzolaLVySME2HTKq
71ycbzj0YK+etCH5nkUCxUiNGKiRJrso7H7R4R1HuAdBvx/MGgST2zL2GUNa54FBB/bK2LACbzZj
yXyLk9DF+Qh+YmAO1C+rqjQ3ZsDp6U8j1KiVIBLUfj67hGobVjCWef6uA8gly30LDWVOaHCF5xP5
0PSW1PYrWYivPbxsD4zxiFmJ5bEYrhEj0q+GqruzCuJ7ebSgS2h0vKzaCDa26wga6rSbMH7BM5l2
II1ldQNGSRNMxPI/jmmQA3nF0RfHAza+v/hiH/leAPJKJiV4e3BfgHlU9+5WivkForxHU6t38dUc
f3iqxHIu4nfYpSFSoHLBQm5R5vUUPJKHbPsDbgxOERPnigk18Sk+g6JHKSIx2ELWB3FRjSZC817a
53rTQtWeOgpqw7BBU3YwGyP/99VvfXkvEsSte/qelKxs9PrqKu7rAPnQuIR5Ze3amfynYMBDoNOk
xF21nOIj62IkZGEipD6pweJW3RSb7JSeS3FG0zjEbcow4VR1xciGlaf1Hhrro/EkbF28OHbTgNse
fz5CpS8S3Zslw7xelvTrJWteoMpDA/vi5TAGDHCD2lBspZpZ7cRvwQxXxlqzn0/E9rsi5XBoTgMz
CNwEpXVhb3nBckFeIXwMjiNjAoek9fYf2VA7wzFbNL4PCYOT4v9oeB/mzfCxcfZMrvI4Z07pfJ0z
fOQgXNUNNaGM+oOQHrtzUObO7TvFrb1ofGgkhBtnOO/A1bCYH0BKeRqRUfVjDFlYQ6VS1ZIcW0tJ
jPIbREtQyfsorPCXir/64QZfut+2NqYImJgK2+3kn716e4EezzXxemDDQUrc7A/D56fZH0PcDziP
7uqVzFCI72BG0EmG7fZgcilFonPR9uX+3h5ZBb9n8B+zLDy34PGVF6BQt25vKfI5NBpvl0NohI7l
su+Bet5FB6O20j4LBdNfFy1uSjz+DZ65nbyDuJYhUxRNDo0yUR2mQ/kTWDsaBISbKo0vgOA+UJ/q
P14fWidwYreKvrY2OJcSWTWhQfZLTwJ5vCfL6b3RHmbD3nxpEmnCLVX2JLQs5cIf6lZfyUkD9MCs
bFKtYNXvVdedgd0mrsC87+U5kT1BZ4uQ5iVyhOjX5RHkp7Z234WQ2Qvq7/Cqa9vqGdsM2s4Dr1sk
b6bTifpRGD0iwbke+cl5YTP6Y4BNuTpJvTvCVkJVVjlrLFHnKEsKrDoZlCa+hvxH68junUumwk9R
3hZB8SfiEIjK8K8yvHxmVtOBrntD0XpiAKPd7g1bKYDaQrtjZvYKHiSmBjqqi1oWeJ11xNE5qE/w
jW9AK/i8RCSslYH9NPVSoZwCZm9AVFV6+It3iYy/xCKTHolvLz5Sp1p4VU+6RMh5MomErI/8+HQr
VgFoTiG6oJtQDgiaPBTpIx+shNu8xE/lD73pNeRwsvz03J2y6su+PTM7zfkiEZjSUYjZWSwEmzGg
Ck2j7A5Kr7LhoH/b6TqAPpyNgiYYX3XV+/+XqQ7pQhwCdA3fWF6l0UuNXkYUFpatDVoSeL6qHEPy
+1J98mP/yWxuRD73GFgbEXFcM1rNikeR7ZoKP+dw/rzhzdK1t6GXr/9bNYkZ5M6dM6oKqd5J26L5
PRlQyZN5fQCldRD1T8xRye3/vMGR8DwiyN9mWsILt0qLfKIO1TYa0occYFETwHLXDBRZw1w6h1P0
WWrf49CR51+fhddQECBPA4SshpbYV/rN3fOM0IhtHcAFmN6LUidHoWc+lxZXyexmkWSuRW4tpQud
72QawKXpwW1n+oaVLr+ezWBWoABhp50ahII+qPUFK6doJFZkGFtTfNk7w/wcGpikYoSYeITtQOBN
ym/QgGH59WSVSgdfbyPf3cYNhyK+f/JUsbJ2h3dnkvGW145uhsAXqRWA4n3mIoRFg3SJKoOZ+o6p
jqtbc1PtPPGqhwMsZOL3lkfxPTUs4+dk1HMYLk4R6NPw6hnVM0+3oHBW3/YW3KD/cXzbwVtqpnAm
ZOXBlkjxj8jO2hOcFaCgiYlckKsfeffQ0XmqXG92YVxjuHSBY3I7rUkD6gTvgYqIFhsqZgjyWUz8
gSoq/bLUETsof8KfvqGCkfiy/BYTzUTtdACFl7YONAkkzQosnkz25MseV3DSlFnQMKP55jZj9TV2
9GHS6v0zYL4diiOdX+MkHDOcuVj2z/e6xsvaCAzSl9Apg2exV0NdTcIeHG6bKR0yHaUQwo9JT5Sm
9xo1wFcQzPJdxx0Kt9uPpuWs0MObVZgOpqUXE8ktD0IJqH+tx2V2qPGRX9rnv8Q9SrNlIfpa/Axn
fGPBDNsVMn+vk8ozG+tK6vkMiICv4YnFg4jxF8sQPVh2hO1l3AFtp2KM8WMROyUwmfhmhuiMyEVW
wEqPHav4XqK8HPQMtik4iAiEOKGDF2lV+xTDgdyEMgwLrdcdn/OMyZpqe1bI1GcaGsWkSOPfL3yY
HDEherkJFLIb/BQ4lZwPUD2grtJJtFMCOZav6Pwlp+UiGN+n1JsdjSf99h1m0bs9LbLBCXBBOsRl
vAfrvZb4IO0fB46l6AF9hFtyUiKEktNNEhyXejI08PV2K9FSrGaHKsp3s3iaCCaDKsRcJ3AET8MY
VyIUzdsooX+Ye2pxjbGCzqTVur0WOkrE3fzWJfONDDutix0lVT48Blkyp7ukIB9Y5+1kGxNiwgjE
PMYwM2hG0Oy0T2i1QMT2uX0Y8OqVddqFCvocDv4CRvdstG9Le+3RUoVYct1HKgwaMsjCSGgUMgsV
JXFPVXyO+iw/7yOkUVDZ0E12TGTk62DBJ9vaFSPl1fnRtDU9ioc8vFqUnipQcCGr8KhPFwh0P+5Y
6Ssc/0x+AOJ9FvENnWtp9x4nzDdrD6SWVWA2PXlQv9vBlZIaSuigR4R+9/tJCQu7NQ2X0wJuJvMX
A4mqf8ELOebNjZNC4jJkGtD+O5fy5cwTG4x3PqChDQ9JG6rGdMM3zjX9ZDoOT28oCWPtoDB00YmU
GNB0njYKvNxQRfhZyZCKRMLJJTqFroaRjxfeK2Y3S6T0ZQuEsSpapxKifZ/AWGqzTJHTzn7+9QoT
FRyfhCeNmyE9fbfq9Ycu6ob4puP+MOjZWXf8eUV62l+O6CBQH5enWoomyz2kqZRDjbRnBXmQwFK/
GcD2u3c35Oo3aIfa3tMcLtGT5NxxyMsV48Tdfyk6GeDJ1cDYRi2CII5bE7WyMPN5Gyyscvqv/zl2
iunB8Bo7QeywwVqeQ6m8l0ib3XGtMSXo6fSLYocbnt4EEUFpDosv4eNXnMMCU9IS51PnBidR3CG9
oXdwGVA8CKSgYeaOuymKUt4rD4Fny8zTdNIoSLhomLNqIzfMKJxgFQeG9KvQ/d6WJBR7wFdBvsKA
cnpZ3+tRbSHrnNOX8VjTwD+elgM9lYXFvkY7q3eWpXFQqHfZ0hKoz8H4rVd/vWiJvRYqbxxXWtqC
w5dwTEadxuLSoGhQQoBNi8GVdbzKwgAhP60rJcKjrRu/hLEpdPnEx7OFJmYW1+eTW/dg+XyBWdk7
Ar5KOBYrEVC6kviyzAN0myefBpU4ng2CESrl3iRHMGugoELsdGnUVxUw9AO/ZhXiluk4K53Fr699
dbg4aKTM2/kzryjP7fz5Q9AIiqS187ctIEkraaKcIr7LRtvJgXimpOliO3+Tu1HDptFyYQz+jUJG
G2WvtULjd/qfNMRMkymrT+bjGfCedoGEcGProRmYBFfiBWf4fDaKiBHTYPqASoesX6jQqwS6Chxr
wmF+ILKjRwiYF6iGVdTh3XI3JGxZlEdfHLsoJcsYS/9rhDS28GpzK2tIU6vGKQ6tyiVXpmwRdUam
ltsIO4Z2pQbfmRGV0uM165MiFxecl0+RhHzLORQamOaA90EwciTxm4qdd0vJCAjJ69nuclzn3kj3
pX/xnRTib+vHcYOABolbwaR1W5bsmGKZCIHz+CblW0rV8VHdU9Tp+Jdx0vE/r1pz9xOauQ9lYvmn
zCqFOoqwNvgO33O45wMG+at8qqyiqAtlON1NMl5AJg0APOHHTVkeq01jdAMVf8E3PwrbTfDR8y2y
gM2omOE3FZmCACL0kOLveljvBSbO6NrY2LTXXUnXEej+GCt5cMVIT8QlfnfP5/HWekUvEMYUtsCf
paesQGv2D0ig/15IC7OR6BQbMQqC9dMsjWTeoegr5ovo+kASlAGnCM53lEfVfuzLMIjdjSnGdP8C
fTp2XGRpRq2otHauZ9Wq1tufKoY8lomZir+VQ/UZZYquRqoiADZ9OQMmnA9yNfo2FLF4srL/Kqz1
LeexxnAlzOlgyK/+ZvYKpQqnut2hF6Qrk0sdzZcX9oxpWb5obf95UUjwNCxeQ7Y5nAujALHWxeC6
YFHaW/yUxlYq+cdvIfBaff/5wH9Pk0yPH1kby5wnfJDFLfNTQ2aJ+WLVvSyyks2WV8SPtTboQjsg
OfVMOrJElMf2sq8lNCyTjASDCW0Py9INZ730SNtxpevXjTAZmdQqV8pBLswuErw0noljnabxqrna
qvwFXHxTUyY+wt4d1Kr9CUQwGCoV70Ts87qSe7nxmnC342qmUS2dRIEpRARKAxyz/w0YHM0gViTY
5CCQ9xLdQ667aIeUbX5wkG6F2zVJadxg5AD13o9uOGUMqcLJ+PVANHt9b714wPv8u6/BHzClnItq
MMTFofssnDGM123Mx/wdeJECOthvxBYy3Uz+YNNNebNHicmr6i+1FlkYs8lCJcCtBWDfF0z2/7VB
mGALCHE9FKBldwVq/PfdBYSEzzxhpglZUruSbVVMKi6SfCjbVSbj0q9oD960Dss6IrAD8WuMI0gY
qEhGsNFvQDTdBwCNkboadIjPnpGXM+sqQJxoUmoEFIdn8N59lP7yIl8x+ekhTMbx0C6BqPIpXdWl
3WIabS+eQJK3lWUthvo4azZ0gNAsodJLTtQ1MmYQBSTFvXqWNPrU2IMpcHkTk681poxw/MbSn0ke
Zcbp5Z4e/xpi4PgSw8RKz/slZcAnTNAuf+Fzwkj7BisBnt+Pf00lveXbCUmCML8iefRznci3GDZy
97Mh8jVmQz+EMsBNR6gDfLjS4uDc7w0WWzJlcuZuvF8SYMYDCviACUvMFnDPTmsoifcTySvXYW5w
omHSZJL4+uNB1IkunhumMxpd0nyfmHutf5OVRBjWPu5ZsOBHe13FURFU/6JDTvbyxOD0zAm4VhDI
gBnqpAh1m6MQdpZMPjk7j0Z4kFSxcVpN38uKnhKtM+gelCLVgh7QD9LZS9kDHopDGVYqZy5VJspR
2WD/fIc8+wJOyKmMq/CCQh5MwJGVLZgtbuiTbEMP0G2xO5Xtydf13c3mqgYKO/cyqQ0fy2YSz9UE
Jq17mReDXNfQqZ0qZJG15sTNT6LoWQl9IbI56Gw7V23Dgpl0QiheBdTC2ObNwqQo/ttjD8IfJOjn
qM1Hh+O67t3pczb+CLLsuB1zu7kZvIRIhLM4w9CV6nWWL82215HyRVatIcazXXrvwdGcX2IbKTnl
aLBa83j3641yvjhtmUqA7OCC7bUeQHiG4WxoKSHS9N5uCcR0HyQmfYmvyRMJDXR2e35WVAR4f0mj
5d5p41mNLNWCGmIOLKSk//RVpblWKdj9wko2dvYF1x6K9SY8hnIBDZq5XpK4jQeeADIyPEfOGqnV
6l3vBBipaX+Rm2bWxbMKk/e+fhM7RYy1pqfDZOtyPDbxgVOVoqgJzh389Q8hplzusTKmF4hCsJaz
Y1z1GzWNGeI2Wdn739+C2Rsb76biJ5OdgLXyyFg3ONDtUT2aCio/AkbwrtONwvEetVYZZtouMh/5
Ehrap0A38hnCRZdjGUMYiTZX/We05Nk+nDcK8g49sNwrkw7PwJFlWAsQVZaelUbRBcItMgj5uKrc
ERNMWv6XezmX6o2Px/3NjmSamfuBM77ebspjP/qSApf0+LlZ89j1aKnunHXzzrgwLwS9WpwT5K4g
uWTB5znc9Nc5Ak31X6de14vauoimarKCn3/Syz6T9eRCm/Cv9X2q876LimxbEdvj98CjHrolnzXp
VIjyNcQe6GCfiEKzkJHlv/DwuYZZw0z1C6bNGS+dcSUKbSVTC7omks+NZQgrcohVAzZWC9NHbjCE
H0BZ2c6H3E3/mGfYv6kyO0dFjcA+sinrbyqG3i5u4HPFoBzrATI6mh316LXcXm6fP1ElAL5oRLih
A7Ms6jA0yC7Ep3SO9i38EmBvzJCGcoBLEWDx9TICkZmh+jP2+TRRc7Ml6fmGN6tI2rrR/ovSrgvs
u1T6YdLuhkclutdu707WO/cVcipD1pL9Ew6kEuT4aVC1uQXDYmzqaoy/qKFf3naje+8hMj/3ulC/
yGPvZfI2J23MDzNw6V+0MxKIEkOXSE/Oy1z40V+fRUn07+B0YsAR2V5NSBiM4eiSCQJ9RPjnJlTY
qLm86Ox4ZaU7gZbeatbfUOXgxa5qQfOHSdYF4uDwFz75RwTBrdXJVMcZ92D1OFLi56wdmF+dEQpA
+diCL3oOZWzwWE7ZLZHOHCYgIa1XiaHHg6bOqO+TBqHZhgpyRBu9ccYuS601qLRGN6C125afVMO6
U+MWc1CNUPTurGljIXJLexzXVtYQiJ8CNoKyyE/rEmk8ZnCkFpnb4LHQBvBZQqVKTg37IuvKDJa7
xO7iU0ZGYYkg4+RGn7cQ/BOWQfCeAoV+mD1ljiPUibL2HpDqgK5QCRWf2JuXG5c73RXzJUjgmMIt
WoQv3jUzTR02sfhtHxHuyRlG0s9r8nETRG53dPLoMOD9lRTKF4A34zi3mz295m8VT6kvdh6zcqCh
jD2UlphQeCjSV8+X2EK7J4ja7EyujBR3eZGINSIxC2/1axw/6K6e1wnxqpCWi7BIaG3/wMcR8JHb
8/dQg0/lThROqBcMtVULuOdKo59ZX7cGpCccKRZg+iWPjXdvvNvqfX+Zn5xx9IzoS4vmiMQf7jTB
qy/fRMWgutAoo/k6VHdw0drH6diTwA9GXTYi8K4jg8HmuNPu6od/J3MBI20HE81IAb210Lz05a3D
AzxwkQYfktZsu8bL1Q1EYNZOVpFYdaoTulNxg/81dOBU26KjZEzPZaGWzMT5LWZkJFDRRROVbL1K
y12ehhBvlp659zk5MvEX+s/dk5yhOBTf8KHLEVzTQ1yk9gfKC0up12xfLOfM0BZSAL3+kGM9h+6G
ynCbtUVKLPJv8l3+APpm7+7m/v7BwcK7JZph26Z/5sYdxDHNxpUhU0UJkWRitAf6bf9ZGroLd5jK
piudVE7WbmCP5xSChrmYp6cH5x8CABSVrgP4dspBx3A4ikAjBXC9EuWXaYWt3OD0msJo2pk57ETE
QV/5+VlmMaVO1d+w6I+tnQ0Ckmia3eYCcUrTb2WVzo3KUMF4RLrX7uAtA1S0eIrjy3CFbLyXM95m
Cs2+PSQaBGIz21HTO9w3EuUBru8ys65zxl/Hq3DM/9hmEA8njEqnjT5NYwXROUMwCQnUhgyW33Nc
ZeVwZUxFvUuGOyn0hzWzdc77lWS9UGBUYam43/TzsTsGTlrjQhVTZRyU1yHEIUGOPMcI/S09nxNq
k1quU21NDtnz2RLCgdcWQd6yur4YsP2Lj6G6anCXgvVwDJRI7xgnPPZoVsNttTzTY96in8jFoCqB
131da8MtaI+ht3A9M2dLFQ3xltwFt4Sxuxs1fzQCeiKbV3KVIUavDnB5d7KNVl+Ew0jLdElCPCD/
FDwvlUPQa+MBLAnIhBlLRgyA0wUwh9bPCV/c3daag7bLvrHfWCjCJaiz3rdYn+XI2IMy47FkzyXG
pMaeaewgwmN6W0F/JiUNRUMhMLlTD45akf2t8ARVtolNjYDovuSC1JGnLen/RqzxNctggXlopOpN
w/2E0O0+PGzkV7ALG0cKM4CXalWAzr/zyd2IR1EH3J5IQMAhqsP//9He0OZlxv7Grjq7CFzXqEy6
G9fCUGVvWKzg8tq2BmiPeHQkNjBIqtxKCgG2AHWyY28qFExaXo9PTvIb1El0VR0SYAbDeTTVs4w4
9wImkKZ6FUqACnsH6xpCXOPA7nD9Jh7o8zTnb0fDlYzwpUBGI78gOPV/TIIQv/F0kQrZSHH0Kz63
4/8XYTE+HqlgF98BrJVSH4eHelsdNVJJYNClpWT1bhyYoIrYn/G5l5d/jDGSS2JchwwxEFpzzCN6
Mrs0LOKGAciuD4DyYrXB06rq8nKMa+gwok2FfgD+P2Z9kcdN2afNMIoZYwAc2E+ok81LH8QtKWn4
Xw1drDqUbin3sEFFyq8dpfxpPTKadJlpmOQAAnCLHlpXoELlBPadBCl/iUMdzTgW5w3pYYVt+cmp
zHsH7CLSYTDYozQgzVA7RP/QWDYBm+cd/H7imqWYKaVJRcUn3oB9b4rZSnZFcW4Pi4w6g1uvRTqM
f0uTAJvj0+7QYcQnKksu9kHGEgLbpEsGpZqS9vMLlqdHrkRL4Ci/cRT9jmylNcSCc3By9iJ1VD/C
IvWqi9U+lSachC1rT3eyZ+tPl+UtPHs92Npt0sKqSjHtZCqJO3R2N/CCi3krFUnlGqrKl00AAZgq
eUtktypISeHdJR4xuseR+UvM3W/W/t/3CcQNhZI6iZqPE5o+/A9smMMMjEilNA0ttTuM/rTmtk+E
2vbrCfVB7OKk7xm6lh/75Po2SR3qXHMQExKqq2fQYgqNR1lZhC/cMdNH880Kv2U9rkQFlrJRkwta
s8VCyiz1OpwFzCfUiZaBlj/tlSK96jaJI0+6v6UkJRNT8Qom6q9tRaPBVup+UzlV6cJ8sT6R/srQ
ysi/FZDYfG12jAb0FuUxNBNmEOLGqKYek9NAE47YQSWLj+d64tp+0vk66Awz8UWpMGCfMc1uv4GK
9wKYwb5+IO3+DniXB0DV3/gS2HfEm4bpXf3eGCA2kcfYDkou3ibnFlEi9OewUy4JaHHjZrzSr2P5
SK3HoCqPZd6aKutvrNbYGPLMQ9k7J3mjSYcL+Hw72ZcphhCXvIoGgSRutlTPkrUxf42ISL2jfV+v
d7MnFoxOjpw51AyKJ95vnp5Mn1sfqf+z7tutHcr5+uT/gIhT1t+oZ9J1VJteXAk6HlC/frswcuzZ
6SQheyenJXHExg18sbK2E8KRbb/CQu58EDFMkWqlxFBZoN+zrkeTDIwZXaf8Rh0Z8OF16klTkGLn
uZ5TUVlmyOt3cQfNTd0qyH3kbHryR32QinA1rsPdJDm4UVLEQ0LU+XPkPz3g9TMXMasDjjgvZySh
a93tsAJcTg8yG/q9NdvF0NDs/OtdTUsfknAxIP1z0GtGwQaRmlQtZDzWa1iruQt9wqyYAyClCC0B
P0I6kAPzgpXUO4rL+SVPYs0tTsalgL/sxuYW4ap/IewCPI1SCPjeafnd39uWNc3dTDdFBMNWKTkt
j7mO/ZAymGsSJvzu3AlZXhZT8mq6mqXZDyMNNooSNCu5uG2RZ7bt009KKboJC7lTYLHlWJXe+1gS
Q7g/9rT3lTFUWJ9U58PNj199pG6NZrpnea+aUTW/FxpuBx662J1nbz0rUk6p8QQv6V86XI5U6cUW
MN2cyHrhy7Uoa3Lw9i902xG+oWArlCfzTXz1MouWHsG2FExFy5iUejDsnRwpUFagOSzaAwQ5whEA
5ADAop+e/V+fMzRnYB4LMawDpsJzWhfWWnfxucZHb6am9e/bs5FH30jVtbO8FON/7vGbkzffALhB
8voMim/X6mN/GslY3bpkvOqummBgZPCCMsfuprmtf00VAYH0Yj6yM655cD2xMt76Mle8UT3iEcTp
oGzAe7L9P2m0j37pgJtV3PeHghTVX7ooip1v1xoXHtXDw1MAFMkMT/42HC9yq/PJyKzTDCqf4xkH
+ukJ5iB9ZACuNi7EbYHxDs1UOYQnIy6u+bVFogKjwptoAra+rpRf9sx4sdgzh79poD8z3Wu/Vu7B
dfmKsudcM4n/OVdNoc1TBZHV0BStUJBhuCwlaVTdUbjqxPb4ur2kDyUXcLAkCPptmCR0vNTCDzfl
c1ep5iguVXt4RVuoPc5vYhZcwvNoxOWgr+GdkLo3ilbqJBBfzKdb98iJa/sgmnD9wWe1tmEVJvhX
WzdmBocON+lxY5nZunkT9I5cDOk5PVzyM/8fnRnqiJwN8hoHybhSBDTu3IwfS6fTaiS0hyeo9luc
YWiBweB65KsTWez4ucdl0x0Yg6Uf7kKHNlMGS9w6VXnlYzI46MP41XVXveHaFen4U5gk6c1FJl+Y
lqsPwFJitKA1fqmWydtEtlv0AMgf6tVQYmlMi309PGAWIkBWR4RpgE2RSutbJpb2LE+aoYwmMHT7
rcTMVnolnnYobtwcRvveA9EO1B4Q079t8JaZFUkIJnxcYHoCC4GNt5DkynvThUFgsZ6hfNk61z10
hfl9l8DxvClZqiDoOan+Oa7Pja+Z0jmMQxb7fZ/WxknxA+X4jwmVTHc3khOY3DfG9xR9PbWJuh/8
Baj5A+5ptyeYfEa7dn3DTWsu/DLXCUxup82H5QuMhCbIj1/ufhThpyt07N6+Cucc2N7Kgh4VaRbA
trR23qMVvy/uxNnQj7z302hsOUiuNB9cFpP4/cIuP2AZhoe603wGfMV8CJ7Za3BtIleoLITOCgbn
GnzvGOA9huh3/JoqGy0B412rFs5dvj4WffSHlgl5SAC+pHSN8Y5tsg0fUXapadG181Gc6mSurBdL
hndwGHS3KwRD2DAppSO5aFTwkcxxtdXRy++gRAG9gs22N+G2owEMuvFb11lFoPrsRy/PsOVBqb1J
QRm8O2mnBRpMmAco2RgP06BC62IvS5sAuS+je29Sqcwu17iXb3yKaSiQH8AUsfUxoWPB7tVVrYZp
LgOFcGaNWnizqYQ6EXaYT9BpDvUr5GDfUsa4OWv7YIkbPSXT6kveek9YCzZal2zmeHCMyk6cyqzu
WCxl+peRSCae9/NY65VvGha81VQBA6paVDo0Cb7GEr0sVB4qTYOhVdcwIgkRTku4UwdJheM8j3Jz
GWw1cj/wec2Jh3/1Hmi2oCatvmbUG5mp4FnYx8xTddsWiT5vrdz4pQXH9Z8HL1v8IuVErev+nmby
Erx7usaiHKSfXr/C56glNZkznmiktgIjO7E7xKncbKHXwuqSSt4VaF2CoqTQBeliRlibsPn931YF
n0IgsoufkePBZwPbqQuK5Ct8ij+axYdeEVeCXw9oUa9pZW5ACyX7HqqD5smYkUsA/3rdFa5xN3rj
d2bCFs1G7Vc5HXyoLBKV0+GMOUJ5cCYAPRKrBfY4q2ZYWJ97RKz7wjK1S7P/MJzXQZsWHib35ev1
RZtznzofBTmI/YLWqFOIs8vGd96Yi2r6w3vXRUmtl6tBCMd2kIt1jOaMpxdf41o/aw4yj/RU21QS
YP8dpQA0OCwuMD6ZYsBfU9w9dw18RPYmlbCB+4mjzjfDgnv/J+HsozeiY8Pnca/X1tB9KRw7d894
0z1IQTHyFxM6ld/q2CNEqppNCJbz2bRk805p0xRBBaHj/lSe0Lf+oG6z3kc1Hm6G89q1htwnXnpR
1pzjRiNSpfSpYgLX+KZqE+gt4eLksinLaCPCE/PhdPoxYx5BCAjoXKL87FxGGDo5TLhdfE2lKjWv
XJ43noaFe54bA1VOXv+019SsWpJg64uE7F2G3p2GQoiTqpa3DtgrKva77MtcIV2ZKK0/vQR8Rf3c
cMsJ+wNhtHfO2VekITtthpxYO4wHcwWCiY/zSvjsXLYmnOvv8Al2XPg/9j/3fBy+AJAskjCIJ4d1
ScT3xvn8QCAonLoR85OyB/RItBOD0fcLl7uqJjZFNR2OGx3Zo7G+0xH7UkWQuluRw5uu9Nwuf2cC
AVlmGh+WSiP2szuAnkRp95MKaXMgfMqpElE1P5zdtNrZXOGCQ2SUaCfPnQKVmayj2co31JPgoWKc
Zck1joTGwRPTc5GutDIObAlAm3sLftOle18DAvjFYLbKgRc5lPyHUs2qmPZ11p+QzOIjxBTOIcwQ
/z2Sj+p8mev4dieeB0Fi/DEDVC1/w93IL5ImEkAmoyGBtnH2KbKamo7syHoeZp62qOs2TXi//hTG
QLCJVN7cWkB43ujFRlquysyxS7qVaeOXQT+w5g679kGKFXVBVODB7shSApAarLiua3nSytgCWSCa
GzXW08rb8YMboy4glcRQ8FLO7j6rfc82sl0UoobjVqJAPNdbtbWGjQG2BffcWDMtgX2ilzgqIJw+
uquIEVQjKfse7uUbnFlAD9L0n114O0Peua+F3Y/zX6h+ew7yxQmje7UX/nSxyjLOky9KSt8BXDQA
xrZg8h680IOM2ulLRIGEMEeiYG+Lg+DjYcQGXjvRz+Us7apTZdbJsJcwY1TeiC/FEIoBV03gg252
FOUsCb+o6a07smRyjAE/+x5uK+ZmaUCM24kK+0CrDEF/WkVA/OtiN9dv31lslvqMrBgAOlEX80av
5PdwFq+kLfznWik/O1ZcMQQ8j87qQ3OG2E+2J3N52BaGWUnHeaO13Clo2Bt6Lon3JPN69LVofJzi
grkkImmBjZm2sII6IlgRTDM0YilMhbmNNZ7IANRXLqf8GjbOdAc3hvOAGQKm50eNaGSRQZLOwgCU
bMC0JP4hpk99EQ07m8JS/QVrabmYV2VhAzmvhruAec8o2wYeJ0BunHq/s4yDYkDrnbogwDzM3Ztu
l7W95bwT9yJNvc6Z2trtD9xHORzsKbkFOb69MLpoLVpfxNBU99KceMX+EXi+7hTZXWcu3dOZK/1t
rXuBszapG1jraiv5BvITyifYOtpFbklIv/wBbQU+w5RWesrye4lJN3L5izepdY7ciwqfrHKQGGJn
jGBol9f7PnNzYuEhJsEqfSFsh6nSRj1tdofe8yqlb3b1EYPF9t0Pu1L1bmUWDe9ba1j2+VRX+t/6
mIiwO+vyWARLCrsTnsY0t8Hrgs99mhshjTx+WPG6Xg6HtbAJGtva2z3rodxiajO4jgCfwiiA+Y++
lSpKz1S58jCyubjQ7w0ATbcuOLhEF2tMVRhZ76SZ81NQSpHYjBi0TF5Wmrq2HyPGvejnqPCxyoBi
dii+PmanhehsLxw6357FONO5LmMXlhkmwaizSxf9FA75cb14Cz7lnRSH5cGAh2rk7+NIGFaptE0K
tZMoMLu8Ab0oT66NDKU9FFOfnJ1aMOw/Okqf+0IAyE7zrGsflTpmvCB3LRvvzxaBat6kfGIR7cFl
WMNAzqcOZLhO4lennz2a8ZcsvHWbwG7Ukjh+CHzY6YL3VyyDCZrGBu2sUrCbjM0CGP1Litxp6gmd
tlxnGlT+XGLfmXW1TCVBGslxxr7OoZsBrFBZ2I8mh/tFPYSW6wRkxsieem2wo03PLiv/Aw4QoqmF
Dzhy8RpjEs+FoKk2b5/0l3n6Nj814xlWJgxcsam27fF8XTgGXxFWdSdUfYAmQx9rtEofyODSBJO1
X/Y/sYMto7A6XSeQ/ROzG1B3bn+co9atjmbeCowej2qDPh6RWF5fFMI1RVdpSrWFvbn1tzR7fIMQ
WI5xKlhtdq/O98fk7szvxliPBPZ0hAa4yF6Y/8sB0bHggM5FQWJYzWWqfWWgrdLk2aqbh/XChibP
3TF7jQugN1lWOsRGszC+VwwudPn7FHr7PD/T9MEjjdF81ScAmPeYKWd4BTALwFWtqwDIjCjTkkBY
XwmRfxVYcNa5hLVPdP/L+UUEk60CL8vstLKWO3qPkV5jEA8OIGlfzA/mhQTXZZMLWqYDCT2MnC0B
CxpDROGGMNgQ797hFL43GzJuJe+S44pTNHQrcQCBDJucTmAhQkGkrRIvqqli/xUouk6yrneBeqwr
/jZgNfNULCEK+hXcwU0E34FAOhwwjb5FOFlafPoZlC7eiOQ121+3giSGd45TQusXCgxrHQA6WGwt
qDqyDBaCtu4Ls9EHeAF1la1yrM/pwghfD1KCyq8h8kCDhm88pV/LiYPcQ5k+Lpci/Yu71LYLGsXj
LCN0OBtMutOVuVWg6spTP8l2CJ52Jee9Zv48uEJH/A4CJt04VCBT9K22MJ7w30tygeAbJGXbq27C
gvdCgjPOuSaF9w/QeRJv+8lqZkVNLrmIqs1RwGH12jPF7W1JsQlhQVT9o/DaOR5oZy4dEsT7Pp0d
VlNSRKm/+ZM3BGXc/AKbVom/Dt8ixH30mVvkW6iT10bH6iAttYl6/BfI94urBr5vOg53pJBct+/G
28QMwiWCiZpi5DC1XQmnetFRxPGJYn45njfQE/UyDkIVgoTmCNUJsb3YaAj2Q0i7PYRsKYs6XEsv
qoy6441jH/En2RNdLAlW+xD3wy8a+iinF8wm8xXyvWluLX6Oz8jl9v7d4Fc9HaaSzDM8s7DT3DiD
JjeUug2e5BWj5KfLqhYUYPjpxzHEFHhGAxUpBKWjiYKc0TfWXHI+Nf4ClwxS5cGSx8dGuqQL651p
pTpLQUSwJXBtzkhgM3A/HJOXgSkROLAEQp5sZ/nJm2uFOepnrJX+ygr3b1d6McdCcF5rEfMiuc4O
/XdnoQU9Ge9ema7jL+SL0O2Iefr0SSRV/6v46LYFIp2jdNLkkrGEwAATuWaLwf52Kl+4A3vLB6e1
yWiC09GIRzHqIZlcamPotj0BfHnDiDVIdaC9VM3Fk06BPyPPpAOOgjnjOSF+Vb6CnEZCVLhhTcyB
VSYdwIisAXBbdi74lT95NNKGFgHMDCQJmyb16n7x4+a6ZBe6ytk8iWtw0iuh/TVyBvNanejBRV9s
CheLk6naUujnbxtzxkOX30g6q+l+TMRYb4WWaEalq4u/ca/npCYMVVq+wncerbNhx14wOsXpyHKm
7/41qf4OXsDN2e4c7aRUCTXiAU3YqbomenPqkBJh3KkE/gRziB4Q3255hpY97BpxcLCqGOnyTY7v
ejgYbHoJcKLuW0S4vIDHEBJN0wH8i4bg56fRj7u1EJsPiCHCcer4+ymsCALTvBLkiWauBtBHUL3M
tZazxGtkdU4tFqU6ogh7DHunUx0G7b4kqiid6Ff+fCDFh5VsBoeqqc48cm080HQ9umbhyH6bcYy9
E8EGEyxqYiKYU22Mmr1QtyTAGmk6czjdfKDtoBI42MVxioiway9j8y9sGauiUtva9Z/q8HyKI1Xx
GlJK3/pLKcT+9g1zAratNhDRg5yr0litZdt7ttp5ttaAwP8YKYtVyJMRM3kuNM9U2ec0BfkXK8WY
Sbx9uNg+Sf/bVa725rDwnbRK6HrUB5R10Jd12TRzMY1qIAWjw97tqixkgPtVhxYyuMsIvi8rgfi4
2MaDZSWaCKfMFdwL83bniIkk7S5SQSW98eoRnn/SQHBNeJSdZtIbGlyRUr94GimKQNy9Q3gHs/vF
ItQUjjgXE3KAJZ4g7yO9rdT0hPhROGj4nOP3MH91DdcM+5LJ4cW12SW0bzm00I8KpK5yM5rJEO8s
Nw4g131NxJVngfPGiX5YsuOcFERYWnzEk/AkDIvUjG7DaHlmp8aNfwzWnmjofRJaa1CLZMmTqn8D
TfaXkdPk+4e4kF21n9ILi6gcwL3NBb+tjfWEsn7WqackMeQQ/W9pCA0jHEpDIupmdddIvB5ThcBs
+YNlRQpUKJYBLBb8DLd5PNbwFEKMa/ltbj9hdRG4lYTHEBn4DNYZG/Npsvybzf2bPEK+ZPQSKvA4
ttE1bprcOPO1T9Iz+dguDKJh4hKDue0/ZMwXUd6bdVxN/f7Qfw9TaK9/RiEsEa5nxjuj6ooGYBcP
OTrwl6vzVvdNqGAJYglKnX3nFSZLhp9oMK4yEpiIvCL4rXeAfiFR9jJF8/Xtvik49OPucEqa0VHS
Ubg+2fG0auzh5wxnloToRVm7+oD8/YO/k4FgONZpikx7WRigBN7BddWw30xpU7s8qV3mRkGALGEx
FuO82G7Y2AZvxVbJ7eVAope137+t+EXS+I7zhGitmU6xZXPQp3xjcaCC/XwIAxXdsaH6D1fEOH8w
EdiHnWNwpE0Z6QC1JCHvzN8EFKRl+Aib2Km7vX066TZiZJndAJod6uVVl9kPQ+Y98MbxOrrA4RiZ
wmtkyZTgZaEkALH32e9h9fZIVb4U70MXCivejrJFQnl3bBY0RK9lQOc8Snv/3dHJyb4jM0Ncqjbr
qhgTMTDCMlRT814p5Dt8gaBWw44wE2gFst5cXICtcaSCjJndQZ5hjLRJGtNqbK2QJ1MuVFBV80oh
cDMhLSX+z1PlGkMKDVKHiF+nnNP827uRH/S5ZrpuU14/0/O1ONdw0VJingihe7/8E+CHKJi8gQdB
1IYqcPTRvTmhj2PWfSFntDP4ZYnIigeJ0AqGLxaKAtG37EJttpTVxQpz//QUX0yBYhk3w/tC/WqY
h5U+2SG/xTUEtzd67qG0UKsZ5kB3LHNJo/dr6biN3rLFxZa5oFUTQKh1d/k2QJFmf8EhIheZQmMo
b05ENNIpX/sc5g0oPbhet6AD8B2MIY/AYH+LZQEouRuwt6MKavneFEymxtA1SjfRIWIIFtjOrt+0
gfQRIo3WlMAfPqTfeXdz+9/3e2rkwsw0fOcCob80KqmjTsMN931uIJkQS3sdliri0/wNhuyYPD3R
OXe09Zp02Deor/WKlkEYb5qsoYsj1QQqaKn2OpxnRB74OEbe9K5RTiAq+lVm50Y0A6WTLNM60abs
jmriN2zRZe4UfV7n7Ys/lZZBS6DLmnc6o0S/HA0eMaxednW08QRZG5RS3Tspwif/tTgYk/eYdjuc
yF+6KxIDnBzrm/bCxQhtGnhNscGG86NW9imPzCh35bcBOtA90w5RjKqMv0KXXxelyef7nopQXSBr
VjQB7EQUTXBPzKG60jU62Nn7pQRLX2/G+1mGUwlgH8dX3w71/Cm2cF6HaYCf5rjPRVW42M1Somu+
ce5obzhP+u//zZQKOgnHasIbtMgrIqGAoCC8plG4VELjGou4CICTLcCkKWM6O6fhHFjU9DuxuXdT
stinuTMztGyenE2dkrCmH2gg/LfEC73HotZjfMAVKogWxUrVsNqh+OHtaTj0GSM/HdQ0tY2yHRdf
FW/BgPFPvMCutf3eRnxqLgvJRs8e158dnASReLo10y3TAvakJLBGzinNxdpmrb+bSN/F21Ida+Em
rnZoW789p4RDsY1/pqSzDrSqGOAxvMDUT7gGUxOZIFJu2naeCptWltK5vnVi7uXlnQGeFfBjlWes
iKcUweY2q9SJmlP1lHhAMWVUgYjac0IeM4t2J7R0TQNiasRrckLmCcVx58B24976/mCDCT8CovyK
txEXpdBSyT+bZvRPKb/dCvCTjGdY6dO9Md0k4KLruQxUSnFew4aK2ShPmqk5c3PiIoqqbWZiH9GL
RpEcDrBnRlx2BCv4oXdH8STwXVtT3sQUDmYNpt1l8Rc44QTcr1/SU+TjNDEz35vO7oMma+IRwg28
DhBJHH/HXkZnEvXZqn/izG/c+Ju2Jw86PtcEICmbn2qePiV5A7IO3oSYwd76PMDDtSKV7AXVjNyf
x20rmn7bBEXc5auFZCLSQTJ46PPrCawyp5NfxB1OFTALBnFmPFvjkBdqY4gcu5/c3VwxK1vNer+S
d6ps2OFT4jfg8Z/DppQMHvRuELVXE3ovDd7wXMn9YqhADGgH4HL9MUml2WT+kyqwycghbuQj0B79
EYdbKIbq36Y1DdCv0nPxHRstv/QnUblpFp0HxkSf6M9lQiLSdHmAwqxLqlKDTImJFTwE5Ag5FHLC
4gY67AmvxPaAjHWXB7mp3ESllpcHnmB9mVQMtLgdDzj2/vZ4RTxx3f/wowHRPHwIAwK6mbSWaKbP
/sow8exZqv1aDUXAaESASJncj5xuXiG/TLqR/MYEYgyvDLgOwZD6OttotPrJ9jsQ9RIgzN8pmyhR
drrP7eJ1LyQU9e8ev/b2lu89HQ/FZGiJ5ha71+uOmkgguxNDzvl0OsWnqAM2rnjxTltaCOQeVAlL
n+7Myzvw6wKV4J1o8gX/h7RtS0QhK9yrGHIwQHiYdfw+zqbeEbVWfufkPLkmjE4/U75+bstF8Bll
kSVrtM4eljFCPpK0OYnKbNFfbaLXQYexgNjgsiXSPTta0xezgN95zT6hgQoDHVNA6LUXRfMax2A5
33GpYZlw0GSvvo54mHg1sE1ma3AMxxFSG/0GvQoCakpSbfko1dZC9FFGyCqhbby71S4d2471Xbm7
HvI9MhHkPbjGy/S9SEHOqDIUv/pwQvbupYN9ZS9n1YD5RDGq6jImC7nTGxJLP18jE6wkqqmbX9us
SJCXg383wiEa0s6edYBU5sm3fiwXJIRekHsBAtAmv2dhj4FlkOKx2z4mT1lotUXLffgLbxYFOFOb
345oZe8sgwWksRH0vVDq1qXq8pkZ3yOmR5ArBWS5C4GDU0DYh0hi32DhvjUbuQ1atnzONlJ+rdpa
Ql5xgLvC9XimEwrwCq01jLy0xzrO7T/BuIu2KpONUECojZu+iKsL1TbMC/PoMDQh9+b11gGRwTxP
uFEYdckD7S8KHl6Ibd1CvTJk5QVPlpGylBXGgDi0zXcvp5d40W41S0FsW1WVUjSHeqWiirrmKAcy
3E4udELbofZBbNALcZw22k8eWp6G6aZjIQUFRFfHz3N2D0sHSRLzZddZn6w8VXRHulV1gmKxfXCl
x+h17L0tMvjKziZ4tLrOJN6WsK9odG1UMIbc/yNGZaIhwONpXf/OERpK2OUfT4N+DBfFt+EB5jBx
bgG2nkyFj1S+9jsCmzXFq/Fo7tMo779EVoLT3EZlAiKcMK7GXlVkcBc4dSajjYphi6HqKEHmubYJ
NMJL6gXTZPu4Ahvz+KoAWZGjoHJasOG7cqOyL5M3ikqpbsicOWYjO8SDVwgWCQWNjSKQFM6YNSR/
CpkG8SK22DGkLfecyH+01HX0VxdLyLNkzMUiv8uWjDQV+F/SYBLNy2xRYcJwE8vmdRdLtKOCAxFL
hsgH8O/LfDE6+PdBId+h3Fc9TTzzHfGsEsmRdXA9fmn6ie1QvFCkEW9r5n3/YdiWNQUSNGwhBQ2z
bcDMDdum68WmqXhf0VpfStpFHICvPihjbtk1qSxfXsKsY+65MBwiv10gJLHLKvbtLnPnBoGqgfms
dTHrzHHQSEeroxyq8ZLomAWUaCSftdXOaV4QUpV5OFV8A8jIaUr2AGvkYv9XCurAYmQKEXw4GO2K
9qvvRd/u6e+PLwnN7iFDznW7i0lpe2vmT+RkWR0OiF3uuLJSCrp8LZ9sWryYKOzIeO/w5uL7XHT1
GeuawQc7suRSI20FbDtUwx4EtXQIYwS9/ODLhN9AqOtqz22fzaWffrr5RAxBhZ+1Vat0Q/E0D63e
1teljGyaQDxkJpgqgBjhhDiNUH6dpkafs1KAlOl32gsB5cTzZngEzxnip+f8n8E0M6rz8PtFMiSK
BBp9HGXt318uEFTW9zw6oE4Rm1ikj9CSdIsQB8pDGWDjxCQvCg5fREcOVe8mvr0zN6w7cErO+gVH
i4yY5tPnCc8hesAQeqrk/OWXaUX+8HvgWGbl0181FTkgO5CTBLY+08df95KY2oJxSAwXGZdFk0x0
PXXmanHCpQDwFPFVlOGD6Iai+rSrZPkCVEwcKq/9MgpJ9GH+mR8Wlz1J5rJnu5PJ79pURxBAr8HN
Ff2dS2Z9HUJOUsnRneH0HiWypBnX+xfB5VxstzSTomASiHQ5+CYbr8qo2I+ccAIRZZ/kg1lN4vEU
XTzfVqquHH8MVkYtwrnzYNnyXIGW53PgT7lEnYfs75C+6+GhrzQgo92WQsGepxwwKPwgzmFX7Kip
q9UG45T5sqpEj9k7iz09ZrS/nxhzEBr6POew9FzxOwUQdriCX72ICOV4Ym11IO7PCS3XTDs8ip+j
V1bnx9UG9OMiOIF5KkO4jL9zKIhwRckn2655CaTtwVllxE+plljVAztWK/gftjTBtEIfY5NBPG7u
wGPrB6rrHglJnbgvTGG/vUM98CSMqgv/LJe7bQhpjdB5NwJlGSfQqqKYALN5TyIc2p6AVhDz9CJK
avWvJIcXSxdM7BddWTTTzJW/g+iiYtTTUHfJtB45ApqpGfDOLeL7NiKPYakQPoeE6GvbnQMnm5PH
Fyizx0LkoDWLmj3xv5jAaKTRGO3rc2/rKydimPkayLB10dFhPHJBp+KSPJlVUPJYygMNRuGTG5MY
vYoVHR36G+QuqfocBHkMXs9bC4o8ys87pdqqxC4aP1E6sPHtWB5lxRn5bDGVmblChmQzjMcL0oQ0
R0qDuK8oRFF3s9s0QdqdWn359SkOZnOsjkbthdI7WCIgSwLHBsF9Epsy5p1I7st75ELfaOnAoePT
7x624Ls4ghVMfT4pMRunhfD77YcYZjOLxzFbf3++EsgeTlGWc/ol/KxpOFu3Cie4Ju/OVeBT8czR
jWrAKeZ2VsVeOJcsxOZ7K1cWKdAFp7Rmc25Qcdw309x6WQbr//i5M1PsxA3oRyuCgxZjRCoRpmoa
CvVcF1V1oeP0KP/yS1g0glZx8ggWqMuedj/d4Wqy+/J5wW3z0EH8l8hUDF4I8O4ZJaAhNKChrn5f
EqNcKQ81w82xKP5IZ9LBSFJrklxtXXkAvlOUkSg1m5AKiZAdo8i3N4wVfIsdHoxDY4U+67VqQAVN
qgjZGdNjuS14wf3A9178gb6Iz26sA68LR/VKm2clGRAqXUWx/GZ4/vsoU//MC+Okj+JdfPSX32ny
kNUsspJPDRY58hl+FX2zChztcZ9JSubTZEbBGh3UpG407N5OKwXljHCsT5tIk556eEDaSug5up/e
2aA8qlr88OS2V3PLYNXoQIxoCz25Hr4VD+YvUeFSQDTgPhMX5DYTRerO+Y46TX1goATRxm49z6m7
LCRqWpKQq6IC5jQ25NBwsB5LetkCzJhIX1hAY1+MqBBxJSk+84xH/3Q70c/cH8j8LB5SHSxe+5Vb
iOr7DMi6edjI3coTuhj7miTKYwySSk5Z58WA8gXfvKiNDWAxH99jtmdOeRmeiygdB3ffgMWJZf+m
nwc2w1UN2TfHFU6GGySz3FDWu3SHz2uwf4E4C+vAhGk0l+WbgjbAoG2i06tXE403Y4SGZpn0AJjr
vQEd5HajHEpaiJSuXqm7tocDO3JPcoRgVfO9d66iz/ENbHOZpLUby+seYH6pUsOFCSb4uMURVe1b
7JQKgfr8nUVlJaZB8MDAq1EuZSAJvnMt4E53P/VDjziqD/ax7EkG3Li2UVU+R0ELOxie7WtyhDcj
xOmYbpmvFf1Eg2M5sAciZHc5XwgM4e1OW5beYP8CvKxMHL4eYa5oV2FyoRHaJT/fFfhK0oFIfh6r
pYdNo/kARqbV0CYLj0OtO6jiY99bKmORXQOmgNUo6sdGfRucLOtj0MThOTzCbyPE0vLoHMhveYLL
hpzCRCAGej+N8XEzFdRj4fDd8wJRgr6C310C2qold+h8FAJuvM3NMuR9nvyKqcnZVFuEfH38pXmJ
nVBWBuoqeMtmB+NpdB7VL0u4RnNbNOejnWFjUnuytkfGshJ089C6bGYzBSAD9trTOqLOg7tdok3t
MkbxtSjYyIF2PC42Mh6lcoUAh3TXoVxo+775IyRDrlnWRBmcNuyeAuiz542phxdO0gSG3z7RuHQH
0R8NDSXnc9QuaIcumCzAWLv/lsM8rwhASzlK8iJ6yjbNsMAS/+IWanGo0mec/xZ9KGEwYdCKHVk4
3H04IWiwXx7it5P6bUK2Ouzwzw4Zg+a7ZBZJLnGGpfgyb1neCgkJR/Jh5e9uZr8j9RD3uKVOFkRH
JHhgMQQtI1t6PguvwXp8hR9vVgclrjgxlTB9z1BMUAXfQ2J35Dq2CvCMGpoJ6M6GoolO5pUT9A4B
qcL7ymS7U+xwdMN09Ljldn45i/2IpLv6jYbMRZ8n3AGbGmbHSpps3Zpq27aE3XXS0hlj20hE7Kl2
CyfeYspQflyqc3Um4QS3yF5p2Hch7+nKEMeAe1q7jZKTwv67AaIImVVKsgjgd+euePzqweY1DSYB
KfxnhCquoit7ucgCLE1uygi9WAYLmyMOxw8dEXggtRxrxngR6mKEaiTULSr66Tgds1EuXvmPA2U1
bcqLavtGPbA1RyOn/x5bcuBTPG28BXcekYEvEPyKcQQ7jUkx6UQlGYzDtrjW3aj9PxjYMtVqdRnq
jMzmqaPoRA0YM2nwfNDVdeQy9Q8zsDkS67PI7q6uiNLdDmGB5gEwfXYZOCfwJGPf/VDP1Vi21j69
N+4ozySpF5xlAKRhrw2yW9tQTrhlxIfAxNCq+BRgeEmZ9jW5LJxrXbBqKH40/E2rzYnE4xtMxFia
PduDEbxRZSckAtYDJ4Z3szZxGWHkHoKiKcYtsR0xh1+XftZzz/YMmNqe+mcexC7LG2bXE/TSSgTA
7yRDpoxUh/qXJq8r8KsjjiMb9IRPqq1/1Iau2V9fggy7LLZP5WbMsYZaMsn3D7yzszbaFWt4r9nX
tJ6s0IZT64E+z5CBotKKy5O3bzg4bNFhLHJmzHiVo1/IWkQr15Pa79e7Vqju//o1nYHHWg7LqU79
aRGXJ5Z0jgCccSd4vJ5xZiynPMGIASXDPXPOxdPIh4ZWD90RYYzx7v3Vgr3yxncL5XnZw4NzAQus
VkBMAA8QZZ8hbDalb+3zHh8petk3ahbqmNJ+TKGMcsw89DkjiQht3eihy7c3GPmb13FSQV3uNn62
QPjWJc2R7Jr5JMw4O6zmICQDZSTVj8+qhXP3bxTSrxTtesj2K4vjqKH02kuu1sAvBaaZ6FzQsVe5
YrBtuFd5sGIkRIeyJw2IkX31/xfWoPKBfaL2zAfjsp/IUuwBUE6Ep7CF/HI/OSzh2sQEiV6D4h1E
7X+frPxNcKjhlaISkEkfeyqMB2jErQf0YYu51Yo2gnUCDoxOgoBA2ypk77FD1N1IUEoPL6FMKnjt
chW/ugED1Wb5lx4rOmNGvP9pq9v8DSKumL+B4xlwJTqA5a+Y0kx2qr4b6Y1O9vLp3yRCNLlD50c6
L+1vwooYtRILGZmxRITXFpqHB+htXF0ULPgFeHmuk8XQldQvDPHOX0/OaAWRESXpF+yF+gy76WDf
YMbSgivziO+mPtq8RTcDjoK3i6BK8+fUe6oA74ax/4dWFqZvIFbwi00IL2SknPJ8g9AZ7yFCceUr
bdvfwMlabaXtbTW5U860OGX4+yOSucdBMDdv+ZAuv3tyvvCJWZZ39zssPJOqTmkF82zn8MnXB8Es
zawF3c/XZpqlJwuZ5xGPlKPjx8P8NB4ko8qvLXkkV1nvqrgz8Y6IfyidbcsF0TXLHmul45/5C+UD
EOhZfvTzyhL4nExfHjEqHSw9A2UmR27llcV8Z1FmkT5CXkDOrPJkT6cl0CONUWGIiL8/Hlu8jwpq
vc49jJAtPZLud9II69xlYQK0shOv9yIS3Us55Hy/cDozBrDuNcEOkkvDHzI1GS2Izwzcgo0GVPn8
qWutcycz2s9JpAQRFfVwGpJIuKc5rfIX+qEJ8IsqJg81N3CEtecMZvCvUyjVtydezFMImijuc3pb
+QOhIuSpO3aJR3+N78Eho6mJxF3TCA1UGaXxYer2NqARgDDSk6aii7pJjBdC0bRJd14jgzuww0pU
qPSuEBL3qAadCV/Dv63tnoQ+P7hOlN9Ay2i2nSE1fqp4S8N/217vN5gGUbfH/547pj29gfVaWxn8
QvytlsNh/V/tSnsKwGmJmNpdzwz09gqDSBtJzyd5eFU2zy671GwvIffDOV39sZY3RbFIeUCbfomZ
jrZ7h34tTqPLuESQXrrXr+8kUREVhIpng4VSS/AzAf7Liw1IFOzi9Wc4mXtScm0a3fzyNYWktmfm
nqnhUnXaiJNWh8sVP6WCexfEyuLYWd5c1Hg96LCmhLu0JvjhLhEreVXEU9uYcQ2nQ2XANbhwuK9u
AK0uJUEKJ7Uos4ICigD4xqca3yLnG3o46dN0Fp2CGyo9f8UPp1rdSuQHn+XuIW6PZP8+W28y60gP
OeBOLZGLmRi4i7w6+xI9x5mB9M0VxZa9Ny8fvYi6Fz49r84B1r5hsN83HvauHtuvvGnA0US1P1/n
KHUdmQ64Ze/MBvfVrsTdzLsd8+i66jvq+i8mk7sNDRBlN/M03pbfT0t/TnFD5ltw1iwYR0qwFQ0k
VZwWFkznKKpL1/zhlntaqlbqbfqQBo5rJYrT1Q5boUfJ+JtQzHcXj5NgXUJ/vriYuc3QyL2NTEHM
2VxVhontxAF9/KT3w6w1VDXg6XbYQdu1XeuHyfFWIo69WeHjXdGy+oO9Os3aYcQgYpokCRQ7mPyI
haYRAiocy+miTeQimPhk+O2Mps1aFxuFTkt8xTnYmQjEIMFrSEijnQyTq9pWAlxin2GgeDUIxvqA
zcFb90fWwaYhwEldtNVq5+NxVbXcrid5eo4c43spOfnTEcnnPQ7mW4HZ7pufVTIeOqkhnbhWhBb5
g/lJMSBajjSRZTcgaYyKFAXo8QcKl3v6wH0b/9P6H4narOtJY3nyRQI++qryPDo5EEaZ+HUltcgZ
7xjpIdr9LiwlBzAglJqvTM1cQ+VCGPvhTbH2/m/jj3Ho3MtCdlXYZy/xna8Bziv2vrnSau9bek93
R7Kqt8Wzmu9bpVfYLrYNWqPD7wSCUsAtyE+3oPEvh/D8qbkXPsw5WBm9Cj4qOD+v0m5bzlPft7Zd
LEbVa+osqKFn/FhBzPILXUivpC5CvHy4BsM56TtOUn/t/bgCMBNfrYpcu3d+YEMHJBG012XxtKAx
OI/C3CbiNtZ+MiYtvfwJlzlrkXn9P8rRj09KtukOsRs+oywrM1aerG+Mf7aT2rhZbuMpNAbIPj0z
BrUQDRADjpXIfoahonqFqBFaRkvhTBXoejuY5kfaelryUKIacUM9mXn5Id6LoJaRQ8qdDkQrMhbc
W/YM+yovIm+EFl3rz3ZuOkP/Le5zCXK25ti53hLtioHPVhBqZ+c9RasaLRUxF3qLtvlRPeZtyht9
TqaHBCdquRAbNwjwgWAx4GnXW2qEKJ8D1c92DBtcFKNjLAsYOWkI4XoeeMZ0CljIC5ZygdwFp4oC
lDCenOfGZQy/SLCPO3eoXKyXY1RKgrAKkeVYRdtYj3C22kZvF/ABmgqMz2rIQVxV6IY3b88jwGFA
a3IragwNhI67oM6IIQx7ilcYTQOr9tzS4q8JLdbBb1gDle4oR6qeJFJwOggQ1nswqwvitqAA3uYr
exF+3Y4+rvV4FdRfW5+cUWXDvJtN1pKIfq3LXd0ZfXOTTSiH0S6Q7TlZrjPyf0EAFeUCpXFptlX6
ZqZ5SrFjzQkuaqSaP281Iml9m7aB1NCSDnrNL1h9uQfo131KsPuOCZ9eeJxLKD0XCM0P4glLib4W
pSE4p/j7ty8k59qxt5n2IyEvCYX0caTmw7+0hcGjTUS0myVC3/RBxC45aN11eZzbTeJaRqgkc/P8
EVm/xpZRZIukEI1BHmO4/IPyjpGmEy3yfGQV+DPPyHhMvsvoRu7LZnDdnzY1z5NLO7GSCUC5YAtL
bDLszhRech3q4Xc1NmSzCi2lshzARkqZ4I8BJuursE7FOa6nhaU9r3iwGFt/2aPCHgshhcVI5Euj
GhxlDUSj4NFGG9SY/gED2dfad6eRR3LDKlQQVQj0uMVyUZIFEkHQuUam71IKsIC5IfTFUjgKeD+N
X1+cgsVWC28FviWnAmsWe53Dfc9OsCPaugJYvKfoIxqeULHLeNGfAhq+Mf26z0I2T9yMQqFlelkW
PAECWxCNnQEeuMPTlvN9AQ6hAGI6I0nnzdoGr3Mw4Qyf8ZSFDyscGdEvUpumZhKY3Hr9fCLHyQzh
ibjw0GCJ93zeUCOrRPF1IKbO79jq0FSZRFghjHNci/GsStaXjbBS8B0Pi7wpAvIXRPC61bJqmp0N
BxXJvm8Yrx5l3IL7qTisbU9Bv7rEqGYG5O+hJm8J2gW6JDCXxbhH5+VJ1ZdocYi47rULzirlZ4Yx
wcfgaTv/shxtdxMgd+fhK4/E2j1xOipWmAXjfW47c+nB0cEKCKnEmcktfX8jV823lWVfsts6SkBt
4rlbQtX67uER00AQ9JA8LS6+j71iin7l0kJLFPPgltDWZsgeNQZenNzZahi3R+1HN9EwZyoTkYOL
A+PWwKrNZyzyOQMOP8SnY7gzKJK4styeU0XOTud8cXp/NdBVE9GEIFXixZdoSIjUPUJpzvFzQbSr
XW3KIqxOXoGS7R0YFWGsuUH7p2RihUY65NLOG9aWMPiqJavfnZuQ79HxstgIjj0e4qOs8uvbsjDZ
k7xEsJHsDCcFlraFAv87r8M6eQSJN9bF9mWpOImXNKhL55GaXlZCic/KlVA4hR+NX7XSfULoa9L+
m8yumSN1l7NtIG6Ja8EW5Qb/lFYqO+7jF9jlPcfPBwJtxwjnbzQhTuLUrLnG36eqPdHhzkeGpFKu
Ol0N8HWXLitk17AlPCgZQAXoMaRT+hHzsELV02IvfvRjVz2kiwHWBoPRPlw9D5hE1ZQ+GGp2xwQY
Okg0fz1emHpQ5tVr85c9qlqTvZGclDOOX5uc592C7s+P1+Qn5dAGtQHql6yf/Yazx7ddCRuEYvqW
/bhaSMAuF+V2nxQMhTpDlkE8WlL9T7ObZygGu1a68KOpLjN9wWdOiMe4RalIRg++lFYdM6ChO6As
tf3v22meFnED30K6GWpuYd3HiQvbd/eRBoW7rgsGnIwnmhAwOOA5kgggo+EvmiVDkDZLzqwE7P3H
UZ8JpiB2Bm89dpHJ1387fEIhswVnEUyw7aPYeoq3CxqvJL+/ZXVCNyw4oJXwSoIMJNwTku3HekG1
5effQREgqnG0SsKiQ8lNyq47uOLaBjcP0MaWqOT1kY0RAgx0mE+fbok0VnBZ9IDeKEAFMbWlU6O0
UjReZGlYy2G3ja52hRJODZ2OZ3dSEzl6VTck9PHoJv2M6YarEtipoY2BP8Zi+o5+o4MNmFtPJLOq
jW+VpqMYq+MPT1fd3uMdfTBfZ4sbGxHoHJ4EoudVsavxUXnxQ0leeDUFx1+15Ozdu/NFdusnvHv6
2Ra/zopCJ/JMVlQnOICM4LgvQZnsmXLDTLdSlqQr8cgU3ib1k3OKoHfsGt26pdCHZNRaKX0Oit99
+8ZjX5huebtmDntJZ8s6DieAUj7ARrgLhHknSLnEE0HWkCe3ksW/KFsC7tgp5gXNmY/giW483NGG
HpAiBmFGu8Fyb4aZMipF5RPOUtLVNl3GhUoD1wRLnnlsILkJHmqyBbtxQd+RJh2JDw1OS2JmpFUE
Cn6VpS3rpgu2+qyPOry9tgNAjlK5cvTCVdRvly21l7A07iw/25QpZC6zD4WCevG7umFXacwQdHgl
j3Vfg5CGNQ9+Ana+bC+bfVXLsI+hysyDlW+xowcLGGC8uN1cLKq3+FIZqEmaR9nNlQ8r67Gpualt
Vn9Ry6DwjD+WdhPCKwINhbsL2hIIWuR3nTGQFMXiZ06WVf3bjt5j4cWFnYLTDi1jAvp91FtLmi1q
4V3GU8L4ywXEX+gfccnVm0dXzDFzKKRTTtEoDbWNkygyoparEQrNrxtiM1Vn0gpCDq4Us1U7rFYg
9bxOcelPAKPrjK123P6zZ7a0sSwi6h5Vk9I9KOIhsiPJhTKKedgHP+5Yjy+b3q3U2kp2xKHJrhBI
NELFPkjiRS/L0sqeGM5958CRdhNjoIDZPZ4imPlm4kep+9wSeVIuaj91tChyg57zc2WG0ixvxlKJ
oZs1ZW64yZFjpq9TMQeFye4RDUqsazcwFl+UwqIDdFXxMM6iG61shSdVKsYiRWDctNfgeDzYBGgt
FCWXXafbJEBhnSxnLsR2gdBrFjLyuQ7X8kmpOryh6+exoRyaazzC9r/qh0p172dxU/vGDu9Tmxj2
zYQr9ieBr1agUOMQ5Yh4lzGFaD+wWciQNzi4XgGqezd8VYq4qEj9FmRoZNxsIUXA0g/4jATTfCyH
yc66a1ue0WUnuTpYeV6KlWoDxuF81KgxCC55IVN2b9TKD0oYWOKZ3W/m3IDiavzd9bsElMrg7YYu
RIFsR0Z79X1KKYUcQ+6CKy+7v0IgqFNnZbp9UlY6iuE1P5/VtGrGDTQZtK5IwGe3KZPTWhq8tX4O
AO2aoJNMr4f1GwbkOzv27xKQtncVCp2iyt16DTNmt535PpTh9J/oj8hSXycDpuhrCEd270ZiKQaC
8+79yDjO7rNjYfXY0a6sJOedBsi7D40yv6eWH4aBZ9UXws5bS6nZmWLHIwXdVvnJvKYnHI1fBAnd
0NQkisGo5hW1Ca2ww3eM1QwNWWj+Hnq9vFmj/h0NK+Od7651SoyQzR/pHXowGCOSXLdQFiQS1ViX
JtTsDMYIx8ilmQ6by0cOk3eF5ArOB9vnBEWg20q0/c5TUoqWVewlAVz9nJpVFYlce8+uorXYgECs
FkigMnlnsSwnw6F2vHuLdB8eiDS3mUOUpagICiCt7rZZW8AbXVvLYBUgbBBzxfwa2ELiS5fh/Sju
uzkVHKq+wQTypjhm9o8BX41liD8tb+Ga0cZF9uUzmByoxdmfwX5gkVsMKvo1YYis+sqFrDeOaBg6
hNsaKCvXSB/AmR9fFSfOkN6wI8D1SOmbcP55MOtU81S+zhePenirvvo+snydba5abiRA4GxuiaMg
Tjn+oH+q4BL1yzedNnfyfHZIwh6lOmnqtkCyc5y3/UZ4OKttShQ/Vs7gdpUQ4Z60ItE5zApkJyvo
tnj3zsj79yUSZOicajERm3YL4hIQqIbCAPKmRKBF8BnBfXlHZAvfZjeI93e7CeyNkHZpN2EaZLjF
h9IqR7aUFoNpXqfSh+uSvUZXqbXoy3O5JFvLDqHS/XdYsbiaYSLtDV9RFmK/T2qS/zP8qAGUKvsN
d45AeVZDryy0EFe4TGfmI5NegBaW/DBm7qWTHST85t58kT4Tk/StnL13f6FQYiXEmn9kVE22ySj9
7oQ/Ml/oFRduQ4lUBfVVFZW/MWJnzJHNlunnuGyx1RCg8Q2gQnCTbSVOSLVbBv6uW4K51Y9fVXMa
O2JgZEfhwRlOHUH+Czh4BEPDbhwUmM5U+WRVSK2PcK+ftEnTB3CS/R4YrkjjCOVSTK+ES4mnZC3K
GivFqjQSTinZEgIawFdI6vt+jGRCYeigWdhAA20yX95BrwDEo9A74C/2dEBe8nPduv+YWGl/k8w5
1UykObKApXs+YiM99CzMEjDRu1LA0WwTB6XqftQ9qWO1qHx5TsYnblRpIumSFCNO9QpuY2EviyAr
mJDFGkHzFN/isXTGDVuo5ITc0tC3BgPVB9B45QPJWE4a3LngSCvuvyFksvHj+aOr4r/LFRY//rnr
Lwh/l1FDbf7Udq1R9w+OLixY79QJJQ7bY1bE7dbE4NEmchnAnG7Ina1ty64kg7HPHevnOqBFb/M9
KGk4v1ca1DsIzGBPknkUHbqQF59f5znbDzDNj2uFenmy0u9n+WrQZhxm0x+VkpcG7th7+fB+5sRH
ir61ZM1+08kLg3IibFOcQyJstCmMJHm050vMrs1r+Rvilb8S+vao3Cxr1OQpfiOc0A8VOU9ZACzV
D/x0LN/ycvI6hWsETI1Ol4ZFaV5nNbL4stSIGK/NJppH6qBReHkKH7hLCPhGA99sX5GmzAg5W4zl
fXHW51faLzre7bSBB8CPZek0tipIi/zpA7daQNov8fn+Ojmr3IKmsimmyvNnr+rizhEzsNRcgauH
Ss4WdbLOY3jkBs5nwiHuFQNspAwOCSUXkRjsnfs0ZQR3gm74Va2AlxkHGpSkrJQ5jk6c0ftrZeuW
QgZlfuQunOLzVEqdBl5UsYl6E8KliPD23bGSn4URfNaHfd5WYur9fzMrzVkkpkctWere6g1Gv+bb
EMKThSG8wGgKrUZrlbEIj5QwEyXZqDXvgYBLLHIq9JXM7w6i3tRTIEs/5j4sqW0OVhWwI15U/5ur
HH437j32+3jr+GZmCtTD+e5UTWeyzSySZG0DeCsEAHw9dZkYhbq0tzVthh3JFcfyZTG5g30+L9AS
mK5iuQv5WnV5rygEIM2o7XY5CeqYzJIPov0fV0uAUmJ0bGWXQc7qqapzIF026l10LXKOTAd/Gc6s
bEYuZzYr1xcKTcaWUbwdX4wWoIPWiZx+oZzsB8xHHhHStUttT01ABX6xsOyRxQDrKPFgOTLR5U8r
X+aFbIAlC0KXxUPyRlp06VcjB2YZUVLD1Ku79LgijSRkmi292ZWUneIf07BXrDIA/E4P+rvdddx6
W2ym5rypr6O194lcd4gdEcR5KJcFqmQMSwjybHICMj8agii6Wo+MB67kaWFqYZyLXZCX2K4TuC23
ImSL1Y7AruglYS5mogwow2ceqaO8w4LoFNf8y7VFfnSZqtrYxTmG3Dlih7nfO3HiWWnGq9Lbom36
l0z8KAadOqAfWbNGnW7UVeFlJ2TNYtfU/ONJ7CAHOrOnhjXaJgNIfFxxTLqpMlLl/nGSlo9FpRe0
SnxQUx+s4u1XOp4NMT1RpXV3ayuT9E3FXR+u2m/gnV3Q2PtnyN03fRtvlOCCFZBxOF7YCSDNsOTC
bGMX3IsDYHzAx19WnX/Mdh/hRncRmeCp2ItqTRNCrcWBIWVzeNDX4o8SRm+OVJovzbL7dW9eiACc
+6v+OfMo3hg21x/sf55+EkEHfLxxX7qFYw/bpqTrk8h9du/v5/mi+ZUyNXFZOjgs/EsY27QLoypP
38EqWljSH0Ka3vx0liza9SKkgvCUnQK7rcxcOttVBBdHwLlIxNrWJ4O1gy7qBXiruSbJjZDGzLhi
hsCuGZ77oBGc/zM/lV797fWS38KOut8q9htn6bDMoZpjs3T2zM4kPtmLFtw87O+Eknj+h98tUyYk
LWAr22NMt5waOf6Lt0O9o/UY99LchakCi6s7Fi10jGX/wUYu/kZ8B6dq13GvReTHNEomenoX1sKz
j7TWDIPJYIKICJT+sKF2n4mYNF87nrRPiJxLdVSXhLP42hy4zHOpa92uvyfJeL7za71NFdg4uaIX
x8P9z1JLqnFSAfOQRlwbHByKu03N2vpaJzZN9wbG18vVi8tTHTVGWvFVsI2UCNPkGfsdLAO1hW96
kzJ4bqnzIJQzKJRUq36jxYrKpIlkMm8lxtsNE6X0lh9FcGYHFdqOkPC7SNPkDpHut+OIquzT9pCu
wstNTzaQbZx8iezQZNYsqFP7e22lHiyQgxj7KPl3swM1U2hXRCqdlgyUGMT5xiXNqE3vV827Rjmm
c+dlfYctEffYRdPuuELx1a2OT5lAgsNcH+ovOPBb/DYKd9SqIJLUE6Q0L8TkDl04Ua6hKG7X7hgc
QlhW4dktYZk/cfsa2gGYXfELYuUr3vUeTYzc+cEzN/oLhRCfTBKo2qhRuxaGozSzKGO2jBwcrqaW
7OfBZ8kY3eAv+4srlZdBpOYMF3JN22KtGBVPLVkNDwt9QoHX0JUnWVQ6FElVbbn5JE3PQrH4pMNG
e/Qn0+iJQLMpA0qBKocdoKOWTGIZPNfevfM5S7MDWjc7jxwdxUlX75IuvxCb0GU49dJDIn80HKPD
bcF0pZrl2aTa1y1RZVs9JFQIYsL2xisr1tZdkePadp1+S83442sBufPJrsHkB6GRu1WWrk0OtggW
yZfVvir/89szDfMFtEZUarq6I9O8ch6uuHIhNqXVGyu2tdhBvaMoH0IxHFjibSMLmMYU6gwAZrDF
u7p19sur3RIGvXvFcOZdWzaNEWct5a/chCY6apPJWvqPHJzsv23i7dgPfciOLKOl3HEAiPXGZ4ws
LcXh98b+KjSy6TweQnN0t9OI1gB6DXHdGw/3+bc8LYeeBC2Z/w14+jB+yX3NDQbCZmGqKjSvl4pH
kA7jfS3AX/ZJ/YAiBcRGqnqs7qptZ6NkxLC5LqLrAILiS3EYmaFE9zSr+Ql8zqCy7AUatm8Ideey
pYZ8h2kpnERtRN7UThcTWyzFWzZPn0V5F37sIy4XnIgxutncivUljcuc+z/gPG8nQvzAsRkTkwEj
IYjZKxYjOCApPBYlmicF2pB3w6YZyTKf6jUk6nJZlcuLRioRFxMD7h1+n3IxI7TVwyINHYR2Ex0d
RmpX2rB4JEN7IGOzZiPuNPLHRkAnr1AMzyDcNOwHE9LNENTUVXEO4Bvw/GLF9vXl54LeFtv8Ov81
d4pdJ/9CNicbyP/4JI8JVD4SPKBDrEq9TUTjoc2NEi4cItbvj/UWU/bOa42yq2vlc65LiWmNIyG4
8cHp76I3j38oji09OXuUVgnn1zjCOMvFywUHwFH7wFLuilLMZWHyrH2Qog21rcQ4bxB1NKYF53kM
B4jOgFUx9wTt/g/P5YnrJKNamxF7yCCSv4RnePcxGTOEI270i4a0Z3Pf9MtRzcMZ5WfO7ROA8/ml
W337/i+GviFLSSA5+goqQGYrtT/Gsi7Jfu0BlOZEXAan8V9vaxc7zy70jfCq44VNiNI3XkamX6JJ
QhQsFgV4iR93rVQWt/iY8cEEMuTFCd/JuDSvWRUd1OjXyS3jwuSpswlCN8drwasSFDyZebhB/y97
/z6krAz9gxCcgD3q9LKCoZLKovaJNgkhJ65eTBOY3Ehi3shx8+YmoKnQAKWrgdQSv0LP6kbyk8BI
d34HC9qtBp0NQcEvANYTwkDUUZ9WLSXfPi5OpzcQXR0TLZA+MlyDeaamKXMtf6wo2YPzEWSWcm0T
glNf4XDtU3PsheM+DopFP1oyYvyN0C7Jx5cZDJot+at40nbM0/0+MIUmp4awH+ktqE1owCVWyBR9
D0WdBvYW8W8jEDCoA+MsBffmdDP1LwWkRjf5OVDyfAVTvXk31E08Y6A5kvvjWoNC04yVsCp/nYuk
tV+dghRTYn7Z1jcbP9Fd1hp7FSy0fvZEl9RaUugkHFNiNcpYmndelnTO1wzJnjLcSZuKeq/NOblk
MU7LyeZhVjoDyLP9vQ8Zi5yot8rVvGfc2bmz4kJn1SvfNRpLu0F149NJsKHs9YQL6d3gYztoNtV2
qvbGbi/kq3WtmIoO8g9QL0ezK5+4rwaKYoNs3UfxUQX9qLGNnJw8Gghn3CY2i+5YXuKWNxfc2hoS
Klhu4Yqc1oeFJ38nnnQ2s7gUaDFlF51rVU1wM5WIIkEWvtvbAycP/nRaaZh4KBN1RvI2EV3w/bZi
TRmtBN4gmq+js/KfJTFzhT1dErQkP59CmDE+pIi19l3zjuLmA/xj/BBYWkR6SttVqj4njOUGQx/x
ErVOWW0STWhFWWZf5AuB7S2dRUjF7K7v4XGxwvsGYhVGll+H9VXumqCU+Zr3clh1B5pkTUGc3H+q
e8dzxWUHaorypHpY6HdewZk2kLMiKG6ThgVCRXCcg+fj9LspJTdTEk9kNJeGk0/Ukjagl1uG9WbF
/+8yga9CZwA1Zt3b8BHvG87S0OEZ6eOIoP++lPEKstk/3Qn50UspCKKkEX5M/3foj43GRSvqYDU9
vZxsQ3gABc5RIS5LW/Hg+XF8QBQqbC2YW8JFXxzYwtcrn+TkNZvnMPLlpS+oPDD61alH+uHe3uLL
xrh1zp01gEaubkLsNc2l/VnlEkOddL4eBvqZ0wF7IcYXGoP1jnI1keC+ejpD+Z3eDYyr80fvrIWz
gw7PAD5tr++UuMcqtnLQ7dzdu1L8rtb4tlPixExeO7Mn4Ckdnwncg3AuxZdAzQA+jzsUuaQmZeAp
scWy+PJmG785h5EI6jzAW0h5ko+Ssy/QKmGLBx6QL7wLpo1klKwKJaUhI7ePMcdIUuzB6smpB3XX
KbPAuwWgw6RY2rFOAfc++Fxp4+x+RvhdBSt+CvPoJUBnolDv7/vR6YngTR+b6zIqy/3rKeN1EXlo
FDrIwDkFBv1hypdCD09VUF9kOrZwlFtU9umLdo0+9dx41vjPA7W5xDlVuu6c2+tr01lgD7ijOwzq
2xoQ+lv8Y2XC6iza02uaIcP1qyfg9XNb5tbjkQoYSSAne/RipkhzgXKcry6LkuBz+IZQZv6pxuMR
U/fnkSo+zDX3nbouu3ZIkCVNpa9CgE5zY8Xs7gmH70gpurT4cz1h9HaGAr6C1sH7sfRC2IrifONL
51k5foABOIwNxzwj4qcaMHRg5mgHZ07tvn/nRGowL8YjQNbj0ZkER7tyYFOON4+vsQg2FQcXyaoF
TFLwZuMkcxthaz2TTATA/de0BNmgRA+jSoo6zFJc8nmYKR/WoH0pkhapjq+49+5/MRr1bDhU/Htr
yW30FDalLx3lYPuhfElIQLEptUz6HLSRBxANYswXo/zO/06dCQsSaJsm07ptuackEEBKClE2AF94
cBDH8YYhWw1URRjSf05hSGuPlOkeSnL+C1AbzsnW94XLpT0Uey8agUvxwoSUdY59YmHK4p8zDAD/
8j8ZSxkGEoap+n+VC9Kh/d4PejB9hY2CZMyR6A0VxMkUx4wXtufzLxuTLixbTCJvTKLxj75fVOUl
oY75Jnv4R97ntWULIoNFLgdyfLurPIOn05QTXF1x/sGrjba7qHd16qgWy3htRycB9fxvj+kvozAf
wcdg7GnFyb7p3s5aPyzNDPOZHvegGcSDc+89xbtSOxWKLhp4hOIBk8RYM5OXFdL2ncEnfaCpZ3Qb
3o7B2F+uY3UHrCaEDFQinmsPKXF8kBvmwFlSmGSJV3bQj4yWI0vCwLEIkerjrbO7IeUz4aq6OEcF
QvY0Yr9QZ1t0VljYCfENYZwRpf7pkJoCJyoe65INnfPDsOm5JwE6dWk4A+rM7xkaeKYtCmN6cvVD
FsSC10t8uHmckxMmfDAyPtO8yoVypRdppCezEwzMb2EIv62MiTjyxjQuGuNAwMSt7ku5kQY8tYZ7
WIoA6nI/qWO7JxpiJw8toFQh8eQuKWoYX31ty3RJoDvG7oLnh8EgdEBA+bXmn12ou7Giqa6hMq0K
oL2+h8yObz4MafEbq4Cr6K/86JZrnPgIKuJNC5/zuq2j1hHdXozArjLWcWtjLZ7tt4kOZCm3WIAo
gr34Gl1VVOWFvBvABkF8UIUQUgH8XfnJVbhhhBhlBazWRF4zWn9OwzeWlJTsQwC5E5xqzEzekypC
mUWTX7bXQPHdmD9TZ3pOOlZrrTDa9+Ad8EDYY6u4roCxkspKv5tvZq71jAacINqhhIiKhtkaAB91
4lE3tzkMGF3FCTG9FIR6Ogfe8NnLkQylv8OnKKK+Lbljv5P2V1PUHrWZOBWK2L5lTzO1GHPrTmC4
Xup4PahyMJjhDhFSIsG1d44iy0BtLRgQV4ZGtpz3xbwcDHlhMv31Qc6B+Leqcts1kn20WzooNo4G
w8pT8ISRDoEwtXtNbRkH6219HRX7ipw+APU8rCV0WyakySEJummVJNiPwcmghkd7NNLLVLz2Hs5/
MG1sItcJeQhzZc5FohQ0vNiD3+Zr5Ad1efQanqzSs2puh9SWpgopHpjsN6y+BAeIcZdnLgwWsPVh
RS7tO5BdMq4OTGnK5C5gXMyU3EClDYiMfFCVPQoGn3gN4w4wut1uZOJgMRBIkkEXJkkBmQyTc/Ku
Qf8BJCvBUJySdIJH6dAE15K+XBzg22ZBUQ/esspVpbbTH3SYvcjAz9K30ocCaDGMBmlCyhAAi/IH
dJqOZHbUbQz1Vjw/olwxqslCGGmIkbqd8is9t/Rz4tg3dbfAgqQ0zPbf40T+1oW7pIYG0ZWqFElc
PsvkKBw8PllMX5Wo/Pptz4H4f0S5Hjw5ALhNloMDYumXIOyzieCnlxQaoDYHlDzqi3+pFzKtRK3t
BUVuwm52Z6bo5vNmz5bhPWa/8uIWO+DLoby06ZpvhDiIHaNzsmJWwPISyc1dt6oGwRHn2Kxkqy5t
CGz9HP3MPyjOHPD3y0+ruVoMRS+whFD1i+LNJuYO41agExoNVFJKNVcFJ4VjbkJji4g70Xsz+LAH
fWFPbR55WZXmQ6s0hSg3idkRFZBcoIIEEbfM8QUXdwqMmSZYiMGTpUP2eiOgvL4HVdGod0F+/oQ/
vYBtMaBHctVEINova3ZCi/s69tMGaWXOa0YpaIJBVJKnHW6sbhtfd7kUkIJJVlL36x0s+XiMgvRZ
lh55dxDcZ62XgraXaF2vLV2h2UPFL0zd8Yab7dnctSlY+LJy6lB+a/RMP7+N3oL1V7BRWiKRkU1m
7NEwbALtwWKEjcgCazR9/Y9WCmLaRj0djCK85DPqlLH8r88dZxgxJNo6s8y/uci+j8hD5iSj6BdB
TZ0/F1SnrNngmDESKCqXBdPMK76sJYLvrEnmxrRQXxXsrMuQcKQMrhxNRnNUcycEs0WW0TsNvYDp
ThlUHE94WON0ri9cXDHH7YMuXnOGHRpu8Og7qpO5UTEeOey9h0ehjPvRxe+DhdpBkczJVf4JjWSH
lAghvA3yxKime1fb+Zk7Alwu0RsWRTaCqybZx/R6npU5mxgJQBGvwfdoFj6fx477niu43CCXqWFb
jihZkOfhSmb39xqI5hqe5iBSEFGCvA0NVfFJeVR1ClxecznMOw+N9eRwIPEJV9z3QX+w+i+bR58e
59TQXJu2Y1ksu1V8DnQbx3eY0gW+WAxg3mLfU7eyio8XTD+2FR3jXU74CbBhTLYok5pN76y3vKw8
uPVXxhGQlODrd+GxQaZRbGLnVhfF450Ux0q2gphUhifksA+LicwwmZjku4d2hi7bmTM8XwSBKhku
CVskGtQecv+12SyrA/YRSenAgPiBpmG1XCaGI6hCBC29XL7nnsEryXWlPsnj4vZ/13rD1hjEfdsq
zFLdJj0+FVZ5gfSSmdnzZ1ml+wm+wwCrHBfIAbzxcCzb0e3AlwCuRBsV7RmVvmM08gPjl+jMSXkg
9m5l6aEHFcMw9knCqOGJYWFaU4c0s4sRdTFhBv9BKnLCQq8uwzMj41Ru7OFSoVMdWq0N99xLWbjn
oKNj+z2uxhfBBIuI/mzeo4kORow7ZCD1MZWg6qW6HhOnxNIi1NGW+NClumNJzPjyGP/FOHG1izCA
NY5DSk+kMzWz1senyXonhnkd0gAJ7pzj1+BgtQfOKzZsYuc8iJxPGV2ffFSJrwNUybicC3IkOoeI
qMYit0k8as+g+WDCwR4ZDkLItoYDwlim+aDftSxCH4ImcVJUE+GKOm6+7nsH3gSADu99O+AcxnZn
evKfWRWO8oN09WzJhNXlzktNlKB2wSi2xrxLlKKVTznXtSBQ+FW/sm6+B9aFWjzFwpT1gKgtzi1Z
YrQKSIM0MJ+ase0QbpQ3WNLXWwGilrk8BHSYVBZVGtM30aWHhP4jlzobTgX6QdFOxUjm26Px5epV
WupDWSFkkoB/omXdH1DcqHtdtt0370opg4UPEIuyNBaCrtxnYjFc2m+b7Ams06hUXpWUkHNb66wi
A6lSyf9CDX7BfNOp4poKdWrhdD4/VyL9dUnL6QDqlylr+uZbPoT6uq8sJWheTDYCDI+SlG/4MDwb
pYbvcbK5r2LOC2h2ROtflwbFarZwsqsryjLzbuiFEx/LROKRTk/ZfFavLX7xgYqWGeCDMPuznD03
r6pv00O8fTgpTwmo/FVXHa1OG8cgavGnySniHqNWZD+KxIALahHyMUPxcW8pb1X83Aeji+AB4Spu
DflVsbvH35hhljMBxpIZr4Ds752VN1bijM5oC42maPuv6CnXSK4ODVkXBZMFzYYJPPkzMpB1NM5P
l7SJEnlG/AUNd9fhS/eYA7y/RqlAIkmqfGaGSYHniREx4arnD4Efta4gvIJTNiEa0VJqWjwEfO23
dr3BcZNyZwV4dRF4jHauf1v67V5FwEBWfvQv+Nhqvlq4YwjlevkJfj0E2reOX1adrr+8X7r9sayu
H6TWUEr1Zte/TrCcKSVpbyPMHJssNGTBfjoBAPlEFajTnTOK+EyKTtnE2a9z5E2xi5iae++3o5e5
XO2hMboErPrrvxsmETHsscbmd6JmZ1nQao1sJyUgi6hKq7efONuP1CkYJ9moGNG8EcMjf9P5pKH/
KfdPJjKr6UJ0JMiRcnHF/WvFMp33iqouxDnmKq1oRN0w9+SS4+O1+XvqULX30Xjf31jxTsO3Gifd
vTa6LKxmSKT+nWH4ZHmmxoAnX9KQxCdgAhqe3rTYyAyKtvMXBnsIMU+fvSFCvOOd1xMN/LM0B2Tu
uQYr39WeqiRiMoWtFgDTwTOQFZHAfEIS1ahLcCYa47JA40pfAaxfmEjhmHH7KhholfmwO09iACP/
NhzrbxUnmhfSEtocsclPrw7uReZObEQ5gd+daYzmYWOLRv/kdZUBLqUt9IwhzKVG/TuiU/LGhIAg
HoS/A0NJLIGmUHgeQqioF3qTPvT4CctL4tKQ+aUIr3nHwhFNL0zKCh13qxk+b/WOkTyVYZthKovf
WdYYsGP73HKjaHkRdLizn3MlEds1qPl+RM+nkUUBIxcsjy9HFLeXTW+g7c+bFTvb0kNre4G4s3L+
dy7DHuSgHwVr6hO87kuXwO3ze8mTYF/JEW/NG4oeFD1jEHWuWJQqCG15LEiPUD814QSIbkI5cBv5
yEq2D8VIzdg1h8zgb4MLnM+qbnEFkbN0TbEQhVS+Z4U9tSZgEMqSFnC5TI362fszi8PACEGsspHE
Aad6MdvGdtnuXEWBwysNUKZotfTTdeDCAaNa5FXZVjOvn0GQsQj4kGLTGfsrLAup+N2UWO4bJQFM
mjEOtWk8pHNbCbHohKm0MWGjtcThCbn7KmmrEsFXpgCuU7XwOClim5wbIE8xFHNGO++GqX2TXFHM
MDetMo5rI64+1bj95ISXMZuaLywzJu6F5qFmKCtgbYybHXLtwxBfIC0a96WcOvgym2nMKpJOjMsC
wtxOyC4Fu7CDRmw242QAbn3retLZ78qN7+a9PG49zCBOc/dBJRutYhAcqTBSoLzSyTraHVYRvv1j
aG7k5GYi9S+6kb4qsKFk5247m9ZmXD9zjdjqjnQSTh63smWe2zyyO3qqJ6TExEmjDYvRDDSrk3q5
OtW+FGQzqNWfuxNAvXAbB37v/ySCp6Mk4uXsti7nR7ugOlpE5AUcDWdXajYM7HkJQByjaMhvthSd
9Am6qB2z+pUMeF3iRUANVuBdrxpMlGRPZ4SB1R/MsZOHty2cMSaKKRHLtjN0N4no9wLkzYihldXE
F1D7c7jDieimg/V3CUa7pXHsQ3UEPCuYS5PDHwAJB7NJkNbGcjQABrMGs9W2yf+l5OeNmMIWU4HI
uURrXzHbEJcdb/YxKuN/oOdi2dVjOTjmcILZAxGS17yl4HMjWP/cJ9sFFmFTWjengmaneM+dfnz3
YomFIWAhidtz8aNIQGeJFeSBZm8CnAa43q8+yOTA1Ei2f4NnTLCfmJi+XC9Alir9tDd8iy+L5x3Z
DFq1xpkiTIYhPNP8wBoJqHjpWRU2MY8SLuVHM1MGnl238zMVOBvbmbI7Niuv6YwKIc8iQGyInfp3
YHIcJsDxw8I9PorM8WcepgyckHIN8yzNb5FAagH6e8ZnD8A4kVagMVsSG4y5CA/Wp9Rik+KOUlCj
ur78niDm4YiBec77NqTizd+ygRmmvaNBn7Lla6ASUJDnUFEjkpBa+j4m3x2Ip1JW18CqzBzlsfVS
hPkSfMdX3EJ/eLyAMSfqzLIiRvGEJKvKdyj1EjIgwoezXDu+VbLuMsx20xUI/IsI08jkxOJRdrKz
DZUjDKGINRbWto44KskurgI/5CLho3JZUtKR2wSu0JWIIhDyb6thkXuun8TkQ6FtahpsnxUKi/gA
87w+gQEdJ570YMf0ELg7due3Xat52+CKeUlAyAvlsU12b1fbZTIru5L1GJJc0oSvM3j9Wrhmxq8p
VuDY/1MdOxT9XGGYBXwBLQkeexMeTO4lHI3H765Zhilnt4ND4VfCR5FlQ1MRVxgyT+qyEzQGW6Zs
t2W4fFJZBl8tOtltdAfn6nceXs1lgx8rJ2zIkxud43mH5b1R2qjb75o+a5nsQnhHKskixIcRPfd7
4fAPRPQ25zGrhEvcvqVFio9gxUCQtJD+mFzScNOhM/kBhkdfDTtDVMbUW+mcPi7ItSEIGWU88cZX
Jqe+5lv0P3ClDkNMMg4QDQ8une3T+HCgiAXVvQfc7Y/ASE4ay1nMDinRfW9nGAiGda87fG68HLBv
XF/fjumgeoR8T613wX6BLh5+ySKtZRU1phzZcqJ8Trui0YYO40ha52NF5o2M0IWU8UuGvQnHNNtC
rfNNB/8vwdk+60QTdA9FzztUFsvJOYbp5DDViHFrAO1O6wC86F3qITWCFdvvKPx3HNfUFdpO2an+
t+ZJZnxfXWxLpfOMLz9bzIz4qoabUEO7ZCKa8+/OLr/VWqZ4MCZ4mEtMuZ7c6aA9jvrYQ6JSGFyx
P8IAmUot23ZXUHCl0A79puSJwoj58JFXMwsQl+ONX6rJquPdlKPBGqM020R0TqykbxaOMCkbBrDE
doxGX7Q5btcHDG3zJgEJN5XSqdz3e+WfVxJMZwpbJKhfrkR/hqO1jtQpaFRa5Jn/h2XS83lphEJq
KlKZuZ7NnqZdDTC+ObxqTdjELUWLFiXmtYiODL6Lz+SH/LLo9DMzr0S+Ss4ImzGK1qTigT6jb6Bn
RHmxeZh/9qbX+PAsdu6zF1uWjzm1sGgaVRye6kYsc3oEbdO17A39OjHr0Q56fzAA3IW386L+1beh
yyfQMuxxJu1Yy1MDy3S/gObve7bH/Ow49RrJLdkMHISy0GjlkIJ6IBDTuLwPoxr94XnEXS31zGQo
0dXitRN22FfGUHOU3KZuIiUoCoNuLnpFojOcffgg6tq5WsmQNRxJiM1iavW2oSmLba3ltBc/JKKh
bWiIaly17uOEH9DA0wdXz2J4dklbjO2PsXebCtUYdM+7uxuoeT9/lHC+tS0wJykSFcWX+GKLO4ma
nmCjE0WaCEGUaghpbkHtKSwYcAaAHk6cBrgGwD4uBt7tBuOpr9HdH9O4u4oMjP3/2ukqkP2R/+Bn
7F98VxzISmr13czFP/02t4c8kFnWnmKmqQwMzzNq6h6+jCBB+0Q5oLjoAJjwp9Y+TFbzL5GV/ArZ
/Vv2Sd0hzNiEsprgqs5WciNaj5x2JvBh1Xt1Tj3JDNpNW9vCa4mQ9BUr2NiqGcZkNLzuzwSymNJ5
E7JNL88UaiOeTVk/pIsgbLYdJE1HgZO36pSFsqN1pDulE4D+gL89nF3OuN7mIuYGr8QR/DSvBrzG
yp9ZyqyFVyOSb1JpmW2MdItfmFPoF2JJliVQoO2TJ9mvX77DicPF/a4pI4gkRsPMJBB+R+FwHxou
Kz7cICMJDYnAUxAJ7s1ytwuTzqkGxGxTXhynlqJkPwiIrBOTnHeUb+tODaooImLmz614ma8q92ne
if+2chXVw78DvwvxrXTdCN65ZNQnABIoZCS2zagwfrfXd8SDlcFukGxJ8KN0gWJkCBN5/ad2rVyX
mzh2zek5Iej4TDLIdEbgCLFllcvL+OruTaytCdRzdpPycQ/Enr5jeHVO+UfpzYQIVNCGK0Bt6UGS
29665GUVdRwbJwBUwzBwNy0hgt6bFq0VSaJVEp26HZBlh0bFnvSHdPPI3r9ETCUNOtLpN20hujDF
45vFAq1whwHqau1cK9rv70QiKk7SgTGrrxKoLX9Gh435Cw5euWLL8K3GRuYNND56JNqJxvyPfaft
vfSs6N/S4c8e9F4z1jax9RnNcqB+Z0Hdua2uB23mCrGEaaETr7Dtnk3hVwlwOAAxKKaXN4OUtOtV
vge03AdH/Z3I9yQTSiTZ4fUPVPO2ENVr7tkCG9ftQ/lE66cfX6uJeyq06UWTGtwXcSALzGaM8Q6w
6nSWlhdqtWWAzb10GTma05lohT+eFuUNW1r6RVN7ekrjQuzFSVTvKGDgsiQKUCr55kaKBYPn16EG
TB/jOCQNjr8Gxt02CbhemV+AgOpYrY3YNUe4k4JJqczfXsCuhLt+BQBT0DKqcFVyicY5UD4zPB/b
GrBFQGpyp1qir0KDLEnGY9vapTitGiPioBKh42yvGy8JSh6X0gWblmzLhZ+P3X3qi/DiddsM0zlZ
fAShgoIC+os5i/1lOv6ttAfanfxNNHmGkLXb0HRSLbmEdnEjhi7SF/g2RgI98WrQmUrRQpJS+JaZ
gxsICZOYoN0h37VX+Yd0XWoJNEKZeAh33Zz/WsZOSRaEHDVa/x7TSqE2Rml+6Xi2iiGgKaiop+Ir
rrS++a7nZjBqS4PL/qh1grmEe96rb0XUvFNLSPRBptIC5Hr34sbjO93bDeYuRO6gbwgmWBe0d3SQ
PG523nxUabETStB2H6IoR5DzKMPh2cVc4TlxUBjNF4Af/2QcsgHXKirK1nhf4kPNXSxJtoOjsp6Q
t+u5skfX9U/Iv8uGuU2eDtbPwIK5wMRcYuKEGrWI/jFy7NJQE3EaOBLYfwj4TsqIOejelJgQv4Ax
rOu56QucFmjkWv8pxOqirg6nqg3k6Eam3DnAzGEpc2npmNM1lrYZguVJrwNbJ2kP7ESXj/Dda4Pu
iEg8PtEIeZha1C0GtGIgZGE5MfAuh4aRjspqhDKy0sEGv7JBbuJxpkd0HF/45cXdUXpzfOUy5pKP
a7Uped4fRJiIMX2FNiJaamana9RRJ4xBy6JlUvcWbSSLYW8cMy4BQs8VwsSq0mR/IImahi3uWmeU
W86t7tuDFXnvZcAf1TbY7fzBNZlNfYdVLqMeLNeyFs0IQao+gAzKF9RgIrsYzYKOnnhNbkkC53Fo
jcQEER8e8tAdKIuTujsZby0iBncEImitWbPZF7lkoOc6rM+HPb6riXpm+WE/UJqW2B1+a0AXXFvA
eLamZUh4CxLE06tnueGPwdGiTNPeg7M6vJSGj03NRAcMf7rgQGMdX2s1/3Phu/84DzEkCULONDeo
gs4MzEgV/tPK8m8E9ZZ5aFD+fz2lRPH9gr1aQxrJOey6qZmw473lMTv7uJyX0IOLc0fjl3G7DuY0
NDOlJG7HEa72/q7kFsK7DJLevW7rYw0GgVgWJHLMy544c7niku7LLBSXqWyaklaqArz3aDyzgoEx
Riy32HlDjf3fqsL9EUepX9w8WOUlbfgcZHI6zdPKFBt+NnKKCamXrYmrQ94UE5uzQ9LoXYSOZ+Sx
U1XT5jx3AEJztNHuZ24gDiyE+BfHWMQy3NgU02hvWQdqiiinIbKhljPgXCu0BI+ebElCUNuWk1OB
Y/UA3rgexCBgggjSAGTcX04Nz4HMu2h643BL7P3BYxZL+6pk9W6MsJ4ULrvsJk3av+Sy3EVY2X8y
Ep8fQVAAI8SkvEtPrgdqSuXc9EfiXKVd9QX+enxBotv2xZQkugMtF6LdCL5ahi6tQLNayxl3xpvM
LzMAzXEj65t/NfisDsXE1YHlcEW7HbSWBkNl+LKNVszrd2hDqmacnebxbgrd4AjZIPg3/eMWIGNd
X7x8bnYKTLbnXFZyws9LtbpJMSyUHM27KTH+vyLdEZFzrVMKCajGfULwtps+vbzDgWa5wzDgROaF
3KQogeSFllUR7SRd0tHzmPDZPvio14qleePPJ+xNHfVU34yKvhPOmgg37MP+3wz4lp6Q1lA2t59C
OExshSrrAwH1gBbv0IfcA8HxoHp8jffnN3UjhvfZGWW1usRfNVunZup4T9yZievOMhn5H56Ri/ZB
hZ56fzoIleZc1hUu1RpTIbWkHAaDHpu/cc9rScdd9Dr8L5UbYaxU/LwMhEUkWWK8jw1GH992dYvk
XF2efsFyc1KqQnwpffBTES4FUoAcDMHzc9i8DIBPcKeqwdMX9ERxpA/SC6XKLn/jqJYvH6OnXsgS
tNUKlvg0lC3qXzklx9uT5pjzSBF1omGNmvkIHYFYyANqKOdxnBdv/BgtkTUuI8O2d0gxJ02zXHQY
OLUTDE88+5ayzW3Cyfn+XcXXlpKi/oU11D0m6hmQcYzuQfL1IEfk+KuMrxx3otNWG1HGt95AXH9h
gr/SyssLjja9HnyELygCKA3Yib7cjnwsdtnJKpoHDkf914NEUhUblZqMRCkQcWbZve+UZ5GfdiL7
2JirsEYEZ2/ufWGDIy523MwJ2qxP+fMzAlNC/MeRKvKBeejJRqofuasfRMYj9m/5vwaLdOFr9C6c
bXKoTchp/oqvp2/Jr3H/1fPCwINxhYvA/6KX80a5CUTEK2ou8Ebpx24BFs6ZplJYx4RqOCB/3ljT
aM/7WhCNNFSPC3J4uuBY9sQ+o3+o23qkOluN7nAym3h2QrvoAcsn0SRX/mhLKv/UOFeW3wZiANZr
LsbkfmAqpNP7wsaGdPxlvOheiZCE7xw0FRlQpW/Cte2l9B56eBM6zmyfiGoZ1VXk2pGAHzdsVc6q
FR8DvN/cPscOgsVhS+tgU4dEKYl0g6IqDZMLy0TO5doR+YfWO60RCoutep6AfMqmnUptYd1BDwlF
Y9WB6EMKRear5oDLfme8T3is1w7rcJXG7ypSMMwtrVjCFqcGYs2iKiH374iEHmJGQJYOP4Z48uBj
lrMJ9+BKPgUgwX682G8X3CRQx1aK6yf5SEMDvIakxFrVBtzIJJDQPUxKo+TjlqAOwBFXm7NF+P2S
Bu4kkWnG2T6Vye6gz/B5nJ7Vc1n/lXgeW7FU+kbLatmI440STzSwr8eh93hQXWOhoCwCFxszI96s
mS0nl8WqNCDtNoZUioyRD4bqWGydT923e1ugYcNRss5QnK9s26Ym7eqqosWKNfGo/A6ryPgoDY2K
gU5z9kQ0m3IsqMWWNMKtGI1w/tzfmVg6XKg+QXuV9Z/uDGpDvFjmpsSlLOhvyM2kYSilNd0eiMPL
hYvOhkMcZOHndr6QSqwS4W7rHiVMkcaf3k4QBQRAyIsOvH5hCTkE2pHCWE9QymNq20vYEjTcalFP
jCxtj1FsB3DC5wqHkVQarPGC+rdcpsOj7llt5inhjHoq7Ggnem/A+zONbtSSFChxYxM2c1QNgtKB
he794gM+6qm747e77GWhbSXVCJYMA5aImpXNXrEL8/4FSNbu8yAHfSOr81puJMUmllgLnmNg9+aI
TCnozjpseUumAUJDQpYJaLnYjWbHfIU/SQ/CKBR+mZupWgtJVp2ePAdpXV62pNsT1eUY2nc6xMip
XH3zk2IPzCxLju+000EKpRuP6jCwY3LoIyRYCJv6upRDEddF+XpmLPXP8fByHr/kkq/51O48/Sho
ZEYRJahtSBdsfAyxZFWi8h6XmgotMdTEJT1KdyLhKKbOT9ugusBjmWUrKFcDHLMzpHX1ojRTbg3r
3bx5VmhcmWqaFIRK6TqyuBAbJTlnxscd61Tb3w+hR8yceIw8tlYHPvkutU0H4kHo7qkf/tnvYpMH
vKXHvbyLcXm2O01NAvUH4emG+JiFfmF6TwWr0i1BgRWc12RioRHcPlQZVFrUf+3mdKUj3vqzmaZ8
vaOQr8eIeF6siQ30FOrl4VLq/y29r6BwHgjRypvi/OJkXdgh6qrewqe68uydHodbfG0tpMoZC7WR
95K9g0cm2cfA2ihjK99DXquIPkp5jSjQ83L0gFOLAbL69/tnfhbdAmYuWRRCYMc4pDV/OO6qQBFH
fhgMh/+qI6GrgPmfHTOkJ4Lv1F5lvHxcRaVEGwAyfGGBOrrRjaJzEV1AswkHmFPADEtaDFIPuP3C
R7wgkf5tsM2WsimRuyUPrDc+1YU8FyBgwml0GvLPNGYAb97+is8eLjx1u1vD5UVUe7vd+465YL7u
geYLLtSBsntLYYHg3Q5zAbDRekLke/DYC2K4IXvpsnTojUwHF1HFU7fdFITorWvLji/Fb1yAsuGF
HYxxhlribjfQFjt//BPr8944EnJMYLmXa91VIQOZcVafAXwK18RuHhW4UzEQ/28lc42SkeCTB0+Q
x+YIWfLEYZKf53dAnW0EObPbyuaLYjtQ0ZJc6KGWcQftSoFX8dCCSTSSS4NwnwCXp+AufBusoavy
68e87eiQa8inzKd0ifxA7bJbWTYsU0uOYd0N4Tx7flJx4iG1l0L+xzK1InlEEUom7OJ69cHSzKmk
4PmzBzO3Kl/ftPEelcLos/KbzvQ5WNUxgBHJHONLYDDuPcWMTz8ZY2ssppQsmjBeMO0IW5RsIf25
vJk8TBAlQBboq8URyglv7pOFUDfqM7V3ZIXbZOq+XUyslAPT466y5B+HC1zi591ksC+ERK1su/az
8WRR9fCbrIMP8nGuQwypnsGf1DDRuHZkeHuXgkFMJhmSd39B51TISPozmrZAWc4PJinj1fZjjs5a
jrnHJEO4lU+DRfcOOdIoCezMSWQaIEOokr+C7k8hU9TdNNuqwJgLbxWupi1IbZhgxp928lKUdJPB
GG0RR5WcBFL0RjVvd8M4KrToxx5kXSNrZ6dvCqkEOttM7/mC2LfjY9kx1CxRPf8neSqmHN2XQiVu
WHNq34LOHY0IU0U7cai2NzwnsNlOpE7RhXpjvA2jdcI1mPhZifI3lvzZrKkO6HbImcgxBoOrRhZm
byH0Jh6emFZk48GoLl6rjTBIOGMin4HNUMDiJs77DgaxVUbk3K3zqphW2Q9utB4NdVUtAdJLXopl
A37OtN+vnFUxacWv6OpN1cQpDt6a6f3W7x6CmwOvqfs262ri5FXQsHbPanPE+MbVPg4yk6tn2HHU
975eICCqgGS0jb8bC5VY9fRo3M+D7yWaJfAi+fQiBVIL9OmM16ix8v04CVTfH2ocT6gR268NWUl1
Xzv2BzReifGW05OZiMIFgKUGNfzBXvwJUjuZfni6mS8aSQcUNfUoMI8++NYFMoMWemKE3CWBQnH/
tJpcTwNbWXBK2X4VM4PwX1WOSBw4aNA/jxVfKu15USOMXyfQRyVZN61Xz7HvlhSXJ0sNelPQ+M+V
6wMda0uf6Fwe9Z0rFeeIZi+EWS2uDNE8qUk7cKGSiiYvCvNZ6zpedRPBsSHDLEaMShTbkQz1BTW+
ps1bwuTsQvaOynxOEIN6Ha5vhdLDZ6mK59ivmMiNGFQtxkfaUa9nQKPQW8SRvDkzNdIkMf6TceU8
0f0j4LU8Mttp/HCtaNm5bT/zDnZMMJ1A2jcFDWjihIENrTErfYSMGfNkQ/QgNGWH7SqNAE56vc7k
BAldhvdPXzSeA/wz/GlFmFFhuImIdypkU6eKXwi8BUL3OrFPS0Ldr6YZmdDD/VTjsCBfSEKmlM/Y
Load3wzcmoA5VRQ98NNRaJzQKh5dLlfBY8MVjR455SeREOo6ukDf9/JJcOePmtnYX8uK7db+0NZk
OA+Lf+0EX+5GuaOtsvxnc9RMnxfLYjfC/37kNY/akzjZQdWPBNx8mfd/0Ex/6EK4jmSwnnJo1XL6
H35DEGE6eXPivgblglO0YgPunFBjWrAbJoYhFzLDTIEblfgSQXMzrNL3snhwNPhQeY2ZAgKkozgc
z0UmNFn6G0wO3sGJ8ZpgrIXOTMWJ3FTLZG0lxI65QJSyHd9B0HUkOdRPLf2Oj/wHI5SOEeS5nmer
usyNgj6vPRhXLv4kpSpRHPtjw4stEHWCTyM3GHrtzVQJXPybDCLM7EtnQdcDt3hn4pNDdIwwa+o9
zubEKziIiBkgWYwAtaxq5qMWdsxNgXxDuTiLTHD1ReAK/xZ4AjnT1oTK3QZdlAwUa9ykup/K154E
pekw1LiBGFXS8uXkyf8RCBfs/oOsbkzZs3KJAhBByNJrupxq0KNN3IoSjIRzMSBjYydcyp8MUvL2
cR2pRAOp0zA3jrhWh/m0GxNZXAzueseUIB/SIJKYXVb1T6Glic2LqXf11/lU2esiIsiwLNE4/H/w
94qkGIpgqEgz481NeRWODzaA/MzdPe9Zp7hEATnM0iBGDTofLlwuNObs0gWk9PJCLMxZ5tU2KRJ1
Va3fhWTYDX/GltkomYmG8dBA+FQ4BVaPtLS7fP8pJhJihmLaFS+XkU4xB+SzqDIvzPAp9gfPESXQ
jrxsVKtnAQkkPDndrAOtu33pj++eazxoHMsnLHz2enpSp0KhnhaeOnbmvBc28KRYy1u7uvTD0eKQ
dxmQxNqQd31rv1Nck4nn7zia5mc8EKonN6qKfv1jwmeXRhI5wH+khw2u7ehEnP/siK6Aip8EEw2j
AJOob9YMILuH/I76eMzFCE1dWPsn19fJ9Rj3Mh6CUItAxJcEY18aW9lidEfwKkhtUMsPflWZYPoU
Ek4It9X7u45xLqOsVu3PsIQunVNJPX6fc/23/kqanTRNa5MTaIm8cLdQNkJTnI0BrNeCjKbRBa2v
zhi1eyhJUaBg+NvDU3XH5BWlqP4Sqr8wACbAncEtoWgarq0UXDN6obRna1GrjzxVS6xobiLS5iEn
kgzHyfA7zm63IXL7fxK4AUC+3nX1JR4JPSkWEwLOTZiXBRo2nh9EJpJcAx32ooEpt9DEty0FP1Mg
THgEEe3EPRTP8rv0v0CHi38DJ54TV211Y0jMy7DflQIkVueHEdZ3aIKI6fRDS8uYtVHS3gR2/zJT
qnW4LHVYnVplKgDSJB2E644apgr8UmU0qDG/8xz+Gpvw9EPDJgpuUkVYyb8e8+1PIgROn3eeIM+i
/ljiqMyc/hFUGD/r0Rdg1J+9I7kcTeGzjrnMUHShnqN+vE287reUoxjZZUchu8kq7RVJB5SlfpFM
wnbr4RVg50Hq6q+YlF9STJd8BKux8NN7j+GOMqoPFJRwZ6/X9V6gBKOrURegqYk9weuHPbGHHLlm
S0Sg57BtX4WuR5bdI59gC17AcRtwrST9YucEngnn2im2Fb8K0SDHKfQFG6rpP8v/SoXysO2JoCH+
ihJTXy8PKJBEgp9jLabFg9bYzajr1k5VaFOnLglTZZ+aCKZANOEf6kt6Hb0kvHEd6Sv/Gr+YgD+4
qMlbAEMDh2Yvk6YYLlODenD85/DcZRpRfvwk6CDp1xzFspnqB7k2e+taN3BgIrEIrxPZKi6ePfu/
VgCcmgbDcIZa8q8AUFyWaJYkWZG+4kGT5PTArzlEepDU44YxEwME9VL4nv+B/T83pb8lHe8hDpw7
3j18mCicNqjdqz4x7hdYm89/lYRx/LnMtExiGqAi9lWKeTNVgbuWtoRi25YCCusGa6sdyXNCvzBx
alnl63i6M48oaOemmFZLVOTWYADSRVcEEkZXBigFe4e0CYOmMEZXSjWMQlUh6MlkQsCP6EE1UwHH
zuM6BQMSIN1NQ3wN1jvq+ExVRQynOZ/FXgYXzW4dMjqezRvezLGe29tit3+yfnsAAKRcr6WdgIpm
jTYxMuzve80PD8y865zcvmNRiHslH2vIuxy1BL8sIFuID0qkOmZ2iEA6XwNs5WMTI/KJkZsbfI9d
f6rSJ7on3OxkmF1a281CNONKaEAC9i3H98HYU934lYsYjn9UJ+MP1SU2sPUyDdMRlrw4h+P7AhtB
vO0OkNEiY10ENtJJQM9nBwFH2ojW3GqZi78EcRU2j515Wz70/YCtC4nrPcbhrMfxs1uA90XUh8nn
lOrrnG+FQcUv+hOUGpGbrWo24Sayvdwujw+9/p7qzVQLkuCydm0uN/lBzFxEk0E/DkB0s87rCrW4
HLMY+iSpeQaYcfJjpfgCygtrgOtEhXWZ08Ee0DSLqD7B82zAOV0WZE5H4gIGbhNY4WQHeDyBDqCH
6MzaFWsxNlstRn0sAd6XT2nsoABduuO8NFzUJfab8a5YeOeEBhj3uoaO4cUebzNV5zsYpxigBfXz
fU3IgX/Z7DFa4ylD5qroHjstbxQKPmlmxmJskZWPb0QLB+ypOcVEvh5GMiX4DZpV/WzUfEojLVyw
OzqQyNWbzJg1cPXSPGdC+jPs5MkuO14Ei6rMQo6zcqtNVsCdgU/wzZ/LfFmkBinlahWkpkLxzZaN
0UAh8VLWb63TXTPq1yq4O99YhppwXRpUeiQsO4oyMjQ9PHkpSarZMSARZpvRaDvqJg3rOzrlctaY
xh/rAYamO2RnFsNX/1NLATJOvbxKQgDOOyVINzzR5FORunKEWIED3jHU0M6dml8glCq76jKz7Xio
8rxyOCaJSQgZ14W7GNs0Or8mtlvJj8yadmvPMuSksJFh99kj/7WTyx5vF9m6PYmfJNMlGl6Z0Njk
fut9HBX4/NLEaavUjY8KT3xuPidC2KP+jYH48balteIzadIoD8PaAl7lT+PKxP/B7XA86T7G5xOZ
aHvsjZ1ta4fEugNdHecnxwpoxe9N9N9Swfs3M22ZFitzxV+dhrPwqDZVbbeTZGfE3strlyCo+1Pd
Ljs79AlPO3sztPVOX+BlUCO2G7kSmY2xZBDZFVTCsD+PWXGG3uhMKUPoeYbPhb7SbJ5kD6Ndaisv
DVfvD+OzYuUmVSPxNav5qMiaVb1XoX9Zs7G7LUEGegwPHXsR/eNMjMsg3Rt0+AdUdgnfNd/1c/45
t2Vizhkxue+NwEInfnxgozCK4FHltAEFuOmQ0JMKOtyCZFk9wbOHVVqdLtXkCZKPIyZ/yPxQd47h
BIUtjtPFEIPx8cBj/EK7yDgNjiDBWrFS0mAwXAWLlHR4BZQlvVBV7Fr5lQYFv/vdiS0zVeLQ/Ail
TSlhvfEFEnLz+S2ChbI7Mjx+g4Y/1KpRBeHLyfh+KDZBD/ce8jkicfxFaNUwxm1Y+s2NW5BqaS7J
dkU6cg6zKyr4nuYCskXaC3h0n5UyFe5T3CT440gEgYo+qdnFOvOCMR4sKUQ22ni4/yfxB+8490rT
2nVSuxUtw1o4zNaf8VEDoLLaFmEbW8464o0iVj+j49gSNfYPshAsF6rjg8OkjT1QzG6b0/L9MHAO
BdTMMFQCFqPsJv0OVMLMwbvutuXefbFCudq0GRhdPrDV1n4UWs4v9QeNk1zSXT+HoAShzNAmSRc8
h42Xt3HjlznXqjUdqnWRktT9GYy2AnmPFJQFfZ552S8Cy+XOB9fyW+iJmozwvlx/+NhAELcuf1EW
KVtz2IbDALQptubExjX4HAVBLAtdDsuD90Dxtv+RNtwkgn5K6vRwIwswnE5ENy2vg6Gv2EhDtTJ2
/EKzf2M4qThCutrfgNWic1QxGRVnSi6q3mghO1DvmJBWDFm3B237/aOFF23RICen5S8/CXYNcpfO
0IevU/5PQCh0tYIfx+mm3CwfWfdZMyAnYWLPpN8OwTvq0lyJ6WMBenJayBf50I27ZnXzJcWKR+U8
TDlfqLYk/7zEZKowFgegQNd4PwDVeOKwgq33WZs8BRezByDXmHbs3imdCi2+ciU164uElsyBV5Fz
l0pd+I4eXj7B3Eh7IYczbNaqTqs50cQvE5qm3YuH3Zn9aD8eW+XurAgWuTc7xKrR6zpeBhKskdzr
jAUKpoaXqFXujHuz6ljechsrv15Tu9aO4Y82yW5RT336P8HmtEO/K1XH2a1gNiEPQd7n+Gor63s5
4H4GPjKKc6hbRDjZ8IdJ6Y1fx9PZQ2Tw1aLDjtOvIc2f4IpvEKdgVj7QBJ4wlBv8ZkFEWHQws0Ng
RUCViGThAR20pmV2UYP9y85pW/wgmj48yM90+maMm+xF4gBqIUsyGm3WA6GHE/+ejZUTLiXw6356
FMq+zrydt/dsUCyr512cXoSTJM5hEHJrG1inFkJ9mOlfteJjG3Hu/o+7KIBkSrv79PINzTkpWVd/
YoViIqghUqI3sL2sUKW+0QEEq41mAcryE7U1smxjyHUQGhWUyJKAFI7V7SwV8D1Ok30PyJUzZrjO
FM2oH4sP6IUuQeqK5+t+MxC2QXPR5HB/MEES0c1kriLjurYgHpwmwCRLfLo1WBhzJmTxZyfQaldw
YnP+er7A2x41769wjtmgxTGJIt1PDEJkiJErsThg006831NXMDPGQJBr3V+SBrZy3Wo7v7RZbbVM
Fm74/J3/USgR4JTi30ctM/CkiiHbtxhjjyOPG6WlqjtenpBe9JJs1SbtHuLfZuhIjRox5wK5HqKp
Kjzlq2wv4+EUomkdDDRR3MlugpiwZozjPT6IaAnkVvrSFvIOSuf3nMl5fONQ7U26J1NgXuGiByFX
U3b6MkwouR84/eelLjrSEAMOKxs/NQonAK8EHu1Fp7VMKNNik9rNlWyLHy3f/lqgSW3kvkGy4bHd
v0AvUoDyOlaFBj8dEFUMAf+9u4Vbc5Hx/VFMGkqCImpGI4FQp/Tg1cGN/wDULn6IXIwPsc7kNcbw
fiuBmwtd4oE8/0+Wat2txXDpx91BmFlpbX9Cv2ddYjX8jkD/XgVhbb+tnrELJGkgBuDasPSFerHy
sL+JPJXZde+koqLqNOHweC+1IrvC8BEB9vlI8kAGtkAiKnsPpDQxYY/TUoOstZ+8w+M72fiMKMW0
FbpVGtR2siaj72yCsRICZloDEsF08CIsRNzXB/TawUHmnqBZqer9VzmMNiVc0xEdOdiW+worYa3p
rVRPc1tcvNJNUQFugLRQh2TPZCR4ExGrEkVMxyO6b36IDnXXplEVd8g6T5UyP4ZUxZje4/VIGw7Q
sDLISTt1BSdIm+L4OfEYrdGygVDPDc9+9e0CO03JzK4/P1B5oAaMWB7N7Y1UIBsevH3JG2z72/JT
Bs7Rk/3dFTKW4QRU9f/vtlILVvveeYeWVydhg/WT000f+EnMgKN3nDiwpUz0mvB9GpRHNX57yB7f
ysvdq9WNH8LAbaBuRejyjFKxwFMbWE7OF8hs3z82C/tGDw4XBllRO35t76vjgQqFSdxTlZx207Eu
1pPpj+48Wr7x2SlFm5QhwgiW5t5o5GdLULi1qTTAeJwl28orlrqzI0XiaGi4RCTp9AUq689FwcUR
1hEcb7f3PbsDSKtCjhy92OucN3uyb5VFEy0pcnijPoAjV9cTqizeXuvbk60vjqALPX/b3VIIX7JI
F2LaCP37KYThCNnlJmDfdBwDhBKfm9FyoxdemAaaQ2P8X9h6wYzizzOHM7dN55xB4T5Uz5zckVA3
WutoqHwSlfxLCed/+rwDiTjQ9+I+ZVQ2jyZ0DeSa8c36JcrKTPYaD8vvF8J1MC0NKXdG0YRQw3Bb
esJR2ecJ4G7zx9LAfbHDGG1BZGuJXeUCLSQlk4tvDGKdlNwrKIo/doIlZMA6kdgv0p7i6AJc6gth
gufspwLKDP/V4In9xDs33tzZ3C3PbmGDqPN0VZr3gfbxUGoBE/2ZJQYnFcXCmhsTXD3Vo2AyV1GY
GcHfS5RKxgQUqDcA+NCxntBD+cq6NHdd6BDrRwbmAHbQkWpFjQjSlBlkhn5ghQOb4rfknM6pPkaq
7uI83A/QIMeUEdqQF/S/VDB6Vb3MwTtAMU8ZCmC8JMRwnkJkkMKRLRpbK6Fe96H43JKQg9aQSvme
888sxSW+7km/ZZ3drGM9KwnxiUvW16marp1EIR5Gaku1QTzGiAWrMvZCAS9dzuc9JaZM8xgteJ+Y
l20p5hfz9GhPvPzlCXLyjHmaOOgC9oz0PW0fCsndlmP7WXWDYcB8U5I1iyPXS8v3C7WOlixsOkoS
FT/SbIFKC4YxR6G394uCOoNIBuDNuS0VY+8Ewzv6n4ktrioKA4lGxsqzEmKkYxsNheC1kEcCjQI2
GjNGNMDEEATE3IKDJRPn+9ySg11NXOaHTpAV5VegUG5UbBynQLZRSCYDbf2Mbg6fGjk2PsTWwR7X
/qOZMTEnYSZTBWfkgAhNMROZwqm06T18nQjrcXwfOLqz/qUkJLaPTNXy1mC+MmDS6fuQWbAbBkOL
VuHOzWd85tpo/YXUVFfOmp6+FjNtQFB6Sl08zb7pC2L3AO8hMVz2G4la3JWRLxy3TLVxWO26y4a2
kxnYqk2gneeOdwHWupNrKVrQptyl/8z4qsj3ealVOknKI5EtOnm0+8YvQiaR0ZPOZzbkg6+R6pPB
1m4xfTTFL0bgR6t2H82+Gh7tGhJ2zek0p7vRjrh6vO5Fpn0lsmIiK1fOZwV2FnArg4pK5vDtoP7U
jEknmG7r4UbrchW/M81/VjG8LXZG6BTzw48mV8MBuycDFsO+7Od8Qu8THMnCSLEXfR0db8SuvlMG
dO+JQTE+yb9gUVLI2t9cxyjNHijDns6wupbDgLLmxheWME+ROhXQdV59zTABJGQ/LCt1Zr249Aci
K77RJ1bk3a9xnVVCT6IBdchdqM+poD2sOzWQC9ME79zracHhlYekP0r5ymG3QlPQZW9DEsHQzEkm
8CIvRafWQgY8aIQyIsxS4uoUdesMqu6VmTRI0FeLSShwjKxIqbNR+7XdfY2QWis368wiuqcgzEqE
RPsInYqtVM03YAuqCGcPfefRYDyuTVy5PbmsQEbZlI1dpH0dgEjn+UZgIkRczX2WPnwad9Ze9Vv8
1N8pc71puqoleZqZJyEK3aFwGHwEZzbmVz8O+wGVw1qj75/l1yIAj27z9HSp6OAFqRIKaIpx7FWx
zSBtYQ9wru0niGJkNeqnEVIq4+vjfFJ2/rEg3LT7h60NMe1PDMgAwMaGZKakT3T2LUYnfEhLqOul
UPPM2wPh4ihZgUhH30DYwaqufcHPtwyz0pvdk9QvdFztTb9nAIBH0lGNVMsLQosB4vqnX8+9q3CZ
wXBxXFVru9j7t0dTjSd3EpZVkuJDoFYIMHmWSRytaiIgej7EahGxUC1YFDDYNAoQv35Dd203iebg
Y63yGLUMjT0DtqEhpdKV0zp4jicXeLvenHCQw4k7H6uT1yJtoGzRec9hTyhLb/v+UP1IB3kiAgsT
Nu+N6EDBITNsz7HxYcLOl/9udpLpfu144YdSbk1XmBGt1amxOmaKAWu6wtRE1MLRPu5Vd2AmvyVk
Z5dMevAou0XyQ6ZhkwZ39sq7Gdjb5GJhEWgYgJtQlZWXFKnpZvRTBdWy1sC9hYgogjkQfyUMfplO
6Wqh9Hf0FaYTAsnb2kSeu8jgp5oK75ND44xZll53WroWeeWEXtVI/ullfCfoD52rxwrRHskYZ25f
XIdNoOY5MxKfX0qc3OClonGvNgWbgB081AAHN6PhPOoFCx9rdQ+nFmmJVQtFnuiw4TNQ1oLRdK4X
5d9ftGROSKGQkKU9FJyauOPnLFkU7g/l1WarYZfyPoUhu6xVf+6FW7aJ+zwTRNmJlpDre8jT5xjg
Y5uCjptl2/edB9fs6GsBb+Lm0WPdlW0bSy+PbXnqT+oO3ekaUh4j3e71gJ3UflZI8rOaV25k9pSL
WRq7fLha5pmzw3AlZ6qVUKQaWGoyyXziOsfPR8vKc3yi4Y2fk27OJpaZ8Y3IsN7tN2XQPhEwl1c0
l93ANJBUqK7s71aEnpHfMCH+WP9LnRp0qJN+duWrM307JD8MBkZ0+ZBUCmEpeAJBdMMjOj9Amu5A
+PHSBQgHVd4994Dt2rQ47dhT//OFOZH78ToGmG0/MqjvPRzxSEqYpp2Wx7uHRwiH8o7llvJ+SHSF
crewOYNB65m/YQtUjKdIIH4+ZphJo6ZdPG1HKR4vc07wQq5WEYEfb/93oenBixAq3k8qwtnAr2v1
5hjHtdu9jN1gadwcwwX2+mL0yIyziHzD/l0fdMlcPb4dzzTHJ5TqvncAQ5o0/8sOMURieLgHAyR8
HJR3uAujmCgFL+XpeRgvKrj9JhBKh0tST4wNliQGwmObTaaD/aJH5Z3oTX6PeuJhjzaN3aat9Nu5
xzvAis1WEo9c40YDk9DNVDrzq9DhR831zOxtjg2UpTAyPpahkdyhfWUfwxDTO+Jl2oxWMXTjoRrm
8aXvKs40bh+PtdfMXxJYPd4inP6hudY0yKA9kxzJIE7C9Q/rGOggb0VoqUBP7LVIyva4fYkQ7isg
xq1/yFA9+pQ0d+y7/5eVvSs1rcaKYfX3GYxvbqlTMjyR70p7x+czjgyhjifzL6eA/lP+chpKU2x+
XEZX14RC0NE4zExi6F2bzKG1Xo12HqsH/X1HMR4HcD93Jl6cSBbsbs0x8E4yHNKGK2hXuhgAqOu7
jjsnnY9TH/NY/b1kJ0TLwAkTojBCY58xa+vybYlIaeuNy59q4oFosNRDnGlKeDyg5jdAyfSM/CUH
Zf7ctJmemEkX0J+4ai00hrTuHeZpRuJvbbw06YyQygiU7PNY3O9iny50rp1wYyx33fxxu+ACi1xd
uyflDTW8ZswgogWzBJ7G2WeqIgXRzsU2Lem9VbBAAIm2VoUykMAhV00UUDbZwqEJhpsIIUx7VapD
ZTSfNeM1b5IZQYg4+VmdRDwNEtW87Y5xZeF7B4oSHImN94l4mE3uwbkuQa0ToYYJS/h4aOH1ZN2y
QpGebbofXz2OL585q97eB0yABDM8Nw1x82dIN9VeYN39rLzqMiI6O4EBje87C1Ecl+I3BeY+w5nU
w0lQXMAodPjM3q/q4Rqkp2+iwh0zssg/5arNAVPeqtChWkqGqoOBzbYu95AXwV7Og81twvN30aWD
QpP5tED6gk+QP7oNxs9runLPeZq1mRRhhV874rgUJgTe2bqxBRsWijSxy3ScoYXNsMc8wKDzm4zZ
x4xKZYnS30w2CydZS6UYUWiBnD0jaXlN/gwwMXtsquDAqyDN397p2UQizVdaLb71BU5RfFyo/E7Q
vhjxyC3fKSb+ccO0OLjK8JSQdOYXgYvL08F0e0LHD8WexDlwoATlIg+GjjK37Oivyrqn0HyHf3ds
zP9pbs29MoMiZt4/955UEZB6ywXCSSex5VdUJjDRrlJWM0OZ09WYJdNvinRl5SIL8cShaFNGIC87
aUxSuJHX83X3+4PE1QOpeayhy9PMa9QlIOEhIQX7GCiUBLCkRgiJaF/18tsbtHUcp8QjGA8cb8fC
SzkVS1fLYcuXk2a2t/EO99B+MegUg2i82Rf08UegjfAyKQhwSELekyQOaUGb92O7G56v33en3RRX
v4T72PdzyX558FE0ySfG74WhR3EhEuzEXF6DXVq8FudKRFj/vpp+8kwpE0bwxP7+R41b7bclzjM8
Fg1YLzGzmz3BBHTUOTBZkxB4VZhMJfPnR5nqDOf/pQtJOVvNSSjvCwzp8Y6ihc1LqZLnIiP0zTSg
fImtrjkPyHWQG9zExPDAv9lsWWlOYSQLd2u3tXH4MOjl8UiRytIqh0/Hm7HCwR2F2sjScs4eSL0j
hlupIQm7Op91bdIXeMjQGQBLXuGoQRdmY96wrEouVXW5iSCeFYS9Sd21ae9W3RhenIVECKZUFJ18
5kIK/JTUHh0a/Kaawkl90qu7Tql3nUQhtYj2pMVi+I37Rt7SV4qxNN1ktdsvbVjNRbG+45BZG4KW
JGXBxeSBFzwGByzUx+csyWqFnSOua2ei9gcU84EaGqAmOpsuuYmUHwzLr/9mTNH4dmsImQKn/qoe
yOTfP02Z+w8tbNrQrz0X+0qzXQzjcnx2DoaMb91ViSVlio0S0NsAyYDSmR5ggD7LNQ4141qdpXqO
j+e6XE56BD8XsZbZVN/nxaXXt6wi23aU9gaDIjdlV7CaarcpBWYHGiedIBMzkDzbrFsVTkboe0BN
Uy3FID78/rzbYYD/OXSHpHNBnGThDQPhclquc6T3aND2669+G3MXq3HxEaTRL5IFRDu2Mk5nfWdU
bv4vHacsg2RgIRDLnYOI9RitZajcskaZRcjdv4Ic+QzwcZY3r1rIZP7+IT1SgBvmhkw/tvXjHWIN
Jt2uzMcEVpsBtiZZRaxfed3zIl98FIarw/Gbm26AOpp1kJ9A/TzxetW91078igLq3PpW2fIQ7CXC
a8KjabOTNl5zf5R5HGCjZPyUqTBTDtf51fJ4q0+x3vOXTuxGNz3zWVSBHl1NbgFVgwazZHXl7F14
CXbvCmCuFQLJGuYL0UEk1pMD4ZPxj3oANPjFTQJy7Xh1UFPhrdiZztFOdVXCfeIQoZM22iOMEWc8
lcADGJAGfH00h17gXq9Gm+oBzGDkKrthOzCAt3KkBbU5ZQy/SNnKDZN1JSbafPGI/tzAeWw5ppTA
/F/TdzaOLlY3inoKvHniXcMnLueiaRz1rvC5w/KJdh9CuCJk0UbfHGxeBr8TqdicGPawb8fc/esv
pHRkCGqUsy8Pc315XxzGIfS9+WeM9+ost6btfKSXxDCYF9dDNe2ArUZU8lmy7qk5alJ3P08F3PMj
Vlvt+KggHTL8FMqePhEvwGPCPvWHaVXW/JdHNO1B59DubsarVlsoSF+iQqVI2sYT5iACNfL3g4+/
oa7kAU6LyRsE34Tz+aassOSEoVy+pBYirsIvzinThSUvskdc/GK8VTGBkLLm43fe/RYx7vtyPrt7
iVQDfD7LUkaR8dh3JbvBEMl6SHlZEip6aZUtg6gtq8D/ucjkjdlZdsEEic0MpVls4S8D9DyLHGdG
L4nW5Bp/Hmr3hy5ttEByUAP6isV1UsMmEH75YgI+5Z6SrOnk7JjtUO51hU64h2F5Am8+22cD0kc4
mJvTtWu+rKTTANt1QOYNzgd5PgLkKDIsrPMpBx/+pk+jyRk4DTmYJXtmoKjxnm1V9nyUKPaA924s
akqiuj3ZNMP9zN74lPD9NJm6YKVLQAVLZ5MxMbAQHlGhvX0CIbbT9LDJLL+6lueCGuVT7CGMEMTI
P7lbx+Sl4dzc27KTKG/njF2LojtMEfjgJ7kN0HUJJepgTMrtHtOcOYje+oUCze730wB5CBQc/xTX
+/4+NlrxTgz+H7+JZqpneC4VE87cwNbRG1fhmrzy/ZLQFnkivoz/zWxmSIhjeClE3Zq1EEDWaBQw
4avbLzsa1sHlFVhH+LyKJeJ790b0dcjhfvJVCjy31IAsblnySYzXK3pDhVpeYRQMndBY81BQSG2o
8z4npk0DMonAgBr1PXlPLuJikYfc1swfrGrnmMcWoUeTVz492XL3/QtyE6hNbbTwP7VLxdE71eLS
SYU7NJiadUBF0HQnQa9CujLT7+5AapjBF0q1F5O2XRUNzva7Wdqkf2SEZ7ECOIBJGQavntl2CxPA
wENr29hxfM18LsweReBnn0R3k0Lyv3XHmXSLCIQMX3PmmR0qAg3462O02ELb467g/krEcXsxoVJS
3S5kQ/cdffySh/UFOdeKCNIl/zRQs5izJr1+7Q1+KfRVyZTKh9Nr8VzO6W1uAoGLGkytCZFiJcXa
xXuPvjRvcPo/17VEYpIcDQYioHcbzGvOPVlAXEO3ig3hpY2Dx1CTKDjMFHK5a8KIXLp0rNcLkkph
n0yVnbYDXnHtscHiDvLgGnewKmF1QjGKYWDQJZenldmkawTYIz/muCccuuLc8Fg7V6E86w2ldcvE
gCz0sS4SgBQy8wY7dCWWaAdepHnPNqu/Ko5+UkEZt3my8gmfSDnqKH9Cv8PJ/n+1YIlAjgFXK0dO
3BySdbt5DWWuV47sbdyNc6b52S6jLOm0VzUmEFvx3V2sqyJTrodO9+3PHDBzSL5eZEoA7MwuNm3i
2CfXKw7e71jGtVIBBh4c72RhHb0OTkcKVp+EVP2wX9GED5jtI6RxwzyoQ7G5Bd9aqWJGmNkY5nUL
kcTSGlkZyscmqpFazDpXX1OUddCca/PuUft3thlvNOAzymse55uVF5zqa6++XS+lLT7yw6Zagl5E
QPLiowZleg/u7ZY0ZLakVExrByA3NiXfRjrzilzM/JG8OOOXFWPV7sGAaUGZO7rNqtOg/s/nD7ys
BrLlkBSW1yb8Wj0WpMHBnnsEaQi12C0+G5coWIz31DOSeAb8rBW7ZQm1lJbowAy4MjnODgIp7OZL
X0mOAN69nK6SWzfiPp/SbpprQ3lydE6w3ETEOFEXMIbAVCQpQKx99KmN3WnLxn1WrH8Juf1h5LY8
4uJgDHtIOEMNSr+sKzswUJboPv+E4SJYcyB1+1qKEnHBA/vAz78Mc0CbyhnXSYpj8kfCeZ3dbNou
v6C+B6SYURmGU/rP0c6i53nMHBECtMKhq60Jcr8eCDDI8uXEkDlkmMqxpt2XJ3EPE8d4V0Hx+mKe
qHfvR48lNi/g8SFKeZmzuwjX9uoJsQNatiYJPNJnAIuMyiamekHmikzhgZ4EkwpyGuOokdVM9gM5
4B/YfDOBaaTIAsv3umIPAsn3uxcgog0E4vN0rgMBa3JMvZxnKVtJjQQ/kWXLrn/6HxKUVDyRPSXW
UEGZLY5z9l2V2EEt6ZaQeXb1O2J1rovRHMg4+MXN+9fe1d3r3c3dzT76B96F/BPU65nV3cuvgQog
T9LQG7Cjm+JimhJdvML+VpggXUMz8fmrQjmFDPpRz4kQSF5Hr7VOtPvBw5xS7mQLVGTkTCv7vmo/
vKZ4fGGF7atLl58jFSH7w3Mjo7wvAqMP2MxPNsqC3EScP5b6MHtsAS3KgUJOJYlMhRgTYr5d0QGT
e+8RM9e/+PhKmB9bS8NQxYCJAnSfMPGj8hOVAp4BnHNEVHvMOUzNV9e75lWEqPrSalmP1zq2RT87
qfxtFPUnnHaSsXJODz87hjkfeggc5yFM1UvzzvXcfMm14Ev15WQ5s+yX5/OudSSomM/HmI4Bynzw
uAzEi9bCmOWDHGkPbCBoUUon3W6LLFPRJAsqnnlUCIV605BjdbGgunHABN1SoQjvJTYZvbIYMMSI
p4aFExhEI8+REFvkrvRmnaTakmk0gJYxu9wzSjgn+CK3KQXyzzKotWHb7FdH7Sp028HSoe4ba+XT
ha0GardNeX0a1E24GFF+vpsUk9uhf5SiniAhx7jlR06j+aWGbVnlETG0iah3BFa8yuBduy8ERIkg
/xqd1QzHORbzAOPSmzgx5omCJdsfAVNOXesi8UxBR12w5NKfhKvRISvKX9AH9RZWimK0EMbfPi2l
6XlmBspT+COC+jLZP+cYf/qo1lOVmQPTZ2HOhubrCfj9p8uOPy8Kxk0sD7T/4HfNr0ht4mvB05Gg
FJOL+tGTN0ozVdu66BDkZqaSob+iyB/1a/vknuHUZ9SIlLnFw0aq8wCIDszRABFPjOpCAHF8cpNA
5jXDgV07/+4ih5xJIHtFhtLrb+5Krogl4vfjkbES1QQ6Vdkxw6t1lcEqSOGfaKzPqepmk6oKGFvr
02JZNXyk8dD1UxXMt4QrcdcZyOpoaO7yipLbfBzuOrjvkpomK6b1UqESgssuMEYxWW6MaU9Gs3Ag
dTmfm8BF+RoCrG3Rd7M8f2QrEHg3504ZmCLHVGd9abHNUyE5cnK9kSFWFmfkvJyW2DOfKD9cnKAM
QFAUD+V7dsoLDBKuuQrzWDkwOrkQy6LueLxVQuXrKWGA5MQ2ywBJRPKKH+g90zMTSB1W3GdKC4Ep
Pis5OeN6TzCGQT1IiNBLefjCgAwUS5hqqFkvee0gt7rqadjDRoEVw1til2fWajSYK4s08q7LQQnf
CgPPeOHMlnIfGM6OD+C3rxZh+v1zKlgontyLBo/uI83Ckx6BWu9rM+ZQy164Bzdp/LQSlDnwbZgW
yCLwd2EfjxV6TqUyvZknmrUHgZ1fz5FX6ehPjB2U10vqM68mK6bAJCnfAA+OldoOQYdffzVqXOba
CnJmZVWVPTviba6Lo8PoqXM4kA0xgTW1+jodmsQ0IMQ/rCkm9IOQM9Cz9UARuvbgsCQGl8N4nFnx
RRYRDaXEANyuIV1QHZnDXNr4JQIy8cwWfWNzk2ObdueRL1YPsX4sHXlM0c3TwnpmrbMLnwpErPv4
0FR2KwFYXYxN7h7NbdeBycGUSQrFouXcw1B1gd72KXj93uXP2uI9N7w7i+Jw0svJI3nLUK2r3mlz
24VQkK0gyk2u0b/0iiIOTjdpF/39bexM7SCPMTdud5i/ySYstYSW6iMR0t39lqufFA5tqVJmLmez
+dOu2o5je/wTQnnlKU2i6vIIhQ90Fvs2fgLQV9wMC6htQJ2V2P02gtWqFfLs00cg8LTx9kGSJFos
21iLlKjOSJzciVORpcshdr5odMnYGlzycDg6NsiY0zM1ogWsqiIguqF03SPDCddJ16sfyAlba3um
Z1aiu3CaKMpsijB8+qzgum/w6y+P1xiJSmI9bihwSQ/wbyz0p7mtJg0bb7nKsYTpcuFwmmfbwVGd
xsAwoxNj6IiNDO6dfm5oRiZILgaspRhVLZEca8nFB+KlhA6+dTp9M04vmSePpE8CsW0qnfUebWMX
hZYlo2AXdhS8/yuYfsnYu6tx1+JzvKAnVYiYE9tKU5TtU5RtlW+F7+TdQhLlwrhsMr/V3MERdAGN
5Ig9+S9mO8XPJElMiF7ifjShHru6i1DInaPEAKebs07gltMaRRsYOimfxHNZ9ojz9yHnWxcB4bkD
VP0A4M5Z46R5QEiKLHyj+WcJ/ipkfFLThKaj91tethlxQUVO97jsfvGH8UAZrzG1c8sjtIKPG/76
PQVdZ5Aaf4wj2RQoDmKhDhz/dm2r50dn3RBpTggD6FKs1keoPWPosZlciPnYKLTAVxrLTSn4m3by
gRlp0OcT651z8Ogz6WhVDh0//6dWE63NkiU22wSfbg252DGqg2DdkpVOMSTAsztrf40YFuNiDnge
n3Bb7TYOAX1HDH/sv+HdgcjrUqEROnfNtrDP4J/wQT6rTk6PCR2NSaDlIEggl3nN73Abjf+MDu8I
f5HXBIVSUU4Dwj8UHNV3kFNmoA2PLxvb/XBxSRAaw5erXYwY06kBHWrTfO4iXJXDzXQ2K3h33t/v
YFKJQG73gLrCDDht5fHbu6Qd0qmwogYvSHBfnXUaGVSRurJ4iziiHj6hfeFXZweCPmoWXQclNccs
w69mq21yAbMElyNJ98c3/eczdPG1Xobqd5F8qI883krEf7f+B3UwWJftQr3iZuY1YYsiUUh8yDAA
4KYoQ5ATIkvs2PVxVPKDgRp27sTO+wWOpMCI1S23WnF0SIWDAPfw9UYJXQBsYZQnu2qlI9vFj/Ww
6ZQx8uXYtusRb9hWbu9TvQgpz3RdvOhlbpepM2fIf7Acs/dlzRHBrqi3qhRo4Q+Yq0uB4dO1R597
4wxf1S4R8jG+ofKfLP1Zyy8TCr5zC5boIgTDtBzVEJu6cog2wH7XxMCi1s0dbtmqM8xqcxnp75wp
iAotNkVB2Slt9PGS+1WYeT8Vn20Rxrx+FZb1vhMx3CWAzeBCCf/VsSIzFwC2jCMPW+191kMM0pdU
exIUUHqdYb8hvOupW9uK+ckqh6GbLA+mpWolISbwOZhMztm78mja2tLRaHSeALcP8dqb1BjhEh5l
eOYIOvpR18f1B54Y5YLx4scBa+/dvEIg3YWalWApEGasqpRTQo2UmVZKvsXskW2ybJ5+wszRgnga
Uj2VAC5rfc+JDJoCFnroXsV72A12YbHGVw/XRsMQDBiQi0VmxMhjIuHw2ycnxFeRES27pacYNrIx
08bCyHwoPIXdPO+BLbKgZJtWMwio0jrsa4NjqKJyfyqvzNRo7iM1JG90YHxaTKbF5eYB0ShZDVS0
0ubw2kqOLFCZME4tfp1Fa39mZJFffowWRJbYPnsYqQIS0inzuMHMZi02d5jYvus0yrorKkcE5I1A
+GZ1JAPD6HDxesTIl5VO11uY8hqyfr1uQjSZyVGJQWnWXtMVnR09vXi8t1MnRP7dFLYRcKcmKayt
trlCR99x7GxQqcQON+CXldS4wjWkvYJzxB7eDRqlDJXS8u4Iva2VtGoJJhqXzvvtJL8yG3GO1cAI
9icGdtE7ohwl64g5gCRFFF8KKquqv7HRjcxF7Kqkk0OlMad8iIDVh5sp2ZDYyv5ev7tgQmzrQkFp
yGP6wmmsjARTJ3YQ0D1vgj138FCYVIE598Xwiqiy6sjwLbQLmZ6Jmic7cKI0gQQ7VX15iKDoutnP
ykMCv3NhfVdaCZtxLrJjFiNI5lMqMVNbnRlMca4h3Ogj5ikurwxmy0q57wKMbplc58/uGrOkaHP3
TnmPmhC7mfZpkAgw6vbD2P3bI3clnnJmPHOf2GQDc9FPXaSQoXNihtbGwJeIsx6vuOtU2DNKdYTW
Z+HaLgcOlYqsZu2pxpOP+coNoE29kV14Kfum5ZYa26WOwRyQO89mgMi3gKryIheKs5Mt8QtBq0CE
6BK6KPgdPeklyf5TvflgeXWhyV6AOiKDxcIp1EGhN+tgUBy7YNSnuCeLpOcXEIC8Y1VJiJTeMGHs
B3FLQw1fz495cZ1VKgIzgXiv2JawWiHrbLBasDTjccETLcZzd44zQ1GSIdPvpzS0ybsL9Z8XOzAx
OXYTejaJILfxtiGDRacrNgHRpciTn3JjduFWwcCYM7YA7XZ1B8L5O8pasQ3pgcU+stibwQCKcW2D
9AXRjcjz4cl2ceOXkHv37BzApHNiQtOjcyR0MUBIi+1X3hVGSLLfaippn9sdfLyWu1f6vFZWfpgC
c4zJgQgpfBE5JOSjS6zx5HTH2ZrZeNRiNDmdWejP2IqpymyVLJk3YLsK4+ew5H1E7o5IOVOsPkFE
EG0QvPCavVTZr46Lf7soWlTTal5Twus/u5WNQYJKHlpDEsvQfDEbnOHIgds2eWF3Ki12QEA3aqD4
W4HrS6SwZzF5Lt9jKH8vD3e/RreitSCuEa/FaxUmnayPZlJgUiVxTL8E1W2trsDIDGBSVEScEc+A
Br75+y6PP7mQFt78aBwP1mAcSdXzLbX9mk++Y4bh5x5iDfWV2/8iu3COUS/+2qnb3VFKGOUG58yE
FM+69oiwy6X/xESiYC5OPG5gj0RpO6WlkefAoNoA5eARka//Yt7+eL+4Q5LO1X3ffemq/vHySebY
PH64/mtb8hK0QcccEkHRxWWgjdqg4WBn1b3WA27LGKbBSgdVAtXtRk0WjpMfgdyeFnm2ucOXcVtF
ZcQg2XNpLT5RGCUPwoYjlQbUj+TyKAFjxZwnZqFYoju885a2YB8Kq6wfvAr8ohppsK/DkUpQXjU8
DhIftx5Ymkcy1gIihpFpUMF4vorHe8yRTAfm8BZ9pmdkqSFh7DCtsY5stKRnI9Zck3gmJ9s5YQoI
eolaGdZ+8QoZiVdrnyoF/miv8paJ6/MilSYYPUsOnaVireA4TcjPN44WnWSspxL+kz4B8o8viNha
sIFPkQKXWarDiyYVo5FIWprlW+XB3d9utP0oXZH2pAKFL0R2FfLsELfHosUc9ttA2ntGXG9Zb/WH
bZmH4VKnMUSDMF9u8hQKTkv7uhPgHbFsMrkAtjo0dOYBjoz9HNk06QJra+t0zUYc7ViZKETLMhLa
e7yEmz31i9M/2cLgf7Rc9ZmJdckqFxbvAP/eURU5ObvjJMvxK9W2Ho2A4M8Dqh5+s94EDdpGQHr5
Q1OrXAXSBm75bUXVFtssnKE2IxwTYZgq5uW20QDtl7arc8MWL15uEGmB/ECCujdNRCnHvogQPIpL
ArYyrTFQFuCzRAlSNNVZelCqrkj0EVd1W8JK2naTYtNF9YoUU+Vlz7Z5IYNdjACIOxyo6C/XzmXh
yEAYeB8aGjNVY7gNW9iNfgAa7DqDBbIXW2v6l33TKok9U/ey5aweQK4H1TgSWoRktOFen6/cR5QH
4dQDTPHY/wruoLXMVsoWQotH7irSzQYeULPALBK85HHWIj0nUKN1hZGB23y/Xnvm17yVmGB4oDuG
mJ1jvmNE8hEYQjGMxLoXky6XJNL/UZkfPt32ZA7D52FzSURafUN2XRMOiG3M2bxFrSgBjm/oI9kY
Y6iVBFtisRqa1NuBadAtIaMJVtIJyO0nAH1h9/Gfn5RYg4maCTQOffpxP9t3OxURoZEA/HGEhuTL
vWwmE864Pgh3Cs6oth/zPm5Lcepep2MSZr+dy29vgrcy+dzvvdhqNKcv8CPJL+wvXmmKPknyBv2/
2WUHE5ocq+zvwf5TSoAteTdCzjc4Yz2aUoBzXajRc1nl3zkIUy5zAAvkNHo2SxDBNLa7pGEUTwDf
78C+h5p7HK5FTZCtBMPOxQKUKA5E15+DpHfQHGnahumocRzGhhUFBL/ZIzu4xt5cThEsLdGNxzzF
A2J7P9M5FfDJWYECIZj0x6XLzkP3HM55I4SWDhUJNbj0lddByHubjm3vz9xfC5lcjGtHO5gRlnA/
CKaTrOmKO/EEF5OjgXSlujDphnqi5oXpWElg0K4JOmGPf0u+qQhPx2aUgx897XvNbrZEs7SBjBfl
A8BQlmXFcv5q8AgXhs0143VC8tr2fbrSKmwHND14Qzl/NKmg1BTvrHLK4ur04Nr9stBsKDFz1jdC
Mw2voTRPdVc4/S489YC3f3qQzIHiHsv0x/FApCvbI/Wc8ZsHW8YfWAwlaWw8nEj6KyAufpLIcQts
WfXcH6QDilDlEM5zjqzqIyWACTFVNAMCAMudRzl2dmeEO3u9/DnM3l0gpaVRNYKC6X6aJf5P5WLa
VOP55DpKzqlVZDkTTuFENMyJ9aPemL6b1CH7aNVGOdihPhZv0KqpK2iNC2Lbu6OhHAxjuyMkqDR1
CvqWn9HQXGfad94/3qKUd8JzWRRQmm/nB2nIoXoofxGnqYtmS7lWYexNIKJr+YKfU9r+5cWks3St
mrCAgy1LRHrXkfTEayDe81Zs4oOHUjheJA6rLYkZWldYXdpS5fICDYQZCh0DUIkBc3FTb8Ysygdx
iEXEzJIYqnTX8Yg7BBwo6Dt3P04VVJVZ8P/iVYC9ReHGPBYTB4wf+egKYQbvyfDHowOWREWsqQOI
tGPRkruNtRQJBhx7tilKM7Xq99XfFC1P++aHH4zw7DG+kCw+kwFFEZoQyp6qMQXDXtbs18KpDgic
QdOBbdGSPIEdUiRAnRWUXuivvso9XG9FFbedooMcw4OVOexlGwaUN++NVOBNDa2IgbrQZWzFc3Wq
yegcK06PHkvn0R97fQzo6DpkFcbz8IRaqTUaPOI4PLbGWCCnrMv+QqVvmQ8DXYsYWiv9XIoDCHpT
4vpPFNGMKlB3HpBYIHUCrHioDa1hJYmoCipsouyjF/BUmoM6LR3QYXER+0GY/AfaRWKw5nVjKGw/
3RAod53I6E/X/JrER2INWJjYi8Wr5qvPLOWRpF/6uDa0wzGBb/kvb730d9aaJX2q6WIIHResJ+BM
gL0SqNwYvKSULDbZ2Bj/yA8AnAssREKpYLNn5x98lvs+aLLnbOFuy5avoicm0UbfhmJAtIzu336b
cWHtO/5p7ULyb8UM8FuCjyDQ8e8ddxKBY/wQYrDA2ytEigIwJi/qQamt0hZCv56teb9rd7Z1BBOz
9A6igySCS4HEReuUaE0gF+UB7WQVt2ajNibzThpZaiQztEh1+5I6oZcamOme302aAvxNZqUmWTUM
SUNai58ahEifS7CNr09PXpZRTOtp/A3a6dPam2GoF6PIoinrTwctcJMda+nWthsti1luHz1JGZtw
CKVdbrCoYL558GEnllVoMyWNusHES1ZRepSfYukS+CQVI9JjOH9I8RVYygh/jdVk9xD1fYZuV5Tc
Md6RAN8P19hqDOk79wb+3nHxowTUmuGj+KtHDJF23a8OYMg9NqvZsrv1Oo/RPs9ZtANFNCPjv+lB
/Ea/WZ8BMFiUzlEiXacW6SaECGOxzChYB8DD9LIoSXQkDqgiiDV086fyrzznIjK6gLQBpzjg0z1e
VLSWWwa65Mf00I1CwpLNBZNYLHgKfZNkSJkqZrmlWWeT/WXLFWLuPRVkF+84nra78rw+uzUltQ57
dpvWn/ErhYAjG95nUQBTuXrwtsEh7xumsXcXBJ1mOl003VWLyD83jIDP0GyutWr14CGY0z6Y693A
mNN8lyZ57Wyo8S5bBebvicBwrWBtzM853+/9p0XjqahyyvrPi5K2NWQwXX7v6aRGY1DHOMUIaG8a
/A4QyWBldiWzTJtZ2p/USkfUMBR5vpaH+sqmcqfhjmMRS+WX8E4vKrd8kualSpISrlCqCCDvx3+A
JL3XFopXwbDl/nGv4LMkeHoysPz/09UqnlOWdjrliJHEy6WrGbrEN5+/Xns4a6FXsbFSk/fwwdEw
kG1xASpV7SjvE+cAA9iWiTIvWDaFUw7bmnoHN7MpDd4fmcG0cJvTK44yWL4pG9HN2qtqNIXPoQtA
p4t7ZoWiepfwZH88h2l1LaYZYzyV3bovUeon0uUIPWlIv80UJ431Ynbdwxp66fQy71sDMPAzg0x7
FymcjoK+VngT9T75hxqjU7CXQzB8t3M40NV954CdXOYLRWEbQvOKXbnZFEfQNbnuLFfaN8R3nW4X
ca8mHNhMSNfZR0T0+Am0DEFkWXNJLZHJezM7zQY7yLYNEgvyagYqyy9SV1PrIZBGYxFCcycPXrcN
eVb98i96oZgXsQhezfvw7EsnYhEs1wbZX02LHKOptnmjy3SJe+aq8H6hgTsordMcW9X/C2Egh92T
7fTSpc4ghFhyUkA5y4DHjizyBOApBGiZ/fgrnd7AxgpLI8XF0I+mnVi0Ml03RcX3N3+JDdSLhkps
i5SPhSAf2p3ZBufl5DaFYwGm98ONIfQ7PFhUgGQdyHli8T3ybj18HNkAH7EF3AzFy6S66oVKkXUo
MX9ISoC41BCqXU2IxG4DGpeG1taZy75crAy05zw1eY49nL9DlB09B1gBVmC8on+rl1xZgloLE48T
bFILrR7d0b33sjDWz9lra21oiLqpVrnk3fApXgTJ5y/SuvpEMxxkgwqdDdgvXUAM4zPiSeznsj1T
oBLJve8mHKVNfVrz7EI+WYkY9TRhTIKrUm0KgN4Yj7TnUur/xjVQUmSI6PMCmQ5gBZ7FXG/2KKuX
pz/tapsgSLkCPpQj9akFoOqEpFU1s4Z7RAMyqho6K0irOPreSzbqW3VcTl+VdjuxSJlvjqe18ROS
wpiLFCALIo92p4VdCa0MLMZF2O+1KDIod+HsKBZcBR2E4B+ZkyplghV7z0XF2D8b3qos+oDbKBsn
df+Z0aQ2WxGrQU+3gEUe4PJZS4ClFA+hYyOPKpO4m3bMiCpYlpvqtsQhXZrFVLMoCZ6QMcKfOcRj
eImdrRXaQdGeRa7gnd7H4Yf4RRd1sMHQnouN39gbXUCE0OJWXJMVdSi7J7DjJzy317jpSuENHNPl
zyyoQZn9GMCwdo+Adv3lziG/EREC5FaPVVnfXgIvBxWnWxhgWWLXcitXWwcqMPl+NahViGhsnIU/
wer3qaPm7vqzpsmvbbKQ4I4Y+XIC9EL0fjpjHC9D+MUtPQ1PkO8ehsUE4yLF//UIDMunJ3JgB7Tr
wJYXtcWsl3LaexmAIa+peny6uXEfYDKLVfoiM0IWdRi2ReARm1f3V8a2lUYLkBhHi1+B+It9MoGT
T5vgp54zV/3uJr4upF8DolXNAlnfwMASoo0GM9Wy37m1MI9uu6KVtXi2VnA1XJt8qqCceb363vRd
dJzqI5iTcWoI8bBRuy/T9gLn50KaIxOct7mGud24P0FtN/g1SyeiN4iIQqZFJvNigWE4CcpUi2ly
zqVWRSDH36H8ZQFX0hBNLcpOgg3GIWNvPPJIpsDt9Z4enTyd5pv8cXixdhSX6/AV2tO5No1UN4Tp
QE/x/1jckH+uLSE+MV9UA5TQK9URI3GdnS6dgL2VQI2LUVw6bCbR0VTSmY6BXFyxInIwyIotmZfy
w1Feq1eMAr6G1U86NHbwpjnlNOzSmzsHNqINftmGRE0bY/vh8vKYo2NoTurDQDWv3+hzw+9UR/Hh
64u+tT7Jro1d2bJI9nL9NRXv7wMFGUoyduL+lt+VGLOM2PmlnAwzBsZ0BgV0sP6mrHlpmfRQiBYA
7o6l1wMdPqpH/eD2XU1Gnn1NVEH6vXxa7ZrvyH7bSYadx2NNcD2TesZt96dWwHJBxIWqjFbDlgxM
daniJEazd05DFPgs9mmXbsZlXs2MoLyPaeClQ17+aD7X3ie6NMv9GhoFKDcPvQNa3HA0hAxD1nIP
BJpxobUHozGZ4Ma9ihqLX1i3YfuTJ41Iv3GHe14y9TT0YOcNEYMRU9aPOzi0EhaarUw8BvsiMDzB
J6wTcutDPOhIFFxCbHkHo6loNVt9KQ7l1/nn6L8kI9rwo/ujCO1xIXo6VV+ztHqjJHAe6nIk7Zgz
gYZDOOBx05g7aa7RDfgzvw96Sx8FCoatNFIH7ktyyNyJYA1DA1jDby9cMsvxn4IWbvIEB16Ep/aj
HcUjhUh7k2Ob9eUuS1MFd4v42ScG5wv4lFFYvc9Qb70m4zdO5MsxJzAMP+rpgdbDxv/xUmMIPd2U
XgZfOfmEb8xf/j3FtOBJc9anwwh1rp9NkaKRe9FvYGIgzXOnRKgdFaqtT0AMsInyfCebVRAbsz+D
m92e1UbEWCBn231hDhlgAVw0qgiCfxGh11jm67bqBZHmqQf4hqSDfgFtLWTP3WdxXaRAAd1aYFq7
rSECnqi3vRgaQbkYbB0q/aQL5xUnIqLZxVRvSFoCLgjqSk4ZQdw+AzqFkiVW2FSFq5SjnPfXMfxr
8CEDOE0lrq021pqMQd1Cf6UZJoAtkjHyu0SaHje2hPUbKI5X8LAZHnnuLQhSVl6uoJ07x7FhwZqS
MGMjpSH0YgotRJlUIacrJo8yzCtOY4EJDw3u1rAC4j23XJARMgTzRb6s+v3q7x7mNM8CpuTPADhl
boAGs8B8sjEBoWnpQ9nN93YsUSUpON55ovN2HINtww06/zrT1a8ATCwC9cAomn5/slcSzXlvZhAQ
4oVJj5QyyorWf2fUQilQRTfGSGdA6X7yjlwnAri3mdW43FhFcAJTEh3dE8BWXV9yUwckhnb36uij
UZeOV0luXUvlz3wWIUxINsRI6O3Z9EuczEPUybXPlO7bB+0km5DSTdFUp0McIn+id1dLCrrvpgmJ
fHFRz4RxvZzAIfuvDoc1tKq5/CIVcQTDLVT6lzLxPwWCoMMk/KZEp3CCRKJ9zwVSq/a8EikJRzTM
pHrMPitS2Y7/3YQ47ThS4++JpbYwHTsBTGEqVNU/O907ZB3u/uVuLsM0EYsr2BnNiZ7sje+NR0ow
WIubSQtIJamRR3bTI4+MYM/E3D6cFzFbRJaP2d/1DKBnRBeEdtZURmQgFynR4+9reh8ahmrbF4fh
qZsNSwmn3mp2ELVl72WY5uROR0zi4VoYT4TpKMvFJ3JF7NaW777yDJnxV2F+N1WZnHGEkaZkz3bm
IuihyuQ635iw572zqOd2aej52012MGcI3rEK5y9BLl+1fbkfwepqw7vJit5xrEpt6OuIrd0hf0DV
weKi5lqdogrHiP/DR7g6zHHvwiucDV7gGvv/QupiEleUu3Ey1PzUrmRRRwKIreAyRFyF0NVoDE6d
hAe0dtAhn79oe8aSYMXstYO8vBN1ppxbOqF3NRkK8CgM+uBWUddiL/ICfD3fNokcQ2iss8A/DC03
l6CVL+kXwUS3cyyBO7oOMPXFCimgr5/xRzenImIII5krjHHcRBW8fGlsdeN1++6rF+kYlCAbMuI+
89nFFqD0oUzAkxCBnz+MdwtXOd78fzZ6JBEhQekzKzF+oBIcQnbc5aFRQorLpTHmLRaE2OHwALG9
Aa5IAh9hb0VUGDZKmUxj81+kJysE6D+L9lb16Y1dsBn9qpyrBi/8yN5Js/4MVgznFp8LWT+FCRgh
8r+mcKTtfoV+DW4Zk7iLFs+QVUVcQwY6w0DhyRJ2tprTQep9M3nvQg9i3z44rDYsfyDGLJee6H6u
w77MGThREim2YyNUn+b/Ud7Ry5kEfmOxXGeTM5hWleoWtkoyoJFjiU53pzg/rsqKnpJywZ+5Q3FE
AlJUOSXEd9ehTCkH0tfgmPOI4PRosq9udEiHMbz/iW5HdIr/oF1VP7Rj1ZHNlB23fGJfqTPNYCCb
IOZMv9br0r3CYQt2MPJHATCb+VCRYZkWyvPJeMf5i5jMyERsKK1pG9bmrnoBL4EM7OgNFUSLLHq/
0UTkpoqVyU9rRE7VUN9cg92v4IJD0QLBidlhVaS67vwypk+UT9/fH5+0Ovy/MJTS6UOvYS11S31Y
G81M8HzX4vwue/W+Lfdvudgbd8EaABgaKPKKiwVXsncceluVD7S2mrHzvBAlBS5nHl8XNO7NKZJ+
fEr4ouAzf5iyUg5pwxxckExMTKjRiX3NIj7iL8KBYwUCNq/WdoIibJ7HVDTVwekNaGyWW6bT7duW
RLdcCVXM9CPpc1+uTQKYaNuG/v8Fi1V97ikz8kZZE9t4zldFJWzm1S6D50/1Svfxlfnni4DxiqDq
a2TegiZB1VnFD6OHR4e964trVnmv0s43F4wa3VhdYoNA8h7SKGW6i5d8V1vYmyLg1LNB2dYlnZsQ
AssIJ4085gGyDWiL1Bti7tgZwHUQ5PUjK/MWaX9wwb0QHnhhaefmcVSmUb2uaPDXEYgOXeUSsN4y
wFU72mVERJ5B35jGoECv+SrIOgb5rQy7VrRWsQrO73g30GRDsuvOKYyXvB/1LO+GfUAhFqZ2gZGn
7Z3vuWq4QxQ5+2W/F7DUORPxt9LvMB8L4+5lRdVWlNA0ofCEU0oOReUhMGYnDmoA8Oaqd6thPtVz
8ddGaD2G6XxNIzpl8Yk1jWFLIV+bMOQabtMpRhabhrxPx0qgfdpw+uTGGxKAI/bue1A3hhMtgIcd
m3G7s6OcyP64ubvHD8WogJJmZQT9/RIa/sZy+MQ7Hgv6hdbVZYXgL53WeOAz7JL54HNDyPVQdo2a
L2G67LTo+Mr8PdcIBCgx+T8ikYys15i/UYR3Z0CnLABpGZrSddeEm1ZDZvueS5GagaUTOsXyp5Rp
XOzSdgWP0mlbsbRHhA3lBuHY8iyZoXfEX4RbGdesGfePSRUvbBA2hZ+M3xHoyIlbKoFzEEluD2pX
pDKRger+p/GC0wKQSpmvuaLeZxdG7SpfaBgJ6OyNHHtMYB0hrQTEpu/2GRDSlNkfji6wUGS8cpfX
yRyUyxNHqEYyCCjulUR+0b5eWsmxN7Bu2jzEXXZc9Ao+fcdrHP8/xrM/m+3yQCDSUtTSGs5EcmpX
nQOZa008RSZwQNpVZ9zTtBek71IcDHJmRLlI1TxA8fcRtJpSAK9DXa7BwjI1GNt2JGeUi6NBz+BA
XMDQZqeHs0NXoqZvdqUuP0pwH1R7oDK4/tgoAu3IMIXC8q7NHu1zeiwdVcVO1KoOCSG7lmpXd3At
zO24b3E+b7pssz/QhHeRQOrACxZ0amMTi5hGA4IdV2AXmNRQ2jfFpZSoSYjSXvpKi4xtbuDdEltU
ijKHUT0ms31Fixm8sMU4i1Zi558sz8GwJSqkjX+sFaoXgqUSD++t0cBpyeqM9er4jxD/lhkVQ2RU
ETCZBI618vP2vhKGE/TKwN69Hl4twNQAKw5paamnrtn5HD9nnEkotRkEGBdugzSxqzCkv5eZvSu9
Qsjdumoh0rrQIHFaz8wGIkWu5gnHYSuxAdDz0h4XaBSyHvGRI0weBfKoYPFKUO+v/NYes5SqQEFY
+JL+SQikfBozQMM3WLh8XVXCPNrFV6HOlhiLSZt0qkaq+dSDK2V1g8OO/kQIl31NYXakAoA65QLd
1552v+w1czBY95d3Kxkq36SmgjA7gzKzleEam10rlguWnO2JRnbIQ4fC2P3ERsM1eRA6t6ZMjb+3
sdEscGUOy6QN45Mb9KB3E6snbEEj/BcijZI8jkSbSr4DK8IqpbiqGe/QdZJ/xqdHdH4tVm/OJgzy
/a1QZqwJ+LVNaG/hz7XPkdM3Dp2tVim0/bEjzPjAid6jiOEYwl4TwONIl2FEUCFEksAvSKpNlPS7
JiFUMuYbhbpejLPkZPN6EXOw2/fvtsfs3biqZ1dCDYEXlLh26jNT8v3X1ZOo8JhTtb4CczEmipcX
x/Vl23Vf+bNcZw1A1OaFbUeJwriXuTy0QeVbtmBIOK47+wns5Nnjwzs7F8aIDb6wAlCXzR/Dorm1
rdDVVrSfbRgdSSmubxlu40QcWp6Jw8UIcnSEjCZUKt1KGEGJ/iLPi1v1Dz+rxfc4qr8LllLWKGhe
YLLM2kvlrBBL0FiMhy0Enh0lTcubaGWLu5cx6Zi5G+oj4XA+aJl3LwBtOSGiAAkscAnUusjINQGw
Zfg9NQdd/piLeoP8QF3imr4cD/cI54dVqpanVYL3umRInvrrJoTClzM9xkt4Qe9O2qZB5IZORZU2
RSfHtMUrO48TSNuSOU044fcQt9ux0jGuqhptr/TksPaowwXG+yOOIj54EdRhNMfre3egBY3lkKR5
todyOe7WLOIuvDHaHJaPkcJ+ennQHLJ9cnSeYe0cWy0dYGb3Otqc8YDylxJQ970Vj4BhbVU0sftz
hkNtt9tgtfwZ8P+OCtzofwG/zNPXDOKih/mH+86LUZu6t3vf/jGlWoStOWkfhjG2M9Qd/br9MLIn
iHvdoY0WITje4anj4hNNoSiH1ochB1InDt96KhzXKrPe5SoI52TTTXUeyZC736NATpefW/diA9C0
s1Lnbj3zCrA6QsQDzZMMnsEyZ0DmTGu+HEoPH2EGPmjkJCMWASA44x5+GDNMDGFU6ffs8jyDLfYC
PJ6uMIeKot9fvkuaKWcwZ9XDaueFON7r9hpqa3jxc9nl3ysAz5Am+zujBy7NUjAzIT77xJofCuDE
RIIzUPgijOz0XerC6RwuhZmBksiVCNYnegVUDVOoX6YfZCOWqixFozBCmPM0v9iDwNw7h8450IqK
qYhXdmjt0GNgwQ6oWLuLiPC7RCCY/jbXhEdRVY+nhKFUcL7DbreAOsZsNzqkruyyQPhOJs1/wkDl
HuSPk8wWz08Xfv9NxIl0vDWUWC9C2B4wZBA7dKXZT5uKJRjvmCBneALsvxGmXfm3wFnvXGHhJW7t
q67PO9ruXiso12dl4tfcbFkBgOS4cdtMmihfwFqsjFNZfeS42adDK9wLGdIb78i9NgLvQsBANsib
ZcuUMaJMeSAx55L7I+7BYlYdj9Dvs+mMjZ5nGQO9vtbNQXceraVORDxrDTQHdrTJjJrQn3aIC0Ya
Ai4dWz2tXoYrtYai5Wa1DtxiTKkFXQjkf3PX26MYP6C0l8a55ixeZ9g0F5BvBQeSAqXTEV+gRQBK
njV3iE4rrF7ZvmCqThdo6333AgIrz6fhdDvKlU5n+mz1UxVSWA+1g1gz0hT6jvxWp85Z3rqCGDgw
ABRUd6gR+o7e3st11h7Ll1t5YO4o+l8h/eH3/lttVBlIAo7tu/R30PvJY0VVjwv+0q/M9IF4Y2vE
NXhy/Jz3VaNM25gTPPgTllx77P5mOVo+KG8CQKSmu+gcFRO8Zgkt+S8gh8nuD03GspYwWFEIaafu
vLuvztf7YPzMSArSiNIZtzIwwzBeB3tZWqKcNgFrL6BIonq7d6GrkPJXHNMFQgVY6GvVpgZeK9Z6
CdNL96HGQdY4UfJqpU+VhB5tYpCWtPMAVujNPW8Q5WC7VRXTn2U74yLp+othki6k1Y4Ih9ddS3K6
RxdZzOTFbUZQtxQ+oASBwI0wExcqk7H+s4WtGG+KVJ6P1teTyFJFZtdJNuS/IbZ076/WENH3Y7ed
woObCMKX/ZP7D3WMoQ5k8bSMu14FWNlI+vH2ciPLkza2dL8QDYnJE+C51LnThQLBzgiwE8MoV2Ju
E881dahGO46I7r10YNhhRtP1PLVhbBltZdaNWd72EjLUjN4RT14qm92IG67Bsh9n0eWyJ+VRC4cE
wS2xERoFkeV9UEG1Tqa2FWq8l7dtUefj30WOlK5WbsHIKmib7uBY+hkOZ0TY+HwfECiXKpORo4Qp
d0Dh5Yu5k/6qnKuaOW9CrXu7qJgH72jNutMDiTMFfTSPerDbkYM35R873DdihNjtGjSE8CTs6P+Z
RFpki54XSGib71vHaelvvEJTLS170PgEjTlsciUedIyJRDGIYD1HMOBoZ54zQdS+HLgQistDSFDq
i2sgXKroHP4qqc0zl189v2nwjPoeai/ewaDWj5OOey2ninmq5vssrrzSBZouiu5pjgcRE29lsbQH
D+EJ5ed5m2VzNVAQ+gR23gDY4ut3fgxFa4+uf67bBmmGgy+TiR0UCCAPSSudVsRargJh5IhFMUPp
zNi6IAfmb/W3yzyXP/fWL4bsitwSbKWvSJ2MDdB6b4ClTSGR0X+CBrTMMOG4Bs86/QMPEKKKCmio
mxUXQ6EEeKEhdzXfN5eHE/j4jfYaKwY2Pd3a7sO7qvzGOPztGLXe/AQTtTu/DbPvSoxs6WKt0ApQ
Bh5YI1vd5YR5xC/bOlW7MQe2xN9xxJ7SDf/kDxTqM0gSzs0PNz1WnERo2yC8yGEPLCFgryENXTAc
BqqC8/2l06EDkjmW0VIvtCIvzYtvQBqM3IHeqJdgYzDHCRVj7+YuISJKNeoh+ISp+f81p2lKyYDd
LMkpTc0sQJYH1K8EL2/3oTzbo+Fmmh2tCJLOng0Ya/ZY2DnZtjygKRWdye33unN619yTgN2lNrpI
R54m4MEKYChXtjTsOtPR2N9WhFpDqPFGXy8T0SBTNL4lj+hS6Hz89p2Vsf1lTlhGWwMfCQRkO4/z
3C6AtaOwtOsK212lUT/eCzYVuLEncv2td5sfe9TIi2dw3A7lMLpPtEC5iu6N+evg7N9ILDSVQ81r
VbzWzgg2mLcydAkV7mUDETFRYXa05y1BToXBqjdIa1MNEmXr9pp6vVY8RzDW55OMRGnhLpDHBr/H
0exldSaxB5GJdLyfvwfLkzm3vVUhSaabKHk/wpbnFFPKJfsIHLEQDSfTg+WsJNaeukn4N356NDzM
BoE9Pj6eZCd0q3tsnMWft5JRC1xekPLDic4p2JiJSD0s9JUYgpK6ohoSVsR5/ZSF4XbDu4a4slyl
DhcuyiIj+Dy0+R/92DB0TG+iwGs9RRAxNhSO0QigqZfkiSGsfWbxrPY1RftQxZp9RtN278aw/8Oc
y3DZ16gehsTJX51mZ1wdQ6F6mjXTzIq8OpVJRLX42DHwA/VMp1NJhopAfgGinCzMVRIMNo5lmrk5
qhBxU9DKTff5CcPe6EicwNQdeu8Xx2Qzsf8JFY9EZEmtY72xPj9R7UJ/z9jA+qoM/gKgWIKNzJ7l
dpyPIvNwBBjrDtAjsUMUyvPsrj7E3AIEm0Et1ZMJhnvWE/fae6GNwdfMbCbqS/+Hkeo7h1YZEdRH
aJ4VxQeM6Cn4+5iKon6ub6KlwuYTaH0QuTzdStPO18yAoq+8is9lO+b896JbeFr1hk9c6/mPeQWc
vSVs39KjtEcNlCkFOAoOW7i2nSjA5XHJ8mrccBJB08OTSi7bBHIK1eSLk5fHLgPJ6dC4qa+cX6Sw
UHEbwnMt9ETn8eilk3PQcnE2GA/qTVANzBaLKDi2UaDbpdSBjqbU+P+2uKvZrKb4JTBVdOIhREt7
vPPi8eS1/OPjg948+KAWn+eetWDF49N/N6eu1AFYhkfJ71e0aWSZBkimGlSB9g7CC6abDLYMSDEo
dOYc6vjikbTmacGlklhcWePsKBbtKvpK1DpidhKJVWOszMSjEAy0tRbCl2XRaUE3YuRckgfsO6rl
hqeOROapTXHQFAyw3KkJSg/IPEE64H31MUpbuz5D+s7XnmicKt6lpj1u9C+wxIh3rt1LMYjfnM5z
JXkfVoWDPEfmUgmknpgeSfs1BW5RWn4p64smGirpOUwebAPevthy/4od2gyB8Wz4DBkeZ65HwFaO
oaYC6GdJcGi7oXvD4rlFgMaParNBwhoqdzpxyq6PzPwN1ObxMycbiqVj8MHEfLagl3D9NOPhDzGQ
uZ4wI0zlXwYgjIrEr5VwggVz1pYi4f1vS13V9sFImDlf8NU+Vi+7Nhlwag55UA7P5hGD5XRkUHLv
eNIkmY/JueRF3Dz1wR+JJDl2lNyfrdUdnf8Ot0Ze7rJtxJ/9ybje01I9DCu18UW9hxESHy+Ca7gv
W4n5dXXSoh/WBJUqyIaicjMQWSpLC1yRn2BirFWmg5kzLDyudK/C46qvifUukshSFimhyDUFxsS0
zp2/JkUdA//myvRFEsw2yHCq809M2F7Mff1528hCURevkVe/VaTRLZ5RFOf5JrAQftYLbi9o/7N8
III50CzZ6pbH/0kzRuFWrmAhKOElhoEsWY4Ut3wvoMyesOm2IHu6xUMdgKxPmvW7nINcI06Ax7HQ
k0exNvnC3BBp8vqCLoljobRa0fHx+edze5V6lTMXAHhsmsidblxulbpQ/QZwyGscGOjCZ+s4WsJ/
o8uFMOdj//soDl/8q4Dc6ljM+Nlbe4ReItcwTB0cLH1GkVdhUDtndSQ6JqdOay8V4Zzf7PYI+1MI
hdJz7qRtGmZi3/IfFXXzmLm+ZWvrZ5c1kcOgTySeq343uGB+weAmVNCp/D6zYLe4bRwl9TZ8vFf1
fn6HIptmbWCIpIHW5rm3ZZ2GQAIVWtUZ8jbfROvtTp5GO7HzQE2Fz7XQvzuWHLwhq2P56VAXt7oW
kK9orwpbjnNIQ7z+OMjHKgQ8ObGnSJ2TS7+yDIez0D0axnmiiBultFpqxTQb0CUXOxy130lTtwV+
H/eA7ucUgpd08K50Ej+zsLo6cvMnX5lZWQ1bmQdK1otP3YsEMwPmWMYGAeSlw+6FVHUQNkqPIOVM
00d6JMqOpK1LihkqVCiO15jiWqk7C7Dr7Xv60S0EYdgJhkK3X0p0AGrtAyBxecLFVPscGn1H6Ago
8NkPBjp3oH24ms/BuLzKLSivI1BB/7oBfoPihpUTwwgL6iIiF91NR/eSPnG2zpPWXtrDxK1bV+jF
+Tf1og4alujgcbRokI/1HYUyJUFNaBHAIlkrjkPvcCN/Mq6sUJWxFo5w4T1mlx146F3tzoJ4YuXB
mA+xuYne+znT5KBb3Am8/8rKXqIgzoK2MgK8wdV6RhMolnMUX8UN9at909jTUDVRjb0ur0AMguCm
0rSUh0I7FnNY1gybq0UBqtVQ8oU9vCJqzixdJ/B0IQNtP86udy8yigCysxPhnHoTrNsFwKdW4cxn
kDtHi2cxJDBbC3TmAa7l09GWzYN5Yj82NdHeygyyZ2IYcN/IKztEcpbuB1XkA2U7pZHOLB4dmQ2i
Hlg33G5He51/LG4dn1xbh3e6yfTeGSMk2gt5gN4dC3hTjLT0gH05Eg6Xgbi3fNHXF3559XTkufR6
aVbS46dvrtXdTJzPNwTwTob8toe77bKLFFx1No/DR+41x/SKikhtuvZ4iBGGYHGsOGAYSeGEmdrC
KI/PqzMKZfrEVgnxvZ7eSqAiQ+fYOIJ23+jcm25po50Vk4iaGNvkoMl7sA70yBe6kgQWOIE53ZnN
uc/12emtDM0VAWsYHNabFqFI0ECGC0ZV2VZdUIHdcyu4DU7yhUW5bxpCs66vk1BoHZXpVrWhU9G8
eaCIiisHP833GPmTQboPtJO2se8bOhE4eF0L6jLj7KKZvhXwc1zbtFTzYcAFW2+GIj7/NdTN/z3M
+F6oI3Tra4aXnIJ10Ndl1ik8TQRK9b9A1aDgFmlVksuFS7C7mUY3hJnWVZgxwR18KLdLm+J6QB5y
9Anr8R9waE0CJ4VCv3WXq5L1iX28cIQ4GrKWcU/ppsuF0RHoRy4nmxDhp4iwpsCh3z3scgr2EcM2
dEhQkus3kJ48AcQLm5w4EWx05V6ynsedCHcwcM8Ve/1HgQ2I1q/H7y9myPO7dSFKs+acXXerI6cn
w4ld/KSGrPX+WAVv3gWXYBswj+A6gkSwub9UpO6Juaiaa4eUPIbAVHzS4qIQrfYdGHWa68X8jNL7
9DaaHwjgwx5RgjBypsdfmQeiZGX/VT4FSaHj0nnCgwSV68DjXtg6euIbyv3r5KtOuiTheTiAjaC1
GdZ0xzJeNtgZIiaa0i39q2Lc6oIXe48YRDzuo20gJDL9uXmz4utGiaTLb+X2tbYZJvIzX+bUnIRw
NP6SSJxRssQ32sFYB2bYvfJieD4brB9IF3IYkxPM8CPBKrCRLTMwasgMmIuMZ9dLS4suirAZ1s//
oOtLedmtnbB9xVih0Op3w2AoQw/waQaRUFOsmaHD/2OIJFyvtCD/F7EcfwYG93eYURPnWOYlrM9T
O05NrppedzWvd5W3DJb07OuL/BDyaqhv//jcAMtXX+dk3A8Jb6JxN5MW1bkqvgBpmolTW2hJDdWi
pq8Qj/xAfEvR5G/IzfHogg3VxJZLN/Zwwqc5769F8WbDSv6u/yKgaMx0wqyt6LFT/eVMsHiQfmqV
cQSj220zBRg5B8L4ACnZBkJNNoPZJLcEa2FTmW72WKNgVn5gsaMA11oZD3xpsr9IsUzDn4TZ43CI
xzE7tUvdmBcSXXR3urFPgD0ouMA7gNgtTxIt22uWW/2IlboqvboNh8I4jNz634K+6NNTFYakB1Wf
0FIbdMxkvIHYR4x62Ir6n7rHiP8gYwoN1wgQ+rwMlP53Vb5K8HGwf8nw3nZuV58sUazbFdN1QKM1
yNMJuvLpQzU85HIbvFMvRnVbfu6c6oyRIp9bLyNtxPECZ6uqfmutFwHEMyc43CHuG/rycz4jtW8c
sFplTzEOH3U2o5qU+3tpUJTcSTypGKv8R2ieLJ2+kEgn4+LM4T3HTOR44GU01lsvbiywkDXINTnF
+odMM0PmusOCc9hvKmmE39tlYvZjAorhW7x82UNWs26YeK7mZWj8v2QXVmiwQkIAzzEUmD2GIk5r
xJGXlBAl3KNXfxwzgNX6DZF+eOP+eM2Xu62aQp+8h/jGGU8rVof47a3y4umhEL/RKvu1r/ypeUEw
DV8FUbaFcg5fbS4D775CilgP0YYM+0fYW/rvQ0x4qljzXbBOGt2ygudmB0hI3c/J1xPbh0H0TunD
96+pjyXaAy4obNYEtk6RJv14dGPjtiobCmHvcEvlmh8qcTr3rKMVDldqJ+gh+I+gjGPmEokZf5vT
xrI55ht/yMxEytkBVzTYl8LKBZAohTsdfoOooz3Mjm91QwDHePTGyqiddgMvqqaW95YlN7p2s7B4
nikJIDBNwYGThUHoeGmvDvolmyD1HWDFlPvYjYI3yrLD2n4NRcU42aidblmOm7q/48lCcUCquxUE
HdeiDqm/hO/WL7ZKX3xREBasOnTinZPzMdbQxitg8YhqLNDUqTA+WP640kG7b25h/l+QH7i3FA+e
c0JGKtSuiUu1jxRDeRgY6J3dHxoshHcUCkv6ahqK+IeV1r5cxGpxBX6kJuw5gjdvi/WbP1y2pg32
OjOJUH2/AnzEFET/zvPwRZuxPfpiz+OMfonqSsvx5M3gensYa0WIH3I+5DA43aDgISg72zIeqRML
9re028qxl28oUvt3Al3dZRE6jb3qF4GXJEwH1dc6lbXMydlgnybQPxKMn+9u0GyKtJpQXHLclWRH
hjzHSphUIReO/zWZPFOR9GTykfca5F57oS8obJMxWA2WtqYDyUyVpT1Y15kHeUtoSyLE8JeE3Crv
+nIxRlkYrw6wKi4FIRQP+gyw6l33GH8ptMvdZmMnnrELNQ7a7/bo9nHnR+0lPSCHcY8la7SK3qMk
SoKx33qEE7de6/RHCCJ/cZKhYfTwcR3YeSOUGiC/sgmAkrGxTAbSoIcSuf24O+LzEYL09oXJExgG
iInwvz1QnW0XB7jwzWvz11YmJobA0c1mFYp/O0KHMDd4aK5rRJx7NRbEJCN8MPelAxlswj/+2P9B
tVMmYabVS7+V+/GCDAkpp1tfwAUmZ6LPD/KF7ExuN4cKOxklzwaaj8TQt9LE/t30XUukwhQx6B7Z
elT9zUUHECKMI5cDzqcDfNxGyIPWg4e+n+OdDlzD/Q+2+GQ6nEb/KMvJL9RXsK26hAVhDqaplAfA
ZHJtR4SX0UVWjOBNrBecxFdodDLryRJ9nuhCjhjHus+hweet2sakdEU+iP8tnb0PwkpkhFHUzz7Q
dAlxLYv5pFb0lXeWGeNfl2ALYKoHbVkQCw9YqiiS0zfxIW+mFa8vSeY6yoeYqyLxmrjZnvwesmu0
w+U4DVAWbMXMSOSqD8jhNpfPATd/tZ6zxIVImW9kWTGUw8dJDKd+SY4rRkk7m61R8k9D/ciq5z2J
UntwDGf3K+9LeBcI+r9SBoCWU5qf4r9XDCO1sayOaaI6HhnA4iol/ZkbFrsdSPotrLbjrjyE8Otz
tcFVlH/vTaWw0XyL5/4e7M6VTloZZZxRCs39HAKjhq5DbxpPcwyWsFGfYo8AZ4GoJ0FVahnL+OzD
/anD1GZUyDHdO4G1KPRqKDxPf7r/EsDSvXcUJrZmZMyD+Pf2vwn1ifKAhyMovuVap8QkPRFpAVcT
H6TjZDbFUK3+Ky9DQGPIiQGylgBPwrrW1BwiFJT4KtcIVeKYkel6QVJEI5vHmEt1FSfDrqOk3/uA
VGvjJOQR4quy2HVJhxSkQfyoaoKss0VFaz+vGGFjK420g466Wwq5rlmvK5k6sIEyJd+fGS6FARXT
SszrUR4x1XS34Odm0nV0rqLs1ZHax8fvht1ui+HjN8BZqJWeikgZvsITPBfxokyF3R68XiJYO5kF
iCmEF6ycQ5vIhKL1pQ34Ew1xk4ok8fRDW9n2s/7pUzRiQXNdNOI+M77VScMaQ3BbtCZSHuDnjObc
Wdj1uw05CI7xLYFZGiMEtTZB66A+Vz/1kvH7oHH/fvBrYSUDzX4STnllCHct4H5sgKxE9LbpMw6s
jzP6FpGa4NAYpRXeksMHFApKaDCe1n0+WNLjSPpLBmXc94glfdFQ2Kry8VZn0JW+Wy+tNGESqzuE
U0fQlyJiEN6oq35T4ECxC4jYU5bXyfhPa1fDzF57jQu5SqbZt5wilWyfDv9RFqHnDkPQJSLhobx4
HefQ7Omt9XkdT5pioTYU9fLtEUIUguOfArpK3ZcDRfZ6ji51wCazJ0GTZtcu9EOcgHUp+KGuzT/2
XJ+V8HKf/9iipReo+hpBG5x03aabsXDDz4ic7LaHyD/g3p7ngAtXqFROuRHE9Ur+KYXlJ6gVxRm5
SlBZFZZV3Vvm/3851bIaaQjreIKJghDJe8QVAo2gnlbyWITSPCMWjrz5kSXTDJm4n6NqAnfslyz8
TXSRxa4s1NrbzfTl0/+o5f+zc+NWKt9mrsDxkdJMNygFsR0gAb1w0p5dY7ZPJssHzuvTVsjTAphe
6yxbFHr3PMrEYYuqsNsgCKTO+DunYFmERCZaiQ101ofbbSolvnfYRI8yw0HSPqzVThPX9PUyzunT
1/6hVGK2rR2kCXN7bwgu2Z3WVcfBLIBWlmBhEald/HAUe2DLNh59FxWgqdnwB/XOnJW9/iZvrZ3q
jvsz8C0zgYrYSR/Qa2zTFsMV6fOjVKDAtOtNYFq6Vm5WxW3TA1aCSNQT1bKTsFheT2ndQ7T6/aPl
CeROEIEmx4ikrWaFB4D7W+2qWm79Z86zM9FDZOtEOnyrnCVSlF6Gp121xewYk2ZCx5iwNwmnyKLx
ybEoYfljn038DAidkJalm6fN9nC/uw4HH/qbUSSaFGHb3yueM4BRb0QLJg1EgwHSphNrkUAopS85
g4NiexLUaEYjD7BDX1LHNYy6Rhb5Ea8qKuKH7xyeoxoKdJwboI2g1rTC/sJFR5nTAUj9fqB9lFll
iKMM1GnW4pNWJCP65w+AVqzcAn1ZXRGAhy2NsSJ7LTcGRBSoIX/4hii2sJyXSwcLkIgi1iet4NhS
ZPcbhAbTSJsnQAaRDexFNjGSKo4qv7GnZDxkwayANnzOu1w7USIHD8+CWDvkesnhOlb+6sJtRZzc
rHxquJTNxY3q7KuwsZ5Oo2bo7E0HplEEFJHa0U1adKBv//2XlFi8Zp8DQV5x3DWpnbNJG8E8Co4x
MXBUy9wyJGxyoJlHjtZTk1Ui0uflOJXib2qbPJJDqaYqsSGiaJFi8NuWe7B6HuiFxHyBZ21mXOpJ
8AEQJSLsxCjjFqCpYYVEGQr8KyoX1B71E9hIN/WfrlJ2XZ2Y9ekQG3nXMjeWXd3GfD99lYA1k7mZ
3AinwW5yglrcBm2nyqiKGwalPozYXZY8UFKV86t7/gu7jdgcn4VB/alg3+k8PAmDSRt8ZJak7uw5
7cOmui4tuP7/Gib44rle1QEJwKuRuRHpZw+kdzGxGlOQt/73zxdNxndSX9twZXIGCwLX/jyIQIJ6
0S3momIDgjmZnyFpPO6PmI3Q4zNT/aE6fE2XRyOTJ1MR3Uu3mvPbSts9CzwHeMgDQonTaJdRCrQ2
wm+mscFfnoaLAwdyN8EzFrDkuWLjXrNVV9eR4Nfay0LrrLXyNLnRy8IKQYCFYmdIX6SM84VHTgg3
mkS0LTII5vj2Y+nYTXqF6S7/k/n8B2oMcSI0MuQqXAhha2G1cxSc+Htv18m4YcixFlkv+SDIQmCY
fmJs41iCv28UNRu+P4ZJ0hTHgKyC0xk3p+XQQ0qOkJpAexNvYMzNZRQYuEOO8j5heI/dczKuBhJc
BgJLG9yA0VBEVIn9htPRjD6NnZpa1umLxiT6mfOZiLBt6miouq5QJdZTuoV2qTJYN0UVVoEBjnB9
A8PWuP8fVEGXm1713NmEXcZ6uVbcyVAVjQp8SE8rjmf3Bi/b0KnbpeN8hfqw3qLHCrG2J9GxR68Y
8t6qQ8MiHkQzC4HLO47ZaG+y1lkGTGxvsLy+KJLD+U7awcgtmCOGQ8/ki9Af6gHrC+LoDuHPrzB1
LRFFmj83F8cmdVT+QgrpUETI2VPjqsOHOV5pQSBY1uDJYGsblXuPoO8byex0GkkBvHGLP9EWX5Ed
yod2VZbX8IITkK6qpOdybH08R2mdifm7VPjfQxwDJ3MILTgvmntYEJfD3weT6/iGqFFPAuJ69OSX
ja2sZ74bWv+k0U6cvLIWjWkwP7Cys8DKS3BOj+mff8K18+hQPQZ2CdNoYw6i3jwH0kD/eAYFvuqp
ONS+W+9YUpxCtY9hveoj67DRrC+gLS9EkAUmbE7bVbwmxuwpzO3LYotVtj+aPKlG/XQBmoNulSvp
SxIsHcshE2SwEjowKsEGV6nu3RRvEjhbpvq6yQwIwXsAIvme74ZwILqCGXOBT7zSCxJUG5EIY/Ks
4FEWF8t2czzddxjNctYPTokmEXO2qEVYJrNKDJbCE1MzNPCveGfK+SfyKA+wFMD8mGt7ydMPAgVS
BVnlxpKfd71QtWUEgsmKVgnKGf1ybNpXDMCFy7skR3g83avbgrCvoQVdrJ/G1Ptgr7vuJgHm/oz+
u7AJdPQAdAF6osx1saT7SmrE4ihT8CiOHBmgIB9+TUhaGa7GSahOHXiCZNxO6V4J7t/OXxRR0inP
sGS3yJ+idGbSSsQnibe6YSWxv79+jmrWT1WQkhStRwtkAz5+8VQ/VZGJid4AutQHmAKOhJsNx89j
JMEBrENr9BBc+zTlK8QI8qSE3fKSGQ8C524AjSR1dFV6QsJKg56YRoglNwz+VtYYmfRrq1Ra1xNJ
vkSid/zld1LAwCDQeWd/iyCCSv3F+bPKMRsAl5qwTQoW7l0pfjAHIPHXjTlc6Art8RK3mAqBAKmn
QslwGSE1EMYDuhj0JYDv1+L0RYRN52xu0gwWZS8s8zRWUaP3pNq+YlezsduwnUJJxRRtiO50T5sR
WoZcnAS3CQD7sYZvkVsZhuehOVL9HfoszpiRVgjuITC65FnOBvKnADg0TKb+eanGjBX+RcPaQyMu
pbo2KbetpD3x88U58LcUob5FvCprTk2lTGO+Zdgg7nm2UqcjsNAzHjdbPVGzZ6YJc40p/Hm5dQTy
Tc3dQejk0Gkr9jJgGm8Okd1i4rS2Ju+GrResLiMkHIejdABgIO1n30Fu8CbHtLy+y2WIAt1Fjm4b
ogk+FMknEqjyEZzTWe+Ebj9ri1fJMxcamaxH+myx4+vV60qcl2STiM4423Kha0yV7QpKvAsI2TJT
7CTI0m/qn/RElHbb/eBzV3pfNK4Qf1bwdjVHkWlv0cfH9fIDzo6ZNMiECuzNhjLI/escSV22LxHg
bN6z9L12VLecmdnC3IIspiv13LA+ExUklJyhIe32eDcoszGE5RtHgPJPKAAeXmnZmk/HkSrd44Wc
1sIL+/IjGFchdZg1fLXvAyyH1HZYvo9bRYd5P2lyvcL3kNjtccdFVgQPeV8mcBO0/gOXKFUn1lmx
WVjcPkrZwmqS95ilbOKPVB0MVyNuhxE0+ToJOES0IzlqvMPVuq2cTvDsnyUEj+xMSiQhxHgXwGev
5sIuG+4Cw57ArGh8XaLX9coRAbgpK3kOoQ5P5rjN3YkXGrcVMcPXthm6XizsKggeNukZ3cAXG+lA
g+Ycd3w+s6NvmSq4U6p12zrbIU0nZoGvWfGCjh0xaD3P6ae1JyBFHQ0r1P2f4B0CsbsnWmKwnro4
vntqFo/WMfBLe+8ACEuvW2H4NB4nuJ0BuNfkSQn3ZnhFwFn/v21H03nmFOH8ep6ChuOapaLfu9Tn
luLgDILM9hZklk/ZuyYFrvVbQsctC6ALTbSs84ehov65xp2TiR0yJPfHd+5ywZuWqeIClTFew6p0
a4hMuEOMOaxtLkAH5dPSjbt05685KezQ95l+UZCPxNlboaNSGMxiaPMIRlJkjCkAzyVJZ1Fl/2v4
eWlexbhkBjZ00zEzL3bJD6OZa+CM+viWgeblZLia4gVobEK+xhpUC4uUAvWsxVUhGy00F+GyScFE
1tk/VbW2SBypo76A8ntvyHULKQ7se+7U5kScEDPu9oQ8Cbt5qyHJCGbEamh8GC8SoapSO7kJV60K
impHFRr79Jbm9awlLkL+xivUvobTW6noS951I4nZDWrfm7D0WULAKLFYgaT3H7DEjg+hTZGeImtx
fpcACYjwHJOo0hD5LKr9dKU2I2txfhgvdwFKjmcT/+nQcD2xeK5QBY3F0eVzselcyOxKHgEslcgZ
LP8DfhoDPhlmbn85xQxcXnvUS7IM4izF2GlFhs9U+r1ep3T+WZxs4BTclatFFJGyqVxnnsBLJTtj
E4pg1f7rpfXIVyipZ5amuZISobEmK3mBrY+IGSRKJSWUmdaOp/2D2Fn4P4ZDJE73AOSR/31Wtv4h
/kl2kGE+nc9MVAJKBZBVN6/Gb6O7uTJ4lMpHLbjndZK1vuSHekZzicl51UOUu6Bmrv1m6CmPqYDq
V7F+RjgXuRumxa0Iaf8A5Asw2wFJ0aonOBTmFbFxPc9VF+a4vHNgRndzuREOe1caaYKhJ8ly8jn2
p8vStad44uTRWZwcDBbUky3qu55zzI0w5UpiGYevaajZ++s/bQrLnpevh7oJg3tBsqXGtiFnbRNV
bUTyg+n90P889Sb5sDO/FMFO23IFz2M1MjCMOX+PPVnM+gaHG2hKd5yM9EHMI1vwfBz3OZ1O1G3B
7lGQWw5gtj2biIV2M7v2qWQyuloYTIHwAEprJqmxdMdie/bpVZPYsFpqY6cfmd+4Lxwb3eXukUPC
YDDz3pYUBYClWyPyJqBoUtRfiFf1LoBRXTJsMRcGos2FaEY4qM08HTd5o1h2HqIpPAB3ugJcuK5A
THkt+WqqTkHBQoccTtKJJ9KynDpBevxXlgu+uBWt9fBsdwnCllLvOw2XOL+g1gblq12RkjQVcHMJ
fUxcccZLdp2tGKthCbnzpnbOjO11gA/7GAQRDgg8Gs8TpNxXn1TneRhZP5lbVzdlm5xwg7K8R2fi
YF3OR72/35fGJn7H2zJp3SGxB/nzfQsPA/Bcty1EWeqSfL1fHbkBebZUuwZ7Z5hBm/g+1/6elRX5
u0n0bX9RTzBY8VHljsyeoxtTx0GAR3upgYq/I7aoGbvLIBLzgwh5oePfKLJ6pJLf7dXiA+2hD3QQ
joguWXs1wbCbKG2fgnRX65pOnjnMTykI+hxsmVC4TYNd8GWofv1QGjEHsl+1IR+QeOCcXssTGbPL
EyVdtRkObdE2C6AGAbv0WnbVOSpryeHytObEsVrGnxVO4UkoDv4o2CfJrIkqyyf67GRjn7LJt1qt
/q2FZbBEguurem7DcUQpS08MOCUP0FeKRD/1QhzjUPAH0XolsUKDAzaPZ5TtcT1l70m3hhAPMoTe
KMR2FbkiJBotMF8m+eSAruzcDib4vIPiQ9TyMpnh67iG91XLqnLl7O0XXhKCMva/3jeze8NI6asW
fF3ZqlVw02seodLZwd8fPHtAwJk0c+1eD9+kBUJrIE0HTWJOuI72FBckucUBEdWoSRs+XHyR9k6b
lYfxksN6y1X4P0EEF872//qvfqCdA2Kkkcr5vW7REs0Egs4joAnthA3w6QwE8n/J6upWFw5YXc3e
zi4SLXBv2VWunQjwhRjOXr/qM0rgaZ/Q0xcqIyMi/a4U+L+zR4rKD4fHCw/nhyBLqrXip3HMYfLl
IU9Uyv7mhIMmyYaZKRLrFDbJiOf7qfErUcFNz9jpdYNK0c/7NvwvrKRjGqc7ceZWgGmBU2g0hkcy
mZb6f/pKnaPbe6VjaRfW2qoI1dqZl/xDTNPFyQ9yP6FWpjsjtYxSNvBWm5xKSqjVy4bKs7u4QI67
hTobV/fKDT4Twb2XvXFIH5MT9LA+5e65W5rStNKgbkjpjcqOVEZIH2+7n3KKbTuE0jN5q1vCYGJu
RdEWvaJQ8adgKwTCOdqtfGo1GJdlyhjzNQbsauS6U3funHB0Vl2Et+9oYx6Wp6409BWXV5CifElt
TYloDo78n7CMvmAs3duvjZsFARlbA+UADPrRA+mqRVCHNW+Nm1Jla/8YG644MUwdx7ENyY5+sJlR
N9geZsuAiTMJUkRwRiox2zcovEAX4hJl2pPPtzKMvxNoWqAvagJkABf+jwj6GwKMf9JNtgx0q/+H
LsLivFb6lykB6nz6PM9W9Vu726JJnOrNWTx25gSBBZ6cGdwHYPx/weNO84JDuR91r99Vbo1f/Kgm
uctpszGwBjO7EJi43YqgjPsSFFT3femMylk/S1c7Nyvlx8Q3r4ezzOuMPz1eDmgXtWIS2TmvS2mI
Z4KTZQYvgvGHDA2DY5la9qHhnjzayq0cpyz11CA2axg8hDkkiXfYrJBT0rt3uFf97tevZtV2JzPR
Dcfl+TH2M2zRaEAfF0Sfj1yFPhQkoJMDeL5AIMcDNLBOLb3DBuwKaTABSs6iClQfBOKXin1jlolh
uue09rcErDjo49ti5+nsih63rx9tptM+R08PvoY+g+pv0WYn6rMSlPgVhYCtLnJFYx0JgnY7XxcQ
iAv9D3Hm8kYYJ/Nl3mzATbgAd8S+/nYy0gE5Pri60PaI+dfiSBJ4MDvPwAcTgPjOJoGnS6fa5D9g
hqf6rY5m6L2opNqpxlVFVXshP1LjEOiZhlL6+vLNxDO6rVHskgsURDmc5FpfZ09YdmLMf/Z1d6Mh
0s5YlfTB6yeGILFg0H4yqK9LrbeDJXet1cjzNpQt5bhjHj4kGKHsNoVYY2MrkRlJr7MC+cSTnQMz
cTtcKOaZGgxxzsLeXEcuTs+mtwVSTU84+FH5d3LN68EQSqsrSjopA2MODSsrM5v5CitaIH1Ed4fP
h/73YXhZgCZ1D5uKz3ijg5y+CPC7nejL5PTd/ErYWqalQ0OUiGVjxm8G78DhWThQB12UsnPHmV+W
buMcF+IoW98EIV6nSfNM+CYIpt2294/XzR5JwAjEB/Drk0OhkhSBC5VHKZVyHsAFke2HLBnMKsSP
ono3lET+2pDdTlcP3ggW3KyBoz7jcL8J077bI5d5JLdynKNNXDWBGkQs04yyCxwYaEOnK9GOHKLE
YDu8W6JnGleqynZcNJ3CTj+D/BgC9+E923570hGiZUd176+ZO8lm7+zSTlqRNzQC2Pd265dlEMvn
x4slSbaczas8BBp2dPb6g9WOLE6iA+4jf6naKALxhLvnR6gHLy94HB4KP6bnPn8m38RJqlqMWGlv
k6QMtESPLIsa/kYP/HfdP4fCVoA8A0GL0Ez3VUtTT1RSO29zSX+3z43uwyI7MYJfza8xh6yAJGyh
kBurMs1CcnEremyD9vWw3wIRhv1sw+Kalm5EBkdOkfsjuXfvBcmTuPPHWV9i1zD1FDLmuVoW5z2J
N146IXl3XebdZQs/6dpVZeuihzhZnyXFqPbMuJbr/mc+4+Fa/LNJ94rzbpy2viweKAvpa/enH86h
YKlB2EYiItFTXgg1xLBwSHeYQjAmHR1jEsC/Gbxg8s9oKTWdXZLgAHzrJVobzqOP+IPVLBk+HYE4
XLm63tFST9yweC2Y51qIEKi0n+A49S7gl7wKFUQyXqQn9IiwQ71NmAcZDDBo5Tus5glqTr5axZG9
FriOb6ZfKT47Ze6CA8puipyLGNgAZkzvURpWe70sh2n8d5RXoKjD8x16gcPTfI+EIN3SzLaQn5M3
E88tb3/BqNEGaxOMPcLIE+0uPzwoS0CUCyhIMEQr+F+ToaKQhrwEYpV00k0nGweuEm+zHKk/Tk2e
6ahVoNBQwn0Y8ftvkxhaeLurB6aBkxsBWc0it9yr6fsk2jPRHpj7+26nxfPtaGXRuepU46KsSpMt
r2JT7BZZZqDc523qp+Y8a85mv3ko7mzXtho5YmYxMhaGWwRIJX8KxgijDDnNFPKCN9Lyc9rYq/2M
uzRPrcQ7PksS08GJGNJ53z1xaTWu6ah7USngOQUg1N9L0ReB/uQhvpyutkmU3IrSVp9zxicpMgca
XFPuH4IeJuQef+UD/8jUp4Ez2o3eF39/wMhOY7hBApQg+0uypqCdqyJtZKOn06iqmVkqLrmfFGha
YsMJl3aWYhPjMOKywKGhP3XCJCQ64R8UlXovauPIwwDV+y6RJ96yMEFibx9ptDuU4bAJCVq1ajHO
cOy4mYyg8qXOu3DIdLyC8YXOo4QI+USRmAb4pmM1eomIiwlXFFGqiogbgrTOt8SU7CfZaCn5tyW3
pIZzAOQCa0AckgpzXAqA6bgBdp5gswSAGc9vmYrx3TB0CQFYD7z0HK1Sp+9gm9KIkVnCn9ueC8fB
ZGpG4/N+ysXLVKav3ABWs6NYp+SUhUanuzBkMhWcNK2VQVUHie4gYUbITPnD+MyYR4Y56Ym575EO
SO8xlzdWwMPV8vqd4hvOPhHv8NXUI6ZjiiC/9sAmg/htPHI0vByQcO3Hq6NDfcIyN+DFeRVtoLmB
DC+yVqgyTw1m0IMtYQ6ooc+NMrG6bB7z9da0xQ6/RkKA4ZmSE3eJXduUOc8uTyncLkGuAJFRjeHQ
jprqpIzzgoJ4s4eD4HJKZFVNwuIjfJ7Z0Ja7lix/4pHA1tiN0DrmWeJTPGHwjNxHdu2LwTklITQY
wM7nZXHrgcY2UFjHzRGJznjxgI5VngL9FlOWbOeD80tM9BkVZQdvREUq72Kbb6Bi339O7kZQkftx
M5EvTDxA5mOIaJDL3W+uQk/wy4CgIv96dsaD+7UvG5pjeMLAbNKNQz+EsmWMy5Sx0nkhi5A4TqyB
GOvcyNN6k3m0KQzv3E5X7ZIP6pKdiBelmpdVp6ji3nK68q45Ysb2kH4GDQpiVYvlCQOJOCU6xdVw
uVyj2PyxxCyZPpmLiEZjBGbMl+arHMJ/tnU78uZyR0gLgzPcXLroaf8cw/ftB9+KxWJSLusJMqoV
wFouOluGV25tVVEPmwniSpMw4bsWaEPdfd6m4mMvZKaGlKzLOhGvrR1Ius0c07RcBpXTnUeHZyUh
B8E9JU9H5i+bqaLPxqbzfuFVB/ikJIrcDoXyXWhM3wZpt7Cx6Oi4Ry6UwG8heNc2ecTi5Pz59o/H
+BSj4YtVwYd+JpHuLR/Qe5NZHgh8qERWLdLPTTQdOYcvdpzzwiwv7ydnqK6iTriWBsQmaNWyZugq
D8X9APcGM32vBr9bSGGn+VeCseSWGmf28tHuGQgUfEaPzvQcubFDvAUmvU/ua2P5yX+kQgiWqT0o
YhaU2+o5DtcNxFMblBe4hf9ZcPYk4XK+CDFeyrfi7o4XRItNzSooCzDlKjp37RvrB9JfMfXu6Slt
IXS8D5ibsuomMwX2jVs/HNJOfkMl0jXDpJZ00abNoPgrlvxeoG1paxSL6SxniaFPBOxjLTE29FJd
Ki1M+M/hmtJyyzAGHfMZjP2mN3rfI/x6KvqYPOj8diYcX4AuJqux9Z/3azTntRGnVHWgbadXz3/F
i1tw84afZF9esWQnEA2HrytWiNHoOP3Fk/viyc1qUHr8rjDjKqphFRqRBH1qvk8b3lxSHEsylOfH
5u44mtmL7RkWD+aorOI6MvfNQshfP1ztlf0aCwiC5NwYxh9NvCh3EgjBK0D2y/CfwjzUYEDcQjqX
wzMBCO4/kr85ru1alm/5b7ExWvfyez+wdpH0F1Z/Vu4Rn5xZv5rCnyjVMp7UjeKAm+8bhJvD8aJB
l50139aVo9byYo390WT8Jge3n6o+IfmI99IgPf9bTaLrIsgYDMqHW8LwjffCNnIstR/gNAGmhcoy
guiE5cnC4DCSgEJ3Cog55M/neChx+8IXEVEjUsiW7UumeIBvaJfneheaGJjR1XbhdK4UHTLs+mtr
qESAN0weKScvD2+akry9XL9d9QEg43W9JZh74SnoKh9Ax/sMrk08vkOjjZsrse+COCs0tdcoGl9k
mnE0En1+cV8GLXJ37AXiSCLZm8O3aM6FDQSAQaFSHkzHQFkDnrlT6W5bSXTUSZdAFMpz/v2LpNfs
jFVMcnHkXe59BJ8dX8nrFM84L+N9Hmp/FKkfKzL2fAGM7K6JnwianPH1ElpNGvv2POoRiY/J3ZLo
pLau7Eo3ttThmZxranrhss64fjc7noAyH90wQrEusxkbkYDRQy3MrAb6DZUzKVvJOIXAE1VrNgAV
QZnAdZZSQRlOW/Q2pR4yxlGf6vuHqF4xweuedSUnquJF7z0zP7k3gq2ADBMoTDhc1P1nJicP7y+L
ntjE2J29eQ7HbYV4WoO+h2xBCeOo2BOCO6jRYtpct3eaq/fKL7Owa06pX1AWjGf6694r2XSog6Qt
7I0VCYfpmfhFDZ8bYCxfPho17sFIUsdzYa/GF2bdERJqxB76qXIcNDstpNkL9pVRtWKc6dBt8my5
WinchtAAYqZV4fVcm54mM9NujcQzmc2TgZpoT8qOgsRgOIQSt3hnhR9j9HXXTmIgCGqWtgQROkFC
BW6hxraXZBR/9tFDtGP3b9a4XFvejkDLHiuhuiyxZ+7Z8Zsk+f142uAs20Yq4YL9mP8xLCd/JVQg
Vs8vfaCqv/BBM/27mr4DP6tu6zpsnb54J4QglXrgygt3CndXbKBduCPx0C6CILyQPWmWu4EhgBuu
5tSpni1Ll6TTJvpeNaXh5/gwoYEyR7VbBRRjEqH+BzrQJqnlQTzE/uvVsTGHm3bWiSP+IbOGjRyI
Y8dnBbEI/YKhR7q77cGDy6SxZzm/6J5IAlak8jn0dfG99o4JGaOABfqOxOE3DtS56lSoUKUemqzY
Pqm0uM2gay0e5hvMhhBNCXWxnMY6+vVinUpCb4wSc8/et4JD2agSaoh8DT0BOPbAkS1+UIE6nIjx
1EOcgGF4MWsEhFcNNulUHJK/jZA+Ul9tdJKMHNW+kXFsc2qkfQsIRPIQDqVTh3tBU9M8ZXWAvjkI
kBVJjP+TJoZniqyMQGNA45NzEzPNXA2wgQ2yQQH8Dudm8gboWGm+bamLonw9lP1pzu73tyY7TXjj
2ae2jk0m4pc2Q4D/1ywSxacqmFweGX5WLQRaRWi2cUApraZAsxsWscuPZ9WPiLIfrMfV7Oi7G8/z
1UhXHencD+DF+aDStlKb5qoyllXNEzWRvzx8zKnQgourG33L94Jwb4f11yCjLlxwOevchlWs4hdP
CwX8apQ6/KwkCyuR89w0VIGiifX87igo7ynR41I6je54autn/ZtexsWuIqnQ1YyKybQImoZL46Ln
3WkIg0OAGAbCTFasdkAVoK4tMa2HlpQ42fAStlTkC4vthzuK7S5DZl0r+0JrflOSaVarbUqTc/NZ
n5tXXXvnnxRT4jcUugNqhcEwQJjwJ+4Vyg+2bzN4azuUUZmxvdM/Hb600ZYtXF0H51GldmiPL63f
weOmIjKyNJXQPBfqu6Vg7GjEpWTat2ub/TOcKusLcmwD5jGLDxw2MHUzC546hAnGSkaIiGiR0Ubn
UToeXtFWBhwaZ1lvSYSZrzn6pTVgiU9LHpy6ARI5wKv4HRocA7z/3STSw7M4eWA9t595RAFc+ugs
H6SK0g2C8BeFkdEJbXJeShNxgKyIpBURdreIYjlinM1RvLnDuuzzZU+8s7Z30lCYCcBYMgN7yYcS
Tuoy9M3lM9eccrXj+JpfAhX09LpA4Y60y87OYg92Sk1fRxc1Mw5nS+krhcmkbYTFyo47U4cF+3Bx
QY0yYpL/65hHLKdP1lbOdsxA2vzge4TvQI6HuDJ2OuJ+yBYn9ZFHdKHv3VlvNlhfd4kANNPjyPz/
bOcp/WCixjxiE6GUMRRXArd2qg9nXSJJyCIBSB1qeOiB6DaOBpDB7am+vpv6lrTBLZ+xAhPQA7iE
jGb4fs1waNl7ticZdmQE/mn93QMQ8vTzZ3YEtJoiwPqAWteW4SQLZ2b15ImA7EqjdXLINAOCHElF
I8zORGl/twubGH8CtgjnTXS7KWxSCioYyEDz8Y7ncAjaJW3voT0Qz8sjhXYODE44Vj6kntJhDzF7
yIoPFjOtA4GQhjQFm1mnniEtxwVxn0loQSfXeXxtqzZWEX5A4BBVAy4z/L+O/0qnDriwlJi+CLXG
UjDOgvoFMyB/PdkJr5lUngwaCcHtxj0IbZ9D5M14RJL5ta2QZ7KuCTW3OVe9qy3Id0efEfbC3QL4
pI/ZvsSLgp0mL8eOaLYfaHjqRGTxXv23aX8I5OiGoOt71QaoxmzMxajSMc0CdzDEieBwqd9O5wdr
Y6MRX10aLWFT77NQ7X/WyiMrH9gmhRGffFZ4CsV6iO4ZHZl5rr8XCujuuY9GW9L+0sjXoK3OXih3
9GPgZWtrGzmjWrnlrN2d/C7VqSqpRCF777ev6fbvP9E08SpP94hWEAgLNCjEdv/yeZtajGVev4A5
F1hxEQq2M9nssScV5Fc37UEHfYVjLVux9mmPs8JTGQqDsyPX5z5CMIZOrVsZToTZVl/sXE3HGuVY
r40o1M91jdhoIlhrU7nYRcnkWH/2KVF9EEbe8ozpJamGqHNy1rH4ONxBbgS7UqkLGHn+UE/q7prR
WLcvmUHK2RtJlNp/T+Wjgu0ZVjH9Zf7goGfI2xekw/ea0ocg+Ee7cPeR6yF052Wm416NlCUPIngK
dMJYnlOzjfFQbnIkU3+BH7hKowng8rNzJPBvc7lbW37Ckf/IxMOLlX3GVIhKTInnrRjODxwGbn78
3yzXMV549zyrDyn/h2Q4KJkSaNtTZdd01FR/LX+nACMkI8+PJboJqoYmz2+Wmm7fSBNzsHeZ9EUB
ES+ADeTb0o8b7otlCx9FR3WK+h/vELDDnZk4gPm8KHG+HTcm4gNaZzOlrSj0OxFTaPDcKbaxGJ/X
nESJw9udUwpVGBgKeXuUyeToni0rMYZJy1xffdb+Lu904zTbg7B5F+lPCcHolYsO9nMlvUxjTPL4
gvSXmMyHRDHMmzYTGevGX2U7nQ6hNJHNpvbMQDlqNgJhDCVvBKMwl6BaDCJUvqlCVksYP9nTS+ed
EY/SxHsEO9qMd86ZHyXg2DbdUbCFXedfsGTvRnuH2+SDiyQgkYpcXzvtWlcfzSpSFL7f+ZqOSFiD
a5own3mubP9BMGDeT4lCPHvZZCdAE9zh6b/7jH9VFBAKGLxkytQ3oPd0IAQrxPC0/LMCH6F1+RNd
LPN17/8WXYzwp0Eb9Lj6unZ6x2jY5a/UElIrPYGWrFVS55xXh6GJ4yaJ7YUyrOh0C7+4ajU3rdSX
vxm2q0K4xHYF8z4846fqZotk6UfvuokFP6ETM1PfefjZRtuO5hLfXts5iy1VzGrLwV5Sqw+Z2xt6
hCjmvszxqBjSbtkTwlYiY357bFiAKXOP9B6M2CskP/ZoJ8I3ltJI4mB23jQ15roLJyCDP4xNu/xV
QQfMXV5DGkezYmFUGK59wwXOplUi5aQqRCAX3k6+bochOG76ihlqAKyU4+Qn6wdzGIiTUHAQG/8o
jKF+X11xmSwUkjSm3mL+SRoopFyqDcvOvpZNL+xC5qQ5XO4jxTJr48XJ6aBswowTuq2emzotUPw5
dhGPlpTz2W8nXMs4eB0JvIWnlSU8h/wbrfQeGb1m6m/ozVHDAEJmpA1w7/nouzdAHYamdaAgAtoF
N4kyqLhF24PT29bF5/UsGh0tgQG8VK0esvc95DGNg4IQ/6VmHvwN0KGOqj93M2DgX7JAlUVEr6R/
KOPmUyXqVLUFgOFeByXHzZFS1MIURkgwPB8YXBXugtvvYb6G52Reg+PGnCINYAxt0RHNWuGrkA1b
ADn+JXVELrMtO+1VUymKMXnqqjmSwyBAx+MfmnOpGn1pEkZe5PqNAAVKtIpY9b7koRRNXuOX+eQ3
r4UNyNw8A+dlm42pXphoF7jYr0/oNLUK2XbvqpXGeVHqkzHEc65YjJQDg7ySjtb2ITKkQ0wn1QVH
/+VcDyUfwi081CT8ZnVyqD9w2vEyXR5VaPtWA7k8OxCywOhtaxLI2pwjvBoGftEUUPckW9eepCnV
IVkquKels9mGuAYXUBrLqihsxjwi7/zB93QgERe5pR32tuE5wegjYPxfg5100hqBUrITrAfj5pJX
ZWa8CDol7oaAzrYf9dEhgYNZ+q5x2p9ekMfmXFc+4+cnlqfyDrp7kodbGr0ur7unDGXQEcbR7kJ8
8bvp13q0/pfxWPaxfdFKF/F/hHXvEMFuImf4/R1gamg8x3kvZTCibzysh3kICBSDCIuzgWuqAxMn
suOsnVevYXstcgJl4a/J5Ov/1x2aNQCOOmbe0ULHkUill5quiis+zpVFKKpnt3pA5rJMYa+kkR+M
TEV8j0JF2Q/jwTSRk588B+yr0z40Pz4oLB9qbaZNMgBtOhLoHYKnuqZAibBSZEGKHCjrLYLVpbl8
6ZwbJkG7y9vYe7t/R9U7IcHLBfgOKzSDSnuS+M0huPC7tBWrTcph85e8j/tvaTGtuByDIBzx/sLY
3BO1tqRMjayeTR5VEusTZPUffCCdhziJyngYnuQ8AzIWfoFMwSmFTtFylMOf44HyX/aEXIteWMCs
1rY7ddsaaVNZgUaF7JttCQuC0RkqCiwFJokSh/FtauWve7r92/b/ur2lGngSjPCT1R2g/2qLlmcA
LH2Dcy2BL6NtpSaiENQILUZkkXnfK5KCHTc5TdL5YVz3hxb6wK2hMG5ZOL1607YuCqWRZ/RbVB+5
/emnWb2HcyfVT/aJuTvQHOeQm/0FUsiewh+BhSuNzbSx0wjHmlNBMKlIr8HJEEORRdzaOeXkP6BP
0ofqhLpB3iJzSTaWRNz5bV2cYLMFsD+svfqOJcvJqUkcoRbtxb9eFfvak0D81eb55jPexUmImBMh
XE4ZP8/UlyzSAdcWUpVu+7FoN5X4VRMlot/yVZe+y8RvmiDe+CC0DCYC61qPFLJASBpZxBtUwiQC
UuEbsJFT/sGvvXKlmeIaWfi+f5cA8l6eNERV7UwQqm1z8sWvyGGY9pR/egopuGJBHFnt95isONUM
fRRDUFP/4kpUF8guzAu91AOHKMEyV1t21h74cGUx4ShQU2TTVQ0ZY39XHsI5mak4mmW5XHMA/4J0
wsujkBBZKclEobi9H9DqrV4lSyCcXYa70o3i9fzK9zHzbvKfMkB4UJ7FCseUGBzCUgDl7QScBsJC
S7mF80ipBbDm2qJ+2F/ylFj/Zg4ZAfqXRVRSv95Lv1YKMBKvGuBrGzfnLTkISufRqU6q4o69MbE4
X2NY4n16lMFOG5W+NW/3uuVBpgq0N7s0cdkiSehB7q/foPw1b9i2WFUwo4wRFgxNDNmFa0w43I9v
DL93JQE3jv5F/rAABjC12E+zsGmEZSxAYI19VTlwxCKrtQ7QY1APyLz2tg3xhWH9muyebCC1oMKJ
BYH9e6MED7/VHG81ajkVgZXTqa5d6WK2zzA1cNaCZgp3xwCabyk9Eo8uoV+vidYB2RJ7zrSrmG9U
8g43yuo0ytYUCbh7KCjbx8l4SmfnOW0S43AJcDb5uy0M6B/Cesrifr8zK59JO6ErJubfla0VpLqT
5WI6XHHq5/SlozjNslskXmJExAARsLhWzHjnHj3RF2PLLf9fa25pi2ojUP3yvv3ziD5a2r/Lqu+x
hOKANqGGG74PfzzCMgIgh42SxDPR5A4I3nJt+nm/dBsON1a8S7vB4IOHRADyMbnYaiLC/ETev1lm
WERIx4dDQhYWcpTzcJjdVZasn/EmDqKvHPfaVk+BhRqDwZDENJUlrWu+EL0UGXHSTwwVg+Ubwo1M
uKqnH5ZsEXKxhXpCHeNC/Xe88mWMSYP/wb2P1cpz49vyJWlGsy5EYGnW9HEPA3Z8eke9Dya1By98
2t4AdHsFhWF+0fOoUZEIQyUsyArKNEQllRX1W/EikjM6Nm2WJGO0Bo7pmpILuOps+OS98kp6wKw2
pqYA6kKI/MFoW2vFz/sc5UW2U/X//YcxwNGoM7zKRijgwDv/J/RQR3tbzQPCxX0zrN7cfXWSQPwp
vWeKS9i5WB72+wAQNaoJFAuwiONZz5rBmmI1io3606OuaaWHkLExSGAVuyhJv9pTG+4K3mqA/Ogc
tQM8cC7M5U0wN4cPKaefEBgjShuGrcbsvawB0ImkqGGo0HB6cqKUYTLvbU0dXcWmkncky7ScWyKV
QAsYkxvgLYnSVBrTPn5O5yhX8PKbjB171pKsbkmYj9rJ7YX37aB9irBYFRJYqzKwYt86yggvLEJt
2XOa1rpgP/G4IY3lKLKCYLsMoNa2OXXR05jvooW531vriSCS23ZwFIMjKy+tFQgQpBCTo+wFX045
cH6gQs8zzJh13GjKQQWEytWPDTbypCa1UvKwgV5IVQWLnynPC94KB3/Yq2UVSuEC+29Z2DVvVyJq
FZEEQDNQOeEFE0TSWfG19C8CnNLSvl4Dwp3EvOA1qVQUB1Qm9qdHSDaLzFiwKRroB/JO88wNArDs
mGHGgFTX61GPvU5oOJU+iLhB2F4mdxZiuArjuUrpFWhJXMM0TO+v4i0pPR7vYn8m2NYATz099Um0
59pRLfMSa/leV6EYqIDOLgsrIR0wlWlvKkzXy3yp+EhxadWW8bcBBG4vzeLOijvCCTOXhMwDuD/M
KmHh2e0dhKM9CVeEVxFQnMkITwu+wAxGLAFwbUHLojWxp8ygI5i7/wMIwR4W6IlOeio48jycKR+4
FkfhzQZ4pV0+JjVztKa8ktwuKj3oxtx5xztiisJqyhCMpxnlLmBVJWmZNfC7ZP/8jjRuK44PB5mL
kb/oYLOReTnPokmuZipl5H2ZwUn9ILLY28qxw5DMIl9xqHPLMRxz2it3IsTws8Xfa/+rxiB78e5O
ec62zuo/Cekh0Y85KR+cKf+Zsmy+Rt7Upw0KVQBtZk7yNhYALINDlvd2zOIOTaZn0n585lJ3071g
qCohVf9u1umTHHwt0vgMSDnAUN3AWnTo/aIz37athhy0jxhcYjo1/Gkw5G24ffkYPGyiKt4JyFDw
PgoYzHeuMX441zYfBefweRMHYJywy/90/9SyKmYALvzicnDQxBXNE3FA1JhriCqtQXjg9h900zIB
FKKmqPVuCbstllahiyl9mmpP7qS+iQZWLribZefSl2CJXUoEQxHUrbBTHnjNiy75aTUsyN4XlayK
d7rf0NOZCNvbUrf0htTvlSeDZW/3YdEShwzL/4lg9fAsb3Raou/IwyVp5PxiR816ZgbL8IHWEnnu
0FhA9IO/eXAputjWUf8hFqgS3zk7PiiRh8jSjz484jvGj2Oi+rl1WHjMsWqDC/204Vupl/+wbkt3
pyEkxZSm6/gOrQel8jjLa0KQjBtjBRBXkss+temYctnmIkC9Q5e7pUe+f/SPtM9gDC7I3yAPEvQm
t8eJ8d1ZFBOsJ5jOadZMiWFrcvXd1ROsEizw20VnA+WqXGHJD0R3WPHV8QVsql1nOjkuBDmgT9fC
mpf1o0a3IbCfgRNEpVCom6hhTQf54dLStudpwJ+gAxcTvRdtdRiB0mt66R8AWC29ksAgbqQEIOev
Vv+3dJ0jXyH/a9p8rHoYSMfKNBara4qduBUkNqLdeszi581yge6bl/W85x7iHJCulk3qiz+D2H2A
4tWksmAwtnB4vDCTHc5Qgya8rsHaHJdfQUiUctVqNhL/n36mz0voXRdlBqrW1iFZaAOH6EZ0FRXn
QRdQ1DL6w0MsYykTYyPJEjiBuY4pVYSFGo055Cb3L0Jdk1iJDBWu7fpuZD1xTJrOM8lBfuzlFiNY
WKpSKlL69aCSIMtSTx04knQvTIOk0LeXF9KRaodmnNyc5QAlU4yDM8Zxppwpy+dA/FDUKzBjYpdU
ERa1V9Pm7Pw/OYJzmJA/xpllkZtDn4tF1zqloSZfT47ZjOD+i12WHMTxHG+chU7k/Cl2xW9uHYDL
xvLEfsMLt9GbPwvWByMCbzNhAbMa01zEjoJEy4zeGJmgxvwWVmSzcKGgc6yt87QrXHUgW2buj374
nz4a5PQX3wM9iiIwU5Mliizf2sJEPNcMGaG9voXzgbjuXh3lmKRMsnv54MahF2/ihJta41aGsR95
vhB3B1J5KyI82u3NQyVv4+6l+/Uu4q137ehZDwXDdfWEZRp1+YZLVy2EGhXi5twYoc7dGQebAwW5
vZW6pE0i/gEBUTC4+oFBlozGb7oh3BHATslwvvSb+AJiBJhGzyc7FsmOSn4mVcUdcFzeUkFbrpFn
hPWGpC+eEY0e/cOxnMtABDYTFkxpEcJoNCRjDWRlstefg+Wikz0w3q9ZQJHm/Lv1crxUKTzp8/c9
DxnzPWy41dhBw/RGIHgXhPHOk3i0gcjdEvJJDGOLKOjh81AjsBvTJog2TAtWaXWNE8Dmt48jDcrN
W1Bz+ag35zxBYGlEqHCrWkjHShoP/Ic84GzLwWXW9tZQnkYLOT+iRdvsGyv5A9L0FNQ2a3+9ZSmV
am+lLT5C20a1q4quC4dwSCh3/aUdHgAKjs/wGLeXLSK+kL5dVc3Ge365rZYaKTCjcd1ryRJoeIUe
bypqDXlljy78+A0G+XNNfdQw8nSRlp0n7TRCmdDx4bBha/npvZ+aFFx9YJchpR1Bkl3wgL+TiLtK
8pEEK2pex6oAL4JS7+dfpm7AuJlfLFFLbPhcrlbdDjG605Bj8CVrz2hKfISPWRTYEc0qbKitNylv
P/KwBiCfO47EoaqneZQ8stZ1UktppZ5yhr2DiOrPynw+7RHgmDpLX26HfOd0Ci4H3q1fcdDimcRT
6BA/bw1+VVU7LPCrLkNj4rSmZgdIqStj7WDGTBUj7BeAoEgcql9ex+GocPbg0tlKwS3SGoNd6fQw
wk0zBD3RWKKX4O8Aeucp73/Hm/UfwxTLfsBC6IohIXnt07AY8vcwDF+yua2LgQVY7BBxcGAxmk6F
j9kEbGaxEe7Uf3oans9vB9rKHxH1/mM/Xi1RPRCLfAtp4FmRAdUPXa1WV+mBbtFyfreLRiOuozpr
pH7/aK1f8F1kfNP4HmG2EvPQszeqg/tPJajMvFACllxOIGqB/4VYuSGuShJqzLhMLlMhp6/0fPCQ
VwLTTUqOsE+RF8qhGb6JFfRg392fi3b3RKpMKCI650gr16VxytWEkJT8POHaqt4EeVuuP/yB8Gmy
aHWNLrEGhvRLzp9FeDZbd1CkmbiDqn+4dyX/7urV6BGL62jkjTTyuA6RsI59/q8/culDj3KiO6L6
1UgLzdL9KAK6JG07AZpNrhWZkvuJecC6CRJpMF/6APvyWQcdo0SR1JLEIchUXxr1LAFgkRE6H4Zq
lmxkqDdGavuL0TRF0csQSmKzZLmLRlHvZkt+XPLxnQOGBkX3qmrrD45gabinSLXsGZh282N7tOSs
qqVsL/Ck3Y0CTez8uDGZFw1r+05DguiqGVLYSBnCg7TaBz74jBuaB0JokfBM0FT0rMbSby5/TuwL
y/JmI6lo600k76i9VUphUlUhYYM+JOf8/dwTPE64DVMTveNLt7VpqNPetSy+COIJqQoSwjXWS5Si
hmV6Zv4Hh8S/7gPmKJx4FSCPyTIAQt8GRBGx3Nu6bCUj7b2pDAbuKoUYsHXVGeTjnaqkFZ/4rKWZ
8su15TYhoRx6MfvHVvajwYNF0u2sttTysvpej63yzhz4Q01lMXFlJFzL3iQVTi6I5lMnM6OqmKOI
f9ljDQENCDwjSBsFJhibxDJYdHEhJVjIzvlTn4a9PNR3OIStMQ4oebyuQ2R6ZOPVk7EKmCOpnnZI
w9yLNAsUQlYoy8maEjF+BC6v6upXYiCdANn5HAY/3RHH6MZ+xfsBkJrhcaVTW4yIkBchvntAb9CJ
2QjRS78nvtqfHbP+tk3ZRGx3rf3FAaBW2HVBIk4yHuK8K+QTfOl16EKzNnUM6wJ3cPuMlK2LS3VR
aX5zJ9K/YTqzTQ5KL3AOyucsNuN1cA7EoVMs5Sl9/c/m8WQw4D9849ANbd0BU7NQDeUK9KgRyzIf
zsXFpw13lIUCpTT5kG3qv1dFy0ypP0l59dL9z8LaFec+dUeLpdVcOSw8nUhj1G+hi+sdANhCsohY
okvBNbl8abWG8Eo4M5gGSgSgqh6SIgrQ/YKTjTvp9oTvVEg6N2M+6bUqnmI5rHZ3Gt85p5yNXuzG
mxMZ8A3Y9m3dQQM013odLm35QSOo6E0YQjSYjej70pidl4yYZWKvvEwlBg1XTS1hGxXPQdV3IHf7
bVr/jcbke55FURfy1minfVCfPavEnpyDgrNCm74FBlWrQWG8tI5q/BuT53naKyyuvMMZYwpa/RrT
0qmvEMXbge3a4zlpZUSEV+0QRpGpFiqTyzUGoluBLR2g3FfBdKt4d7zaXtrMHG23PIbPICuQwN87
LrVg+RrXKoJX+sLiOzibbfrVrO2Ua7apCZJ6pBmWnnPjF+2GBERgsNVzezb27ANqknr10KBcVwY+
7ni9bI5z435lLg3wSGO/9oz7IDLlh5AkbFQVzimP71fLWd1NCWLyd0aT3NqRG2SgJNUnDy6HIG+t
zTUYAbluzY7bGv73823qAeM2KGHcadj0Vqi9w9KjVjKcamuuhwYMkuOgARzaCcLKx6A4ei/xMvjc
d33F834AHls/og3AvzUMD17RIepY/PyjFu3iDqSgtYstjVdgDQeIy4OebH54z0gQOAvfjRnff/vO
Q7olHxjkGrbREySwi4Npc9sim3OtNQcpFGg4jo/5l+41yo5Z1IysTC4wet+oyNU+j0RhVbWa76Ln
CQ0Z0HvLX/M/iIAMJOgF+JYq1NBXUo/LWHcF7h4WW4JsADatb4PGJCg3AUuD14uT+ytEp6yxAd17
uerdTVX4P0Udlkk+OWKUcEX68mLkJ4j04EO44IG0U5c70ZWWdUMjF6u9huWF9ldbRahOsSX/F+qq
J7dK5qC03SxixnjvD8TW1jdjJADEww7c9sivk3BeTwqZADXSEPSB6ItUhTtx1V/pSi+vxYBxiVeJ
/cR6+O+ZIk3JZTyDdhsonFOrIFbdFRCI2qGkRX9pupcjn7YEWVqKrFVJad3PDA/vAORxu2e4YBA+
lJHF7v+tB0EPEkBO6F3ZEgGw9MU48e19yOQUj758TTia67Jg9tXi3C9XTsJzJYAdk7KhCSMRsa0y
+4JmaPRUkTnRUwJrvfXbhcM0gCZiFlYg7+IMq0UPscXiUYVdG6A3EBt72liiDV1Al6tQdBo6tIl0
zs3UuV8ptBab3LYE1lu7BJxiUvP+SyoRBGvPHmefUlJFu8oEUV/zmKSLsRlhYrxNKeUTAKpUXCER
og6E25pGuJONG7XfgqvMJebQfOCMOi+O/Sf2eNMT/8AgNdS11Il5apAkaZJT5oQf3GXQ4/1fQZ5f
FIotfBG40NQGV9vMJEILAmB1MG/BFjFC+9E6p+wGGmuCcU8Eqs3LE/kBDGQhKpEB32/U2KMbhaeO
nJunwnuqiJtbO+P/2m4FKTTUJUKD6Apbo860qS263jpN++E41HMUCjbahygAjaDz70rzT5+VeuuL
6TpuZTZ+lj/Bk4NJJlsjvh83+0qBmrroeR7Ja5CjnEbRQY2i4rZlV1CTLivVj2dBhRWv8Wlzz7W1
wq+g5NNWrAtJ781jl4i/AqxRD8Uh7kB67YB3xkTDFyMB6GTNhwbSZVt0ryVqgJ8EaWeuU9nBGtGb
hyJJqTO6Oh6RFeBZztR1gsfO788JZ4GLZoEhs+pt3KVKlqWK/2bPN/zZ5WnFJLmShQkkUIz4pc+8
R3TYfpXKTezMN7k6ZdI6wSAoq+HJXnvp1pp/qd93CvfK793wANiUh3eJ7wpijQIPznujixq0LJVp
pL+kxOJRNPBmXBMvqKtYVVQ1ulAFHWY79IWtUF/RkF7w7jiNdhDUHhkeJBtQlDZnB1doA8xdjgb/
1eRq6AmnLrVKBpGqVLQFUJO2M2iycQnAf0apqT+9VJMXJN9bGRYwBTmp0m1PCUS3f92wU4rcE58H
LS8uEB1LZK2M93ZtdvxEl6Yu7LbBf8+Ixv31SOgdYPjtcugF6Jx8MevJIY0n9jr1eNYE9Ow/4FjJ
x0jWV0RfzYNCuwtIYTR01FxMlYDx8vmp0CR2QgVLL10D9aoa0w5lXl3XpRCtzH6dP53TDncby6Qz
41n4+ZjicTTehQN9ko8nkHPyfNXPoXFpwMHZ9+ojSvz3OlTMOiI5/7JsKvQ9AUt2GLB+9cUJjpli
uTBum9BUU5i9ocV+LXSqG4lVSbUMf8i2tFcfKxNEmONgBmrY8phRBiWuN3O/YVuyOWKVyx+lkirl
oi1mio9c6aeqqWUfocObyj95xj9/KtJpNrdD0cWS4FFWzQmjIwDu0VmhBwUwJ1kxtieI2rkscEq6
XH/12Sy/NIkC/HI1m1wsRPdQ0cDIoyQEXIxAlc6LmgTHM6nbJ/v+Me5mODkZPqft/xuWzEMsnfj9
0hvCPsjS/qT3CrxRWV+kPJA7l3An9A5ABb/Ve4AKDYFtnNZEvxQbdQw+iMQSFarBu3BJjLG6PWRf
zGjMnjUzq1BGM1HdCdpI12AMXxmRXU8GBWJmIG9jJw1fPTca+EN8e9TBEPfyzvRlpJKDHjcYXQJC
UhkHLHV/UOLuh9oKnrMOk0XusCznj9rYKpq8ivCF8oDGzzWPGxU4DeFf+piPmcMkfGWZEouXzGis
nU4amLszC2v4tBBpag4Nr+7sQ3wasGFVeGSxAwALt06+HA9Qou+8Ylso57hNhH3/Z6Z2pP/MmUJU
a7UQALcy7Dxl9IC4sU6WlKh6DlizRDSa4ZSv6tO2cUw+Xx81stqiHDB4NOeqy2QFgqB6ySkxcctg
MlNpOCWwk9SansaDCM+gRahXoSr/80G8HXWWkg1jRthI5eiZ3wSGjOjzR37ntW+tp4EGhUocAgEz
m8bsKlTh1C7wZPwgyuAnJrdW9dc/oSD+18Tr/ZB2jwzlWQdhvh3f3qvFCf4WIllkAQeZxZvXq6Ke
4jVO/qvQnJRupcvNnSFK06TOz6i6AGUA/dzYslFVEghy/CIdYOq9TolBHoa2BwC0H1VCjoC5Zn0y
9SKbR/3ffAQ9XuBVDYT0stWJwu3tKgfcknr2z8PBFEKO/7gwhKyf72IgtUtbKMPrhBiBTeFPAsUL
doY9jjrLAjpl4b0OrzIblW48zZA/VIEae74lfXpxU9ldO0xEXDU+VT/Fhn8JREdz6+S/+RgMIA+l
CbMFdSXYKyk1RzylGOpk0vb0SO1G6BlDAqgylX8QL0vEi2/oRQcTJHzhskZ/2TVjFpx+P6RdRAuM
XWJzygI1qacda+AUgiiRcQMuijNzxmyGS3qZ/y/fLApaLhzE2FpxEV9a70e4JiUXgyB7NFaORYTf
H1y65NKfHUFhv0YpCRoCXSa9btsn3lbTg1uZLJmV/tn4Q6d4+KMoEE2N8WzqhK+aK85h7cit+EUH
kDEKvPgHhNz8V7fRYiTx2VUYMug9gyWYEeIaUJ3RSbTH1JJ9RPp942IsESa12QZhEJMzymDuowp8
RdOBHt++8j6C6tqfaAcIpSq7NWW1P0En0FRJaacdO777dOheo///8DjCjB1Vm1xzJ3Yf/DXIlymj
sZqIkEHP77MkEOCz6JS46OJbCYfFBi+ze0AFnJCh9Cv4yW/z7y7H6uQDGjnQrtEnOE1l9Yh5zd7z
z58RflfYUP0r+3Yf4gevPgyS820nrypsP++pLY3HruDh9rL84goxctsy7kMved7wBfyMXJGaV8xW
ZpA8fjzAfaCvqV7B+s13t1TsvazqUAxpxbTaT4W5t7xBww272ChDynXF+uYw51UQ2bGa/eQGB6Tq
jnfnZtwCka3fr2eXksRWlWaNgZZ2+e3j51TuwAGyfwnTg6FuQjbDEo1PNpR6ZfmwI4cuJsw0Nc9S
rlMw3Kz+G/vvUgWvkp+e3G7MWYSYIpN7x7gbNzh5rszxIziL7BYV29OzZKdcMqrR1mJz3FHVgkws
aU1+iqfMNYxXjN/lba0olhqapS1xCA36Yz7A4lZEuY0PKm/DS9OC46U+cmavYMGzmX4LLwrZ7Qe4
rg2RIU02vQpS3T1VY1HgLA26zYSfs93oGDfLwTY9KTDH7wFbrhYeJZOqhWIBEHn7FakkZUaJ6haf
uWdMYGMwfMeMjYyzbC9ZfiNv3P0iEg8e2ltle1g0X3FZiZ47Est9LD1h3+atFn4wOHe3O4Dcb+a0
7tufk2ZrAqgHVfqaY/1UMWRFpbbPU3tNWKbZ0jHwxZWjCOOtHU67BMpa5D7GlsibZup7D+apWqVc
IEGsZD+nKxt8ZjjDIBHRlKXOadE9amgcgaWMjmWDC+0Jfes3xna3KrDkERmsnaLiEIqbqlTzi09k
n2OstHAOkCGAT14WHcgWRT8v1vikCHHFMGcihrzWbjYmROMiK8KfP37pfGK4dKkn0vCaBK7SeylD
pH4j4QSemfZCsjETsyB/044hv4YTcSHPZ1WSEk6hjcK5eLJVLY3ooP4+GxKfSxzA36uDlVvixoxO
LlTrQVfkO2G/xpEfyn0IZ0vyimVkteL7NiScpTddEhXjiz+lSUsAVkG0ZtvuHDhpZ46MaLPtlHbp
Ko9YnQ+d/+Jz90v7dRn+I7z+HoZ0du50kvBUeGNDVtct+wAkqtXs5Hu/EblEN15SnvgS8jHiTY+9
X1TF7d5OCa0Xjwby0pZU0b4f6jbkzME8NP2/Qou2E5sPh54otuRiCiAQKGYA8/BmsiQgkU/jUW39
dwDngSv4nL8Iw2DLgMUwNn5pYhhVdTS5ztTVYjrdLm6I1/JpTUqv8+f7KktO5C75GD2VBqJTNrrR
loi9YI/PzBa7T1Ri34rEQktNqpZEKh9Svmxsc0xMViV1/SIfCulKH7EL/7vCV/F5PaAm0+iD3Sob
qdMPIloDBMdWApoSZVAYjPIDzurh+Bi54AUewrFcB/W2DOVheODRQc6hD9qQG1D/0jMvEYY1sY2n
XzLqqcccH43GTds/XG0FyQbPzQGcuUwYX+EDqNjHS+4i62qCd1bW9QJVHxzJyV+oR3wpaVs2kFIj
QLs6XCfNJyzodF8BIB331i5JXzTW3Xc22qAmYV8ZIQjKU6pNwYeBLgynurcuFbA7quWK2xklPFJn
OtyX9rzK9qwZQNCdyy1FaA4T1W+CK6VsNdFJ3KKIjjNY/iGJxz2ZRJSwnxq/cebEE/8sMIdxYxaD
RUQg/Eq5cR2xO20VcB+QuH5puh3FBkee9MMTi7uBSiwK+UiCHm6xgFFm+YAAjISKI5VKdUc3CiZt
HaxWt5YAc5vZAUg3Tx8XHbQWKg8eUdIu3OxL9H30mZlifUna7mM1s1fBkHJZvzfu/W4+mzVOgXjC
k4dFd8Qgm0zGqamb0PauMoP5ANslThpFcrZLmDHzxM0q8WpNv6eGoThgpTD2B8RHPxZ51f2ukQ/6
YF1AP18Mzrf5GFA4rjWVhCoGAqDqM3FuCpj4cEMGP3wkjotj0qK84wirLbzYyyi/rkIis5NZjcZY
x8N97SylK9zEAqi0DQqNP9OcknWyGwGvB82oi4mxgyoxy7ibByUoaic1rp6fefWm5MY4+C7ghDOp
NlA9sWy+KOWSDrd+/GG5Y2MLJacqFw0klSkzAwiHAblVOXFpqDo+AgvRgq7jhzYD5CAQ9tGNy2V6
pyPVLh6UlMpMdCUT+ZsRDQyytT2Kzb6EbDekIXolM9vN7qgBt8mV+mu3xuaT0oH9m7/R5Nblp0Mj
FEKzSfd9Gp/E+LkEAltUThCd0R6hDljNgcpauuZrkb2jUDdYqikoRSFrCct2MT/tTbEEWrvdAbG2
hSsOle7Rvt7gAuZXqzGMQvn2rIMQ2v0KPKMibBHGEOfv3i8kMVTzJY7sDg687B+zYjRAWIdxo/or
vCdGnBFGmGxzJM2cyWpn8siTbNCgZw8u9btLvI2fqepN5I7O8fI7riEsj3VQ0HrE+p+/3IoLaJDv
1dEYZ/fVaK8YCSU4hb+6+Vu+cg4JlV9Fr0VgHIcJdg7IFM7JuJTHAlGw/xr3HcLtV/2g7idh5Cie
3lO6w2ux+h0tc2yw7vlXqtQlRLgoLIttwJErODsi0E0v9yPE1nhWjJlvYJROioqyL0JdVdiQCT3u
iwT4PxvSqnRhbuQPqai6AoPVGnI/R+W+1vjWb6AHRoe4am3pHRfbzcSO0zVWn0uBfBOe7ONWJ+0o
UzZ5SopC6TuPCZj+AGAcVbmIOtMWHjD122QwGwH+T0vvvPaSPo0Dp5j0SrrUCENBwqmixE+8Q8BN
2hgXYZ0PHLP56R/GkWe3dR2hO+ILNiEirWDP6cZYy8DAxnhmvMo/jtDCjVdH4zyzfkjR91aACdFt
Vy+PVU29O55xnymiuKIbmovlg2lxa83N7z/HYI8jjoMj8X2WbXN6YdLXgyQ8dTu4jH+lKuP6IYyq
u2yaivwv6Y6lPgn703aX4RgfcjfLuWuxnBhgZD7gG90cdpj2+SQYcrb5aO9HsIg8chGrVTb/eFTB
mx+6PbT8yTNIeJzNCBjsjql1DcBlRfy5Py9TWobIZLWdrmkjArI25TehsEwIr/uU3L6ws6qhOTl4
Mfz535wpHwxmciwS7VpqU6n06nfOyjyagWLmWEoH4tIg6Ufcmum47K/ptGOBgO98E8bB4+0EgwW7
IOB4gomSl96WdCybq8f+B61UUiix/XxeOQ9B51+XKE9cv3viGi1cZptPfhBVuhhuDrIjJOXN4hVB
l0RNjLAheDMG49fH764wOP9ivwK2Sv4r79uTfKaUVkPOeYbQZlRKXGcFTLHvy7QKZ+F5UzwjcpZr
6NW/gc103Zh1P5EYMvye+q5iP1kAmMaOx5b4rvM5HVFLGj7YSCAWzJ1H8CcgRlNnREFsMbpRRYXo
IfLimjRfGH6orq/fMcXcRAKt8488xgvcZt9wTc8T72Pzen9Ef8IB/BcJgJrzi8oMHHY1Zhgxllk8
TfuekyXKHEbM4K1CpLT0ZBkj9qgzDsRQK2kSkafaj1WDCaJkv0pokmqQxDh+jWD5+alHYFlAa+MS
sGC9kuCMshbhHJxT2E+/o2BzBlUuXK3FoABh7Y1qJ+bN4z3wS0FWNwjT3eY846Ze9R9sLs9V3TLm
RcsbKDXn3/uQUsW0MnvGir0rs+KWxUcXO9qc1jvoBYXg//aB/JLgjvjzoOUDQEbhcBdn3XHvHZ+0
6YrL2nbYMd/B4L8aHsh9h0S5YiPAI6i9st15G/AheZf8ozlHHZMeUZUhfRzFEUzzh9e3BjjRgolL
E6PKfAqWILlP+KbAqzVHwHqlmL4bBL2oKj4ceL9VXR62lvZYA/FkU6BmFQ0sMrnhjLVmwHB+dGQL
xOIH3Gr5oGumLyDV8ac2cThlABEUa6fv+O+CMGDG2AF1FogSLpw2iPXEFMXbaxOneG/bGq/lUuJK
dkedeSSOrFBkWK2xaDguTGwBWxSiBklIc8FrTDjKbtoHdM4mgi8WHTEv4Z44+j1UJjt2q8gWOJl+
20pkehsmlcR86Ge9XOKIXa2Z1iWdU9WHDE03zwheBvSOY+jVAjzHKZbpeOfr51Ctx7voC46wBCV3
KXU6NtnKII+OX9JBzTn/eZxnSxIVUh+tpCSQ3UfX/74adKW+qp0fWI2SLzCVUKDf7ZJkbsCpkUJR
Y+gNxtsYPt4bD4MhX3tefry4dq/NDziZXSnhXwaWaZ57SjpvQOHc0iabujSiV9TnFUgEw31BSW9D
iJnIcZkuiQh1DZzJgBBbWnt9+d1q5i4/VvRh1iQH874nWwxN/RSrwUAs6QFWTOAQox4Unm2OPJMa
iTy2rCgMCPPnCjFZVCzlt4Seo4xLwDBGcX+yvyBfzLP67OkUvdHxeFtfnHCGQULrNK60t63fUmY1
FhZ+NIqTFn1nNo/x70btF8Z1sIDGOzsQVOYfBpw8s6JCY80bADyKboLT2Ln/mUljcKwIiaCVlwr7
PqkzIiHPkbWFXKu2L+Zk9fUd+im3Ywa8L2S6HiK6iKsngqcVaXBLAFJeDqCBZ1JtQfuD+XBALnHj
PgeuWrnUrTkIHuD4siyVbU8AAC6aHqUyMHuZ/GnJZWsgVt+TWlZmvGoGIB6dhQPZs/D3O6YZhQXE
AxSgSeXW6vIu2M8Yi4aUkHjhZppo2FYgCO9MyiLaErEtseefJi5oFB8fdm905ymrzIsxoOwZX+mn
Jn52lSI/tTnSyftUlX3/gIx+w+Dxb39z9S8E7gpib2Q3PQR5lu7O/V4lS+Gcd1OyxbRtjIpW3Rhc
nkYt0ZgDAGI6OPQ34RRLxjuxfmB1MV8X53pfTvRkMvhfY32bZS8CGXcWmNC3VQliybYbP5japz6w
YpEcBkaRId0Z1d8PNbVxgq9sjZMstrRy2iga7x2jshFr7Oju437jXuh8a052xHqn68fiMxvSyEX2
AAopwB80jFkg9iKJDKtvvv/EToo2D/N7L9SZcHcI1WY9+KjSa9R82RKnk6qcULqEOPPOrcMBJQnt
uiiZtzzeNIPL3Wm2bcRCP+RGOe/IBkW5EbIo7BxFskIHCSn9SZKO1vuH6OOOMk7rHQimarh/Vee4
+6xtd3Mu7VJeRjky9kCcUkHmcUHZIn2ZUukQzwqYBholWu1/sF1md9rKhz0w1Yqu0qVlO2i0pKu0
eTsBLxX/5nZbQ55EggUMukDkMCco8j7dGdqywovtVV4nXdNSxoF2x7TBjW3oIC8SLDtRxeMtWlBz
Sb5tjPPHyn10fq85Lg/uqYhx1tFB51wXj9YbBK2Ff2g6J2NvQze7pG55hsg/LBx0yy844kYzrWZY
MbVNyUv5+7kZ0M06/0P3sIYO5rPrNOPWQFhuJ44JaWeAPej6sif7nh640IrnW8OFjG3ZpqYrpatx
hvwDTbzayikA47j1uAgNi/wRkSyLFbC60vL30RP2J3oQpQPAfulI4YFzLaYfb0guavqPqi27Yoi4
9itKkh8uGOC/xjAqiHu8F36OnmhTCi++cDUJaU9KYX5P0rvuXqHiUPkX5Cr3X2G4WuuHzZR6ByKk
rXpye3IIPJhSINgGQey2HOj+LiTurR/Q8QA42MP1gUMTRQaE/qVHF3MnvVmdD5IkxkZveYC8wPaE
GviZMfWUpWU9eAfPuO2IDXbl+jBu1YYX6iOTbZtuZLDwBLkUCU/To+CFL2JXa9LmzondUCjSjysC
bLWlznVSzDWeb6ovAnOAegQ5IjhpPdju7ck5qPBGMHF0kDf2eRe2uALR1MPEnZ0XH1suASLNG4B3
FcXiOuQwm+f3IzK94T0ogDYRg9BNWjYgFIxxJDL1ShPVB3LpY82aOu5PIdYR4SGIp/hMBZmB7CgF
UGJbPGNa325pXbtCT9+s4VKj4R6R+JuKE8vb8IYCyKgrvK1N9HQyu66qFw0aCFRgLS6aw/NIL4g+
hYh2vzdPN6En1njxpcnQyJlyhCUDYWjzvdsi4p+gmM8Iah8EtIwDqDN1Dvs/RDAybm6PenPsss/G
zL9tqUo/Tho7vZlEBRWArMU3hMghImLM8DwTGNm4ibRpbfrwhiwvZYObIwchniYzPsFZ9wNNsmNe
NZvABQkYLunsYXgePemJC3FGUkPzW0L1zYWRP+Gc26EeNMMKF9fagsvAwOgBgieQ+BziNj3PhK1V
AZ5ogbY42k1FR0kcJB1w65iPgjZefSCs205ZWXwi9T5jw74H+VHDcrLn5JMgs7cNFi86bLWTf2O8
Aqlr4ju9vtuUGovCNG69lgFPn9T7M9MvsMACw6z4Z5ry77SvN6LuPea5t+p/GQeTMVQAmmYdPVH5
YQoDFTqL+2YTEwvQp9pTVRDUPTJxikTsc9IQTLGdjf+WyH+ItLKFNYS2wUJsIIDzb2DPUhp4tH9v
7EEPRIO7dkcVKAbs9kVNt6rz7TUc+8cJ6wSFPai/YL3y7kvIBL4jDCYOJqmelb98XY78Kf2Ej3l0
70PaSRPxoznPVaEQM/QpLshj/uPYTtTTCdwaiyf5P0+YOQDEJMmWQtrsiIjjsD6XMycSNQwsMl9P
xex5QQpzsKvfDZvQZlXaNTw+pjym+BB8DbDfb+8HjpaRmSvOPGlxt1t+H1g98UvmoCjk6GHQTumv
rRtB064rDXuh7jlndKuXPam+bSeJB3dsjWepdeyjpUJBJVhWX2iM7TPmXJ/YTMzPgDylhY4+QBbx
NKTUx6T+Y6v+h2Y1AxXRnZdozl3/BPiQRRSFAHsD58RBteYpJW3r2vEZgmGt9PhxYJiX/ksDspM0
W24X+uDxqoBD+YaDzCCsLy4Ie338FEwmhKF+14rH5Dnapvwwb6OeXO47FS2CuGwJe695Yu2ribtY
YZH9NVzQ10rdB3gRALR6vFnWkTLSFYtu7LJkiRbxvZarPEFntOipNcyVpO4OKQLqAfU+7Y/3wLAH
LnolEXW3ahsIIYnpHqQiPqiXfWCtrSSd/aLEop2vi7e5FLkNSPZqi+b2haAtcxFY3uG/m4CzrdAh
yq81PPeG5dmF7HUnMku8dXFRsgoAmAhvRpppUETJ9fpMcMxVp72h+QMFBMu7/y+8ws/kRZ4RDxqk
gx8a+bo21w4hhtpER9lyhLRm3nPKVdTjxYzCHp1eiQS5TuhEY6qsY1qwItUOZSBmLeBXT1Un95CD
CuyP3wag1gMwmd1waDwDteQ5cctX62CULhE+96UmdfUxmfZop+/mJfNWvsoaoSjHCCfzZR8vFG6y
ZwBHQswFVafcDRgRVeFX6A4l7Xs096+LziWooLE6ep+6SW0N6E1kuz/AYRXCvPy4a0H0pyuv4oyo
Vdh6Ye+z6wt9vcb1I1jK7/3h95Mdx8kJ9TX9RRjPbeukMD/xN8y5FHzpEUxtcpwqvfKYisOV3PxA
aYW7MGOYDKt/0sR/AGJJTTGTLIV0cHtpQA3QS6zS8bt3L61cfYKoB1zB7c63y7oBSiZdIdFWErxN
Hvz5dbqTzCU/HmXzKluCSmY0oxaPgJ1o4MMR34jrslWHKujmUq3P27/58y1JoMUnAt9+EczS2iAB
z9xpHddECL7UJLvXnzn2I+Whl4wXSGg3GbR7ndFfXD9jFZx+u1VsmeHc6JE8KkfedBbLbBpdXhEK
BpW9AijIe++2UmVs3S612kew2y0UB/tHJtz/9wcbloO/OS+7izBzNH179KhSnGMS8RuFW5mqHDvv
t8yMcHFlm96V8zCTOIX/xQx3x9T9xqENhm1rVYt6eV8qfJAAzCruY2wH96y9XWwAQPllNRFw071X
tssz01cdoM/fN+AcbsWdeSpdRzj9g23mlEf74j8VHaZfj/3dFagBuPGI3u0+nHypFv5ohLvG/IjU
Jb+Brw6nGc3XZrKKjNITA9HqV/I7aUFIpLY7+xla3Ty5gkeipHLr+dXn27ZsU5vwyGPN3vpTK3oj
Y6ydU0lCIJa2TYQ4Nz/Oxrw3M0wbufA4hF/4XRRoN8jSjoPr7hxYt9T+4rMGc0v52LD59fyFQ8j0
NMWHJfJ0Eo015L58z5ipXmuTc9fBDNhCKznSIUT8e/3gwXh7l69WE96zEG3bM6en8K5MhiR8UFsw
7BMc5Xh0b/L1JkWsDg2h+CGNh023EpvNFcby8XYiqKf4VWinCKNX13bxQd2+pXmAGyuxA/9jk62v
i+Js1CBY7bl/myMH6mhSYxa9IHqhDM34eI4N0bP8xZWgxjhhvNI/Mglh2/mrFZmTGDdDBynzwy7t
nGseQaoH14dBHX3tv3WPtwNkO8XZflbmGCyFRgOygtatmo+Z+nn9mrKarcQFran+NlY5EOfgwruG
T/r282JOzmUB7WQDtwF0Vaw5V8zp2Q0rDxRIyrhw6PVpgLdN6fJbqASP9Jz72XLe1Ur+9Fl0P6vl
eXoF3EAb3YVXSPOWcTAXNpS68QB3h4NuYGZU1kcfwsv9MK9T5dyjKvUSJchW94uIy5c3dvH9hHlT
UXxKZsKgohyVaDj8YmJ90SiSBacrduFR/tH6DnrvlrfoV04fnoCCtoXtO2fxKN+c0vhT4pGkajeB
q4LxzfH5mdw2v3vEJ7MXeB3mUInI2ecogNdbkQ7t9icVoag87cyAwLxPRUzGhnizPQZva1SY/XgU
im+BYAvFr+hysc6rJ+Z7sr/50ZwAxziTay7WQGyNc+BgDKsLD/t4EUVYSNaOV2wEEGRGa2NYbeYL
CzZNFGKNuYPw6a3dQmeDV4RD/ocNN62X601vy7ITVbPX7OBSySOOSj2bHw5fxi9vRUqvYokk1HNR
Mit8qdeVuLhjm8qgMFDTB8mBgqEI2dnCkCLEpYYyRz/SCHmc7KJTpkU+UoFoes7rneSBdP83aT8Z
fJny+9pDnCJ3xDiOyVICVYoUBuTyZVdO3C6FzHgwavARPYzpX+eonx4QtmLDMbdzzTCMVnJRrSsi
wvyd7LuZPkNJO/nAbD6JVnZ2bJKSGiuzrXaxu+yXNy0BQr/TrqrFp/Hll7qD2j50pZqP4GWqmfQ0
carAppPWMnGHX8F3j8LL0etF+zhN/H7yRH2q4tyyI0Dkod+WiFlVTsKU0qa4HI401iAlbhJo1oYH
D/zKH9XUXr54G0RIsYzvbYZuyCMl+uTiLksH7xlnjkZzwZyeFqTHbgcpedSCsUAUmmBUu6zTygOp
xOGg6EpJSjvIYrUOrLvOv3J0hvi9HEwzUkAUYxLmA9TKdwkvNQYg9ZCRgUyWPzeHs4cUC0l2FpGu
BbKkCK7EGO86H7sFeK7m3hPfg0f8SspoiH9vruib0/3xI1bt90oHEdUngUT8/0WNPC8ifDfbZERZ
ZrcbncjDseUfRkEdnGp64UIMcdzs7MiwsE0blvUlP5pAFc1gTnsOFkVFrO8YwtB+X35sxlRsMuuw
hFUieNZgLodGT/NznMhzC9T46sASI2N9hMboXKgq0K0hKVSUmG36Exjji/PrY+bihnnWiFdu1qJo
1dLtyXLnclD7tj+lB0wDaUw0fwuxOZ9Y+/0PAmzguo9owWidLCtPQ4PTv9Drfx08eWlty6K0kiyH
HaY+O8KozKpv0Fv0uKzh3hwzqK2NFV44/gk9HtcxLrsuqTWRxaSpfW9zu0TGyWXh5aKIEuXe5HIP
n+Ej/3BHgV/s7WjhGS6WzRFq6wUyq/a8anfedBKEw3K7TGHszedeiw7ZefjRgJJQMInZKGVrmz5g
/q7ItCZCd42hPm4XlOjgkhBJPF8b2iRqgoLdMejCkITYl3z8cFaVoVw/l3XUstHbTIyWTJA/3lAL
t/6Ek4Q/YSgYoX9nfgV1WagaqVs2G0uFy1K5/6p3R6B+XxjxvwXc9TmVocevCh+VHugAkbka5MPe
58l76CFRaksxcRZZFzG3ACyk+Z6+bb+H93yPa6P6D8W9uGWNoWCDZlkJjoaxS0imsGyL2k8AQGKz
1lRClM/wrsuQBl0G6MOPXa03su+ofe8VMnwg8Cq6Y+kK8ESV6XjFww798ofpUnu8Dmql9lZ7i7Qy
SZBzqyLsZr/NSzNMGMaFPsmRzJRMFbRFmG/zA6YFu/31H48zft4uO5+cgc1iCq6WZ955jnecvybA
RpFDojr7AU4oq798N6IrhuF/ANGa2vDQ+i2TiY1zzfG48hdtX5K65sBzrDt1NwEbsg7GZlCtrj38
NAkuQ71rwmebhpqtBbOwUFm3L73Itym1bqdEKTj3ZrY2QkxvhYOPFiCMAqpFs9iW2taUyI07tUoa
U4Rdxc2Obz86h9MXYhwK5mTcp63toU2FMbUlu2ZfPmo6WoL3ivqhsmJya0c/h12y6jZXU9xJ7UQA
QN+OFE1iiBQ4Lih/rb8ZBm6vI8gmx4HfqekUjYBHlJ2+/PHQHA0wAHAePQ9ruNymZD8dvTASSLZc
WJHWxvp0qgj8rZSUc77uph+sELX1upiP4mJ91m5//ZaqFBk/Ho09hP04OsgWmAhbyXZFnlKQrgLV
LqKU0dBOHk64uJw0LNxpV0KYf0prG7QbT4BpXu+z3p1Y9odB7FP26la/HlGZXmXPrNBoU1cNUMoX
HjYiWsnsrNJreaIryAQbV1J50zkG2QIYQU2bLCI7YU7RdNidMpsCScjh+BLZo6267FsriFnAXYI5
jgiQNjruHp2ta9ofK1EYLU9Gf0PDO7Bw2cybVAJxN/AmSVi8spSXstnkn/Za0ruhNG008ki4OkLT
MUGa1UVFxsbADMzUekZPwFYqnSNFXPORyIi5c4rC8c89ktpR2dPlwQH3kVfCeNu/ncYX2bxMjS3h
0AxBI/6++M7QzpT5DXZyn+xplMy/mZhkkpsJVH9LhkIpBQRSQEHcTdOukQwKPDTMerRfGfWRG+y9
Ptj02TwtdK1Mn2Fy4D5oe0rl2gAiIP8EZD8FCiQ4mWz1d41F+gLrRD2tMhPl7FGV60WCIfWuYnBW
NRLoVxRQ7CiEP6ou4kqEqXK+/8njTn59UwQuUHdojfYGgX6803yNd/+67Th4g/B+Wmy+9EUviYRP
78pvxmEgRdnFhNPeY5C8CM+2D91MoZS+WmlJ4+evgCLARK8bsiIWNu9/3ISiwQWHx6+9F1KLEpop
rxCHFOQrMsAvjx7QsVTEMIOWsIYJuichNdLSx5k7MI57eKteSTBcoJBBNq6nbpY/eNgwJ+kKPYGF
OIIqlt2r0b6yQ8Cv1Y9V5gzBbVkc4fkfLLyObbaHJMJg0E45Qn3u7b6lSWNhQJ3ohvMU8NE7y9Rn
nNd3UwB+A2RhXZG5vBlKrw0TxYijCPz3ttEKuCwIi4KsKOsD3dptlWxV54xIvob3qH1DPEVIbOJa
+EUju3I6RLZQ0mZTO3k1cL472o0fAT/9I3bXFJ0rPJZua526au870nMI1n2YCdD4dzV+hFm2iD4s
dsjUwbhp7h8R+me5E0G46tDVez3CRXbcN3v1c/jBjLmcxqjS8l+j1H8syaHS/M3zvayL2u6ImHWa
w4mEJUqWYDu45gYeN31IOFBobYiu3bIhnLsEZIFmvmGYHLMjZti1LouJichfTRioDFk/R8QuJR5+
6lJLbZU3hsbbrZWD7AKLJZY58P34xtpXxwe8g7MegH7W8rVBzKpslF75eeHa7n7k+ZPj/J1rbUA7
FunCRYGXQyselHUv50pEZFABl188eJDuNKhk0/X7/YUFu7+WpnVbyyR/9VGlwdzfng9ju5V9seUm
O11nUEp0CAfpf45MEjBVwRQCyK6vGrKymQoA0ZiBBwzk8DiOK2X5AdCpAUM8p6+CtFG8Egqq046P
Vw2VSLJAhVz/ooOsRtPY+Ns80FPR4sBsk7MiJrHjRXlsmJhJ1FNAW85VftvJ+16gC6lGASuXUbca
wqGXxPeYViQu0ihC3U88Z0uDnBdcFU/ria3coJ8JnzuSUqz1fBlqWpdURAH+Mf4KHJGtQ8MBVsP2
XUFwDCHDNpmQfR7TvDHXc1EGzhlKyVqVJOWmbZW+vnWaBzj66XDyYN1uub/vnDcIyYINNrBPOyvR
T4Xyj5dRASxqRYbq+IfHsijTtx0LMdF/mKCd+WjQLobhYaUWYCUfxre5sD1ekMnJuRt+tt2Nj7gW
nKOaxC5wY2bE2JnzIe5SN2LSnyf3ZERQ+OmzOt+EPsJE4TU0gpt47TIMsmM3O0kyQSzMll69VmdE
EcwbZ1QXhSHlEz6fM/UV04Zn6d6BrxA5uTzWTB0ZUmRLZC0lzsoiBhZ4KG1Dql8hVD1blY43KAvR
dLsfyox+5eGKrPUTZHPlrZrSOO4SwHfts71RcntgEJIVcrhbLWGRmArZFlvCC13FYaldnyXI8Sx+
gPcqY408ODtqkcNgo8zu5dPAO/FBoQnBSu5D8/JeCX7oKfr/D+cKIuUpEwbJOjyxnoHq0w34gmTH
VtKz7mi9aeuOOTvOuA4PYy/PKqAUP4u0AidY6taBMjTS+iN4Bw34QsknToSpaeR906zvr2GHFnf3
AaKkAM9J47t73+ZEZNvCI00Iw+HN6WGHzse3tGJnkPA6b8gXflVnGUux0xXYQEmS1Hb7DVFTJVKa
k9EMrBfhusA1e2Ni0LrqWaPK02XkdpAy7ok7Ulv3+1VY/BK1hkpBhKVjSAktHo7W6E6gTqbmdM7W
74xzzi3t1gz66+BdMOAQstfEbKYG7BUdhyoYIqkIExBj2YTnkj9yu8Wm0rON1pXH18Secr9LQpVw
IPVGml8BPHH7ldHLxsv6aknc5qwBvSe7zzzfTU8zOB+rfOyxJH7jXUPdvVrNCIgJhh2Oewml5dtZ
/8RH1HU64NxtoKOMg/AU7K6rPg902WFgcmPh8gv42jhqJG9lk/v4R/bO8GpNkgtjeYny72Rpqmy7
g7NzvU/FcoQUITQ4jXfHKA4Tw3Bw5KhNs6PHBOJ12NX67tq/z9UvcocGB3gwkTdr4MYDXD5ZNG6W
XIwH/jtbEF64Mi9bIlg07pbVpDsL5UEDyDtjHCqFiWP1mJs3KZ56eFLOkgUNumNDYo5efcaIpoBG
ChB7fmwzEdz3L4/GpAfKUWHFhSeo/EA42kve4Tb8H0GRFlTvGzMW/YmtKytt2YUirFw5XtASloM7
YZlgCs4+exwX1FIQTG4GTsPR7h9UDZ2RkiZI/PoKZiF7s2MjgxPoKl/9FdTM+7cY+XEaf3YXtAts
JuQ07HkIUT+4GWmUQMkj63NvTjJ7gjsH4S28p6Fg09vzhH5I5a3MKKa0+U7k7EDs4PtGMAI4XiKM
K1I46ZPaQtCR1iy9NKxluboGhKrnnqAcLSx36cWTBKiqnYOFk/Q4J4ez/CQSr0T+v+4vL1sJ5snz
o5gYhMkpGvnVNz0qjlijCznNTOmwf5kQY94R72Aix9o64ru8Q1+SjvMeMxbnYFmmSNnbmT7gkjLR
Lz9rKuA0932Y75CpNbGMsHwWsOYFpOyoOMOtmaNqwXQg6MlHL0ue0fQNl+hHdWNak0d/xjX9G5T8
MbFUHhn4Z4hfrnbtoSWgT4VXWmXgiymAcdrq3yVUY7V6i4UcayrklEB5LD0kItQOkUuArYoqMVhy
BD0FdreN/Yr3MtvAKmX9XuT7k1+aI8Lavs2wTxv9jYnm1r4YOxmP6qDZMcbwURS31EENDQbY8iVU
HZE18aJLGTkb+nFkMsr+sAoG/5BGS7uEnSTPPXH9tGi8O5TXku9jXmTCP4fWBONyYmDojdJT91Fj
DR8l2UvhFNU/+bMmPZx0qW15+xGRBC2qLlUdxihiU1D4R+WMIzzAUN6hWGVzVBig0C+IJr7wBBv9
GZabrx5lymuL1yDrIxxkzH/EBJSAFVYUnNTVKgmbjWetoI6nOcwff03AYhZrN47DYOIgMRCoRbRv
vXRLH2Tcy0oNDkvx41AgKY5JVu+iIFRNeDNRd7AKppTnxCAqz6GAH3F7n1WWfHm1eewf1YHG9Lib
lMw6B0jf0ymDkh78SSmcAhjfBRGGPI/KaH8fZwJ0tJoGCsxKl0hODNEnW6kN+2AZEAC344Q+ihI0
tZ1WC53hC+sfuyYw/tfwLP5d551ey1jlFZljABXumbynrgmhuB/RCyefAqEkzalVTXHvPtmmuwWh
zFrGKw4uD2Y93/iI0flPPU6rmLkk3m6ogrGkcdTf4XNyHDGFa6OYhXeTZSj4VZyHPd3Q8CzXEN1Y
sSVbP9EwhZC+0HxtDrERG5IT6STwbtutVQzdyyNeeEQh8mAhKM7kVXgamjKf4cBdpFfWYN709iQf
726I6pBYA9NEdEs41QX79ZBLBCujE0NmtuDSpNlUfItUOwB4Mf22ZV9HuhCxfo0uR6MJs+6NWo8u
s5MLUdomu4he9yYLPUxrCtbVgXJuBDmn2xSpNxQ9rovXYFk9lmk4B49veC0ydq63jTtItp0A+YQZ
aJbjtkp1Tl8HzNoQuYJOls1dKXh0DXOcsiB7Tp+T1yXfKajjN0sYUuBFWwy4YPdyWNmPU9f9LXJr
ei4mn/JHKpGaKyoCMogC6UFwUfP20R2lQj39cI3st+4GN2iKShq6hi/b3+SVgRIXqRTMFMe6/mQ4
ofghbJ0IdfKXODoGO3eNpvHcGDgjWWjgsfLPJeoaODDGQaHlidq92+gUeYeq++eEUCtNIdR43DTs
8HOSR8INmhTCJ+6b13QF6Vo24F75LlakzfJT6/bOSC4Eu9Z73n1yXvaLtAYuxYwTV1Q9Qg7XkTrv
OclGx/F7xcWcmAVrQUPwN3k/knkxVwxNPdPI40Bax947woG775ZERfVSFcAyuvRZRg5Te7dFw+GY
051GTkfeeUzWV3zAI4YtRhQSCRBM4LHiroGkl4r7LLmRr5dpt+HDtcUOO83yNS2xDAIhL7kDdnvK
lPSeyA2Wfv/bB04+kmgOcw2nK9JHmn2sq2CDJb6OxrTzgUKAwU8IhCqygZiuq4JgdcP3b3H18dNX
Mcur4bzhlNiswKSEoTeLQ9wukHymOo+evTIc0pMfftag4JSAaQd+DQ+1V7kelSR5w2bTKWz4heQY
QmnIzY1lxA1cc6IE3rxX9PohqRoATyy4PZjZr71dXK/U7ZDUbDMUyq8roJUxKoLBitr1w8YLsyB+
0oNMeJPQAta14Y8tZR9sMSBPiToFlaCxV174PIamD8OQHNnIojgwCPOxLjcO9VoURLWa1FjCC90z
A/j/anl+NgovT46XAKa4m5nYP82PALU2GDDPjLukSqr0UMrMuUEZO7QqKIqWy5C4CsZq1dXIL/ED
rIMU9T4rhj+GJCoF5TofJXFTDfQinUlddcrBV6Uw1pNy7ox/GDjGTg9MzQzjc9EoJUL2anll8Xf5
xkP4Mu869lVMP7XRrrb3EzZzgsa+iKfgUfF42dZ9jZG1s1aRMXBoplNZUEeXhBZhAs3pB5EdR7Al
cP2fBUDT9JAMeII4dvE2BXwKmIJOrZQ9KiZCk9XEj8DuedExm/mOoTClwtEotibfT5f6XQRtOYmH
bW25+VZof5qW/R9LUZMKAztwhkBNzH1P1eQiCSCkz100LXP16OZNoB93AsdT4qn9cRXbZtwJHkF3
ZaoghrMv7yvVzbUbF283LeUhtfbtvgDH3Vi2WYWa2TGfpB7wE7WcExIDUVDUVl9nSM6IygzaZD/6
BRK7qsgyLYFQgnIgCfFR1glVcZskFxCfTrpmhDYhTKLN+th0HEA9aQ/zDJyxH48HpmRn/HEPfPt+
mLhmdMhOTSgWWrYSDuLpHJzs7zu7C7EhJj/IvUbSKySdz6aQ39XTrT1Thq1glMyfxgD+sZ4SWHm0
BuM32e+w/Uw1OPVKkDFHQiOssEx5Xf+HsOTiquim87Rc5T/J+pSFHulLx/NJ2246NcHQz9GlmwVL
63znN75+RWQgB+n8ptH3p/YYJrvOYkht/bOEEWTA0mfH4VTwqrN22k2jMEKnXanJXx9n8Zz1Y5Dh
356EVmAc800Dq9ArBKTaQLundH1fckG1mJIYidlWhFyPE2C4jlTl9Qw3rm47S1XkPLh4WjSS+9Rz
AaziorygVjt3snryZl7Wt8Bi8q6qTyZHi3As7NPFHpB9SZcwr5bvXrHHEPpWRhu20jAiOMagvHSG
C1VV5Z0OxVj1Ylb1tk9GD5aLe5wp36mqQ0W7flshbsSF9xXQTDL8uD2Enqy7sxxSFajQQefu1Kgo
nJoz7u7Rcwigi9TiL0qwuLbWse0Nsc6rTZkMWaEAqnNAdmDwSn1TkertGeXuQNSqGcNVgkhkcmTv
XUK9Z1zGsbXZCP1Ims8G1aVRMLfhFbR6PXmseAIHeawYGzoMQIv8jsQtO+zZ4FigIf+9o07EOglr
fbwoGrAUP/KqOb8tvSlZVHR2Uay8Hb2d/1J19UsHpyKVhl4z0aD0xvecfiUPo8VS0bUoyY0PvzUz
U2NQ7Hp8fnmoAMl5XLuaJY483OFo3OBfZRVdjoEtAYnIKZ/HMWS9omDpVT7cPP3r/kbEqRkfD5zB
TgjYaP+hpr0e9PxVNvgArIhHxEFcZTlp96Noq2K5qbOdvS5x/PcGr14lveMfJ4d9l/EVv27bCL0J
Gip8j/20s6LRnbpTB2je97w/qsAxd+QapafAov1iMjkKCISDkPZZCIJngBnJa8eHcxqGsmyenAIZ
AbC5ugXl/2UCE1x8J8wphRJadzRkXTSZipcwJM+ZTlEGzbWfcQI1gCEm6WhEhDneIIt2ZvDr3BB+
qtN/nGRkbvl1aAL5kQTFka1e+Of3NSY4TzZzGRoF7XKN3VxRjA/pdE1Q6LPKg+FMIluXJqM+sYNu
4nszUCiWzWVvi2FLKzvusuOjFVbzH/D95+JAoqJP5ENejTHiVR8MGYt8x1Hz+w1KHEpC6PTmD7DF
yn234wzqBFgde42/2dIPXP0AW2Nz40MJmgJRB1QdPT5VECztUGVUwsouXf8RrBwXksod8TpkYZxl
IVV+bWFqFiHxsJDvqdLv+V3npXjh6+zEZDtIq2c2sMWLfWPl/aH1I/TAgioVtBTnCTFwaikQnvYN
G0n6/u7BUwLr6FkgZEzfgJiK/lnOaXiT+e4VxCyaOo+gJobz5IL+S5qaiWlBCqxupTu1zHBW3QHv
wOmbzSq7UvW+yuUU9O9GVlEYZ7vBpGbIh5KLt2Vx15OPnAEFvJn5r74HXeZYANzCcFnJH8t4j53s
/RQe74M30JnpPjri/P45CgAy5tbwg5uiWyWbru2FviwqhsiIt/92lnd/yh1K+5nSiHkGlKXJ1g+i
FZCOSrfQxsnda6O1fHc49wOR1uZnJm1SsaPgr4jq9sciOkZVc9uUQG5xTiYrjn2yVY6MTUculadI
C4g/gsOtOUr/elcPUgPNIbL2vpd7yXziL87PzHHjJwWp6Y+gPSxDsvdUnPiBDVTdQYs1Y+saQLw/
YxEIwfVL3hsWfkKvGIe9pk5ISVN+ppIVQTpkYZFGCy/3OdA3UCNpHsdG41We+fLwRW73HqngXVNG
SbZGAqdjJYuN/HuLmGS5g0vz+hP4oiHiHTifU6o+3bkHA5Ysbz+Dx+mEpLyJ8ouQoeXkM54/P3Pd
vqOGn1sLso1PqiAr6A4J2ltYTgkHv5oCWNCvWEqmXhr3BAGFjVNHSqlMGlvfdfwy8w+pJveS4Yqa
0LCaGf6BD75pGxO0OIT/0GR694eE6Y67woWT5EUpY0q5oWeMyq/4YdeR7OorXAXkZZAdOAYA1RG/
EizYjhK0+68rgaPCOAmyStn8G7oFQd78PDdyFyEMsS+VOaLgzG+HuJygLmT/LMKeKgajeHLBsFUD
cwClGxnr0Od8BS+LXBFxRpw/FK7zVrPKkqIoM/PzFce6YEiflNWNtdPkUJeCt9XJtSQ1CIRspcmx
hglfqUCBIHzV5On3eEndfFbbDS0+SjOQx7cXlQx5KyclKofyQmJ4SqobcLE0XgpRwd98M0XxID32
KaxqRPXsm330qw4LFQ+WcBh/FI8islgHNW5FCQOaU27cjKSqU9G7QzBylqXvkMBALAltYnMmLde2
MQoahyZc9L2EAeoMYhxHYBWBucYi6B8va9/Aa1anViKkL8NVsCC0TueQuylYlPEezGzQxhcJKU+w
F1qT5+5P2xaiCNQX5x6+lVCZeJ5SkrkjkXUgclBBy9uWC3s+wCjAi84jPTwSi3RFXP5LQQn5MmAA
BkbwGyA7wLB483bQZFGrQE/YWGinE0JUMt8H0z4v8N8zHWis7S+B/Hq2rjNkr5CQvsAAhclgqrVw
25dcwj9wpH445OtMLh9Q4kPuyRR+82fO8Hoqax7a6f19Py65olDXuVzxEus1mBC/PffCkCMii6ac
GoU4tgQbgBe4kEUUZY3WQfzkN0SDC7nX+mKX3JYtcE31drWbKKtYI6WKpCED/+PnL3dFDnnEjE2Z
nyf7Q3JshwGUQoEum+uKHLnzaF3p2rdGAecRw5p3/iOOeNtbsAE9Lu2QoLZbcRsfG45lttJnU4JW
h9ctL0M9INn5+bukAKthB/YIyYTbc/hZCfwJgC4DFeyBcVCwR/9Eb3eB7tfPn2JLhNkoNpudHjM8
VInA6VubwhzIY+NaK+Z4lt2Pd3fHjEs9iPLL5V354gIPHL7Ze9nQ4NxYtlkjkrrsFK8V0SBb8xrq
uOQRVO+RIMWpmTY8uHmKi7siHv92VuVqxW2Ywyg+kN543QmFWtzRxg95I2KWe1RtW0Wln0CI9t42
yFRll2CkNzAPKLp85b0VSfETHdQWgpLJI+9PnO3jge+fmRinYEREw6N2mecdNWM4qFw0g85+eIyI
W40/P0KagyVChgef4l6LfvMtNQlzXAB5iCfen7tkw4acc6v+hCQCBJRq5dQ6eNncJCV5i0lgKGfW
URTtcy2OOk9Bu9Ss3+QRp7YOlM1dEwXLwjSFppODixAWdIBPNtuC6LNMhBQBcDtnCsvpkJAmidjx
BZiX5kGa4c719gYcYOvuw7uMHMvQqAsNR0NDCAwCzMhkP4iwT8H1aOhzF1NhCokTmk95PbY2gNZI
twGytps/XUI/FtA/hQulJ2GLn1egCKhkPi5DV0tW1TMSm8uylUaZWIeOU7Y/iTZhgJRQzAR3XupZ
zKDLLIMUAtVXbjipLnBFKYUT4XQBU24DLgwUr57V67fkJcFmjbBDBLogPLrNZx5VxVqEq1a1tgNe
gg1mrL/BP9EhMayAzUHuGodEzOHjWpEel6pOuVAlxx7txfRX2E+PlfPzkse60nw61RKqDIIL7hm4
1XAAVu7Btd29nmf1KI00NqDBBXLB/r9anzdJnzrT+rFRiNJtbKtXzAAzDS1TOYa5grc7N1nI/bW0
vHlC/2IkAq7+PJewbbZ6BQNyuofVGIcITROtNkdv3YZdNz6Jc21HILzCWP0PD3fZjmifllHje2m+
DOxwunAbEIAagxIkxbHGWr06i5LzNYeCv7JFBxIvWZG9mKcYfPmIiJHKhO9mCuIJYL9av9Cvhpjn
8H9mjOaqdEVtypJwT0rqe7vpHLmj3xfV30bmpAm68G12kEnjZ8c26YHnFtrfbEyvMcx3yptxsAY9
WfC6dwnE7qV48zthVH/mjk5BpFEkjpkM4IgBjZ6mZmXNVx+zs6mrJ8EU+uW00GxnpdVhi8DaJ583
KRutTIMAuLZLpD7ws23FspbzdD5rnUNPHIWTSIGaCFQjOgU8TIrwtvu5v5q/OjExXX+Q0VOnUmGU
YSwwTnnZCKJiCe/sTt5ryavjn+abbe/3FH2bxzCm2C+B/gw3gb6tPuxmlMPfNkq9pG9hDlNPx3jf
ww43aoWo5tdRgCdZEtD9k/I4Hr4XhiC7pj8TLmZjFmtZXGzQTpFn2Ujd/bo7/dHA4vbkZWBm7lsu
cU7GLzX6n7K7XRhliV5VhdyKneAo3xvdYZiE2szF9Km62OiTBwx1xm1uH9TRdYLSMnhNSrxAZ9Ta
pxNGaDWFjS1sq+1zCdOeGNeUqQSKI7RRe6VEqF4yJlhdwzZ7IJDQO+0ZWcoYw0EeHBRUDqW4bfEp
xgdG+B5DwCIcVzCJ+1r1rjmI1p0ZAB7kKi45+SwRmkcOCGpue5XGgvu/c+13sT+M3PWaRmyxE0Ee
GT2ne5ONjieXGjxEww7AqwodFUph7vhtakSi+fIJpc9WC2Lm02BLmAuq+0ZG/q1a4IeQ3lLefKPZ
/q2i8+bdCDu1M0CD2BSjACqJ4QsYVu5wKRWo8YzlxKLavhG8e+aMs1cZTQrQV9FSy3k3yZ/TBwlf
SqVWFceisZgUBFCYzs6BNQL24zoPnTNC84jETmMa1rDnKUPw0eE+AEgrR68kP1sUwQYFmKZDj+bW
XarrCTFNWdRzFpTj4O77JpXg69zv/DlNIXkCIuYz/D9o7DjhMA0dfUEUb1eYuXkWSbLW+eEzYLUP
7iaYyLfkKTeTPrIM2Z30fI1sz5bE7wxBxNtqFNFVUd2WRk1iRm4ihSgD6hDII/plVUK03KJ4boLC
SZq942DpI7bHRgPsDHLeHEg3cc+BbyZEqifL1gJxFyKuoVmdyMs4jKA4bdlFw/43rOTu5cYq7J/7
tFGpjpae98Nti/boTEyRZtdn/0ugy576QvaSYO7Wg4LQDaat5xDlK7eUziNPbeV0sWoOX4kplk6t
fVGu00bvwSl3u2OMqhs5yuHrFeV9bVudknjxLCkALo8dAcbi2gNrXFGNnoid+wxtIJYnCVihUBag
VPJFhJJIVXHLQe6IrfdICDuZgByOhpEmrIm1AtgTE5M99SlnyWzdhB0mFFXd+n4Dr+8KM5E6Bmis
xPkC/oQhFmQzK6kdvVhCk26HEYpvkKzjt5e67E1yVhwmkJwsvtC2eO6X2MJOtTljq6gHS2XnVmqf
hUtwcewHA71+Hjx9P3kHjinHbW+S68Zawnp+1Q4sDtxuxieHA5wFcAq9ZWkl9eQFgN3J88E1qlxP
2rqHoF8Dy+3v9uQuQs/TDhoP4yCJOxJHRMr6e4cTtvYHmPyXC76e7LDijje3AN7x4Lz2zNdG06fj
qWsEkmO5hqvZznNtuB5+T8EvxMDMO+UaGnez7fEljWU8RoZDkL5iABgeYQwbWeC1R7cpSaxkOVcO
MiL6K1vFdBwFLZJfK9O/xA6M/wvL2zVtJ85qZSnZG4dVaCghPrC8dCHzqBM1x3dUaAYHA8SQYPXv
4hj/fJFX9z9aODGwz6KxUOwJ1JdGQ/JBAQ8/YBsEXmRgHX/2lTTNT2H6vA9+swqyasjFUTzIy+fo
vRTPom38h3nCH4Khy6ed6jVMy23AZY5doNgWaWD8DP2gne4oZNwSuKcAtHrcRSQAAcLbV2sZ5XeD
WRD5C1+U3uWezNZ6/JZxYAim7WxZulRk9l7bMvviZTScEtsktD2IDf1HvLyDiMfKJ53ZRrFkqUGp
eSbYdj4GDTbxMyKF4e6rEoXcXK8iuW7Sumr0kAJfFzFSW+1zzsIRAxAuQSPWWAgdw9DQm3hN+VG5
qu2oThymwoBP8aHEt0Vam1aFQpX13uQqJAIfxoinY42On6mgnECjJiVioa9LSp/yr7ugLeag6P0z
SppZMobZojZYg4/OP/oeHraqnkhhLPiJdYficn0K8grEAXO6514vpRGNSdaeYjX2ugNbGJjWdPqX
BMWXsUN+soAepHFiQuTrHeFKMd5ZOROpuWAypCxfPU0+dAmkXSXnnBX4CcJoCRAkwqnph/eMfA0E
HNCMnz04z9klfgIsSpz/C3hdsqDTOAv5SvA95ByYkKWSO3sQn3u4iTQNPkNv5ZoJUngIaFghQW00
3swa8u4prLH2cAKGUtnxQr9Y4WnLzaLMH2lm54FGd9t3xKDJIg01FU0hHRjxR99QhhYBmal0nknF
g2Xgffw5V2Sg7z8l8v/le4R1Na9oiVsasGEfLg3l7o0Pdw/pdhq6fFjvfR/+QF2f8sxDr9IQI1+e
j2uffKHWH6JpwOExE4h95P7ShdeB/pBlh6jV06TgawizJ5+3nfXDkkoR3+c+ahG+wjFvAMGdG13v
fEeO868X9T9om2k9AcXZn1Y/eB7ZoAaQukFrZD/a+cyBNY5fVY7lyI+Z5SjgfbTQSNB8tQVuYA85
j//7K0A6rheJzjka5J2eemQ2TXdfuBG+3ns5DS1/xly0kAPU7uSfh/BDHLymAEDa6rNTfQ9xyAdK
enjKKUej7njgXzN72A0ePz9FT2WCYFzE8WHsCmPQLIKMzXzjCCU7ky0AQvq/BEVeh3lFUbxTHb9O
AU8zMAlZkJ/Xo5H2fPpNIvtAxshGh+vV99godRXHkTLwNUxDi6zEneZiW96ynUnMyNM3Cpe5FClw
Srn7jbiWXWZsQXbhz9h+OOxq6WHevW5/Xz5+IbSYt/GpAFFWKHW+k/NIL6NhCloK7IgCSQV7GjiY
Cniw2lb4Zt4dhKhbwSMrGbDADNvUy9TJtsCT5ncOU+5A45tkTK6eLx3929H93e1l+ya5/a62MLLv
xqtLzBjQx+y2BS49y5n4eRR37xotHlS5wWKOTORCa1IElaahUI86umyHG7msLUTG5Uy8R/geW6xN
DW7X3pHRRi7yf6knPLG9qDMdw2mUdC8ScF4Rs0YoXLaxcR6vqYd8mhQ8LDKhmpIOkiliB1F2aQVd
HSZDznPn5q+zgQMtWiVdz74yG9vqFX1zNeJDkvKlqF5jTZ4HAHWSMIYCpIjKdUU3dZAb/hE/wydG
vAQiVW7t7nE1r8z6ZLJeupXFiAHJ+su1fVxVZOxyOWmlI43NAjq3WjZvUC9O7oyJ0Tcc2uRghMMd
poC4iyKzbg3AxHgJlfC7q94PcA9HUxWezQdhBi4oL2PuGWjAXmK+ToYnPjGCm300rUHwu2ENP8Bg
o+e48XjuireTazQ8yQd/HjJwoUV+C8kiWmoNkyKUqISoBthuuBiX0GjyE+DuO4TUy7rVf+0WMDF/
T3nP9AZy7rfhl9awYTUKeQYob+wRRdnxSRm4EgkWzxosFyA2e+69DuTvRaZ9CHE+eehNhIrGNY1U
OQOgBaiiDlcX5DCY35zAwdGW1cltBqG/kDHv4cGXrcybBHPrBcPwkzScyGd7ZEchJtewrnDx5RiT
JQZQMpb6VMTgerYyo5uGbxKVseXutCx0+0UkjV9/kYqoFBU/j5W3hs4c4pO42QxC0xzGVW0OXf6b
w0/ITVMa4J/8DO5JIf8K7BuuNKWE4IY4aNjvVwBGvEsXYDdoir3H530rXuRRj1wc4hg1kj8+368o
tRY0xH7EG5G3jI++zTeK9Ixs1Eb4Z5gU7GEPRdu9V+mNWTqf9pudeF2mn2jZ3HNe8tpw86FheSKH
tOKJWJUC7zUH4CrbX/beFYmX0YDr+XYCFJJqKV8rJqbje9m59suaO7v11dTNJlrVOvtQFiWa0HsR
2X5owel7C48XDvyxngipmMBG0CZGLbPwb+AdiUbLCgSlJA4h5Hd3Q10evZKhB6xP+Z9nz458bYpe
f1wgihdEvgKsCUjSEuX2ClV5GifH+13Wl7cHZy4ARVyNJicBEaghLPhH1JheqtQgof6gzLn5JkEs
oyUk1UgCRf4l0URQzGq8FxToVUtJosQNGoLCRB3bZFc99nAziKwYnoLxU/R5ZdCsfjpn6yPZGYfD
sUD31D9c8GVcYLJswa+kWL2QItjClR+jKIZFl1g/B6Q7excO3AsAAru9qN3h6N9/bw+vUHeeozg3
9GlzTTaWAgZfq/ZADLnI66pxRNAIZSCiFUczrEk7KOlC/Yo4PmI/Ei66IvUG5a0d2R/aOG/1Y3wJ
on3A9xDwOVRcORlua4mmUondNkDQ+yJAPgAZd85urDuveaTzFtFqtfv49MG0jjrKAEFvGc7/ao/a
c+H8/153TlGGezJVLrXXLyH1qVP5zMhmQZDcDIGhWQnH1EErVEx6SKAurrv2JO4+FnkHr5PFPW3m
kuRIMfyhbrm1iRWqSeXyICgwJ+ACm/PiEExSsy2LsaXgxe9vdY6EcJUKPWhJEr3IDLpNfXzS3wfX
Wu0/xhj5Ps49RDePsWJfBynt6WAI0B64rG5PBNCFe5TRXE0izZgVKsTgMsmR3C0GEm8yqKRour7v
oeTwAtBI4QhvqHMRO9PViDZHSYO2K14YjGHOE/JPXt3tdPlK0s7tIkawa3ozJxCTtJ3jjlNnGgIV
zkf8dmurOUfOepVNPDld/fYqX8DL5wwuIGia/tdKXOKNxcJKBEM7stlQeJEoSiPqyeZacS1fQx7l
9Jfh6Sm6u+4XouJYEMMpia960JC5qPFNmXRsa4uXJCb9Fz4WO0I0OkbrhV4H4SafRUEk4FtwhwdO
Llytlf4GxdlYSn1py3n6nlsovJoT5dxwrLlnxOY8hy3eDau9GYclz02KtaWFt7h8ume6oDN83AOX
fu7+N+7fD3CEHazqDvHIQVdKAVQGGQ34fNsfLTMRjv3WoHx2tqyFl3WEcytmWn6kvKQA74y3jsSx
h5A+3NJ/yeSCOobXQjoDnEh/pfe0N9SdLIQ8GpnV6B/ZYFcS7zMzP5dn1E8EMUWFCjq9tDueDHWw
3UBiDg7Ns+DD+jD8zJfpbnTvxDAxVV98wowanjFx255A4x5YQRpiB0XY7QmQth1E18cAxObfUvxE
gbbj+lGstYgOT21Qw0rncS4J9kXPrc4HUSyojGx2gQPj1mwd7+w7XyjaDRWbn9tfO+IsN2q60f5k
Wq+LYeowNheQn0/cAMbAIt71mp8WRw4cPk+UkZCjy+XRhByjw9lMAC2yYxEZzaRNfRAE5nahp27o
IDwVVdx6+c7KW4WbyH60pbXugCl6NYK5g9O+F2XI2AFyr6lG99zuVuLJ1yjM2+tFfpn5D9IUJ7xk
v0pj2LnTdeV+rlzhmGTBoRUkVFKL4lO3MC6B0DxPfraYHngW80vVnwLBiY8SB2AZWTEzbNhA3aZo
xojnieA1J5g1TaG1mPhbHQolkvdS7X+43WJnYzuPsc+dP8a18dKaLHR8osAuspIaPSBINW+h+PYP
5cYECLmLRFm3W9R8vcEtaY9PCYjger/Yc8RZNA1bp2novFaG6Pkw3RQCtDIBwWrmYONhX75+7FkI
4V7u+FgTLgM91tmMU1U/hfNx0qrOihNE+SGdQxLcsmcZXtBAUwERSg55pKSEkuQN3Y2C7XE2Mc7R
N2Krl0TlpHq1S/Qnyxtqxac4pWh4P9GyWWD1J85N6AsEWv1wZNlUg7ZkeAc1UTJRlnqlykaxSGET
Ffhxhiy9xYNKcWYpMjUI1Xz3gofIBRU9nlEjs7bEgdFnHumbhP5BRHnd9RXe+cf9DzKLyp5mvlL1
FL5c4zWHT1oaAOXLLJs8iea7GcZUZPHCI7nZP1ComHNzEA8YxJf48X5uQOCvLjVSIOaMvwqeFE2H
/HqVKnDBPbYmj8teKYHS187IJapxs2Cxge9/4UGc/X1EaWQmBrGJyp7Mscs3c40PEeG3ghLY79vq
4azCdFhLxNBIoxzPasmIyqNvlvXjsWCiDYILIwpA0nP6SLwpFoBjHIXb2HBuT6Lh5/mHSF0ysskE
M2KHwhCeCDz/zWmYd/nyUUePFM+S88RNVh0r4tzEt0ay+XrLWaUBiyq9Wzcury7qbmBpGSuMoEl5
uuw0d0Cle3gy7WFrLt+TrVKvpW5GGZZ58sGhUoKoH9RAzZqiXuHIoRZHZMRBTtWIJryDAlfWOevj
g2rAJkHESX+pMdG0Hsn0EYegVn59P1GRH5HInZ+Dm6s75ilQAdr77HeRDmuX6ZbBq0fODyJJxfp5
1mr3XQLcpL03JAhamRbMuTl5VHdWXdxReMgSKJNA9k6H59T3mSVefUUJz9OY7PsNGdtW6H2TwqoL
XWm8Vkv0xlS7QTRJj807+UCCvVckCj0/yQPQytDTzjLHkU2K460LGyrUPFONshSAQjjwCbj5D2wD
+5gqtMPFajNCc7AnS/letXQcS53Lmmnpj/JVyxlBecavb3acY9sZI2znyLajv+elDt9WrAzKTmw6
sIy1JppobzsnfDF3mZUgdpgUrCuJPK6bxzXhv3foV1T7nLRR/AqMISbup5YQ0aKzpT8DtqChVTcL
OZcn0kVeVhIRWez/JES+fTmUmkmXT2Zg1pj/sHyJxUHKmg5wa4mjcPuVkOX68+dJkiO0wSj/pAR2
Zr+AT3rSfWs6ZwJGI5zhrAXOq/la0bIjfbNITlaTT4buhgHTXjIrQmjbXd1D0Fi2KaAQszDvJxh0
cV4u85/m/A44YzpF12W3iDfHAsXw6UrP/vO1CMW+iC03dkOwvAhqhPa6GJikhD60lTe2zouejPYH
SbDLnNOu/gS/TLBnPKbfBkYmM8AiRmyVs2s0rb+ArzLK9TsLJaLvgGAGJEER0QQJjz1SAHSQzz5A
GD4UWf2VyR0rk2V4u84Fr2QVi7b6DMsU0SSCNTwJAWaIGkOu3H60o9k/Nj0CeFWb9A3agd/ccZ9n
NeP0nLeXHm6CXdM8bDv3/rCtmN3nJtt9IId+P8Cs4cKOwuCDBvewuHYS5mj/ioOV4uHfn6wgoahv
yfrSYy5GT59OZlAVTYPxGdqNz7JNpJadMRohKYdJLUs1njOjyj+MgzpcL2S6lJMzjX3+nmjHu7rf
K7kyLCQXS8tqv6Tf+RO3N/PETaBIGBbSeTH2EyUoDnoNEBWTBeY38SmDVJ52udXJJCaiX/Cbluu7
CAch72HK0XitKWhKrqfTN8Wb0m/HOJ8ykRsSI+wARXd7A1TL6Ujh12cp+pH0yP0SiKOTUjBqJMAs
utpTyPZpQxkJ9ljCnXV9aiLaSmU8uHTeG7X82d6r0ivZLT0LznioT+zLtE/qLMpBEK6jfHlId0Aj
E2gWWB5+NKehjcAEtKKW6yBAC4WggsHckLmjdTr0B59KzQI4WFts7M/RfkdcCLnNoDH7TGKCfxf8
tJIwfUxxajMUoarKYZuwyEB+9ScFneyfuXpBRPbRhjHZC1CjfKFwAiSCkF/CkB0V3vJOHf+jjP8V
7HyUFy5vwRWUemuQ6srSU9sTrGWY8B2I7GvJ9Mj87ZBeZ7qm8jBZK6IvHpTH8jGV7oIVkFIdHAXq
lZMnWdn0VtCcG/NsUFDQzqlOY7d92iDlNUDD9jFoCo/mkD8zeDBtduY/swW9Uc+bNSXTJRhZvuFU
N1RbRZR6PKSVfqBMHtLmpGW5bXd4zU+j2uXPauSd1lg2moqk9P/1KRQ/VrQ78fISpvKzvqu6qE+6
UWesIylrt0tvk4Xb4LQa68uCWH4MyVtyFejhFDacVf2KSWnZ1ny5wTFKdpyeXFEuVUjEaSq9xFwc
2Dh/t0/OiPtdaP98GRLoTibPoxdkWIHZyZavAa89c7gzfglUCMTyE+kxrArZEbeAZBeAHyJwmI/L
1nq/knZsIs3Ct99aFWCPF9CxhYUd+QB6w6+xTY4hewm0zDgJyvB1yAZ7+xWJIykiVIse2Vuw2iqC
rzmnVRpu+BFVzXRzQiuWzL8JwNREXAg1r5OGveDVZ0mxt/fjIkn/AhHe30WZOXIpKv/TDqWAk18+
7nwXZjm5HUxH1Y1CoXydXFc9khsStsUt0jQnn8SySxmhFgWIUARuugfI68egJcmgaYIB9D5JvDQc
IaQ6lVLamFe8dU0Bl6L2byGqOvX8vVIdt8OGpqBh5pMihjWlJHXlzXgVrcxNknzjCSGAi5L4K61n
du5GOrQGy+K2xh10BvOwmuU78/a2uOJjElEA3OF2l1bUegWEGpT801tKC7YG1exHYUOoNlBkhesp
+UNCmoyNhPHPu+oQLJGBw909gbFxt1Z1OBwWnNbS4yL/t5xzg4rk7tjHnkVi26tDYJOtzGFyc67V
LsFTwjDgV0azKC9qUxmUvMHxZZyFb34KBa7Ag/0gc1XohqhY6rts3QMa7mRdWZywM4Nh63WF4Bvn
yEUZXgL7dmCGKcO1rRu/EIU6GV3qhqI2oKXLvQbG99ansOMleqD4oZh+Vz3Tq4YGRgvwhI0tvMwL
4wPiFUR5ziqKT2phNcDT2Otn1BAZuiYRXnk8GAhjLNXxFxiKrw2lfB2gVEoPagmyNnOPHcVDdbxU
4BzYzsWLeas3yefg3HytyFHIia+cdHTdM0QW9OPa2dK8ir43JcYxXsMmrs4U96jkICy26z+Pq3kR
NUamrW9aSJ3Mj4TXqEzKx5pDrBxOMsXjMmUNWrqTouXH1vVn7OhaZPMT9l6i6OLWUhaaJmttZ4gT
WX1KHpbRhRaEU6vVc9T90TpXRc+VhjYvgQwdqcGVY7/yQ5Mz9SQDAWn4kBu25s2DVTkv/Vibq48n
WGydLx/wHShHtv56Zihk67WhOsX5CsoUSglu6eMvissX4e3hRng/8cCpIn4EEEDt6qVFtn1RDlI1
FjxXFIxl7eKGhoL/hTMlZ3fePpqo70FyTSSSA019n69s61ztLM3GMerXqAXVDAn6JtOL/3o5Lr6Z
s0YG9oFt5NmfM0oyjfmSy8K5YbWXWM4K7y/XqiZRBdGHPk4egvbSdw66jOb4ox4b0Zd3p0XHGlcd
X9PMfSYafeLyVun+kJ2pQNLj2UkLzTcbCK/pR+cdFJFNxXEK5ICI3bQkYBkFHq/IPYD8krrVzz2q
KGOoNzpvWnR3f7JtR9v7xUaQMdd2lAMcxiRSzBVJWYSe7wCEl3omc1NaxLsUowV3EjNJX6tAME5Z
1AEZCsHsf1NSc8sURB+w0YV5/cFhmN71+DYxed0L8WZY7MElUZyvwyE4HRz6gyncHxghCVBjrdQ2
fVSrXRzfWkP7dy2b99MdFkLRteOYM4S6NAz9oRWRSAsZ/XlfA2hf1E5+Da61nkv4BwcFKqnrBHyF
ttbUd1+toe5zlK6KTVXtOSeZn70eOPZJg7N+6IfjQy0yvHbV1DvDosyDlPLtj/GKzEuPpTbziyf6
zacYD2bWVVDpv4PYqQWV1rd35IFoYauMLA6eNGvhyH52KfC2gFaUcYLkP6OSqGv8i8tNf1HrK7Oh
0wLwh+tMDXpY2bXBSdPn+R8SSp+hNXijG+ElTMWgjB3T1F7d68l4AaojiK/WourQkVVndn7ksX0D
Ha/u2pzNPxl7uFG2X7DD0Q3vbBpI5kAlT/TSirGxohh+/EMhMS7+gLJWvMs9euasrZhTkAr0Wr2e
cLRGAzaKLINSCwRaInoO8Ei2ONdNNyb0EoUH31Q5+pzviil+KA8ysna9y8EkAdWdHDuF1fJ0NkVc
nN0s1r5jXIDYmYfRRyvSyMNzD+AupZFam4lqbRAQwD/rGyMYZQe3qF9Bi7Ai9rn6hlvnDyA3WyFL
CWLsf9g5EjfwFDpZhJyTFfXIdJCsLTrPcVBNWtG8DzNRVDCznHJPmoUldDKfPZSLREqyto8tiT8x
AMsSJ/1BPZsOhU2lIG3PqihpBnDzR7FyHVUboqWrixq41pE4o09K6LhFCYN+wECH87J/b2a+0Wf5
tDbbQjL72ju+nC4OQdbs1c9QFN8820TTPAYz5PIvB/8PYvmYknn0XjWZ2An7/+tnYM5Ls1maf0yQ
bekDolqiDfzUluLNTCWRQlm3wGCbj5niaZqNRbPjHcRBaiDJfUdr2KoI2kltJycODJTFWe5O93Mi
xiv1naSPTjkIx8uuoCYRSslzKF94DQUgJXWUYJgUlmez9BC4UOq7jHfjASIQc0+t3ihqEmOkBKi/
vnf9X5rATSUQukl6gsk7TfTZ16rXOkt5dn9jqLvWIN3reBNXp5At2S2Y8rVfEXV0Fe4YtKva2bur
uL2V/Jvd69IK5k2HsFV9ArA0Y/iGWOX7/9g7LAenP2i37NRjJS2mhAPCM1N3k8dM+y3AHSGvUkSp
+/CykpsTjKKcn5Jo9IHsgjS+3ysmTNiYXYHunQ1wpti88DhpfkU0fEN5TJPOlRPJVGuCrNrXq3Wi
E/QINOe22rnHrhulwx1mMAEdi0DhFWVevZNXIEuV9g25vpdhFuPE4XIu4YLJRTY2/TLGnrjg07KG
Z+5oWHOTRd1hXWlcNI3ckk1gH/4Q9t0cK/837mmFsJMemfCEi9sWjOs+iMe9f2r520jMwM4W3SXT
jIl7yz+CdCj3/uaFgZAoaXAXklZ9SXB1f1PsffvUTrGvSxGnsouGCtM0kMV7zrcqxQUbczHsmM+w
tD7G3hk94rmRDS8B5lAgHjUI6ft3zxVdq3DtEVqnSw+YNDV9NsaxyDbM+bsy+DH+Z6chlVJVG5cM
VS78VtE47SE/QFp365kOWu9oaLwJFd5HDGrcgXFU9XJQCwxT91xdPwaN51jIdeYnQTi2tM8ESrjz
T7nfHCnomKXaJUxdIvJOHNNl5gR+U7ZedRC3R3RPdNMvOYHgQhZlXfDJQ7491npd6Xzdiuphtq18
ZsOvyMVhQUnUz0hfuwoHz/dciq3cEo/LpYHlao1Adh2Wn335/kz3TNaMWXj904Cg+sasVeoI2YnD
Sg/aZKt+hh3MY2nglObaF19kaNQFG7DKIZmaWSsxaqm59yD05c7pIUPC7LeK2oogw85LIpPWu068
gP8ovm7ERoDuL1BQd1eC70LY9HLr4+o0ZirgPs/1T6ZiQrz3s1+D1xC+K2mc7eS9iO8GtCQdQfYN
Lzz9yXHihWwUt3VJo8PA9/YcUNfEUQpCQELYM/p/gB6xuIYI+bBP7UPtjCigblGzJQC6mv78mwBQ
pzONZXfwA8XKcys91KC2HUpQZvsVB3Oi9q0eCHSMaeHgPQ7kyRqmpi7eNnD+uV46szfERhXT2zLr
nJN4feRD8OGi8PuozQ6BmJ2J0NXVCBstWbumSNJSCEbCH3pS9iDo+asTTUvlD9V6QXOHMYDr9nev
zi+PDVcLvDng3Ucl5C3+Gh7sJ9CaMAur0hX62tjndJDqLHsW3ca8kUen9ucG4QjmCv+QpTLxGxi8
iG28bIxPiZm2z30IwLsfTy5448YTdMfxTcFwuWx0VPMfQln+TRs7A5Q3apudyeo4IxIQfmjmm3Jo
VolDzj6LOogeOnWEUw+wlhveodovQ5hu6LlWIhCA0wzsPM6Lpl4CnN9TV7kaIOfTCJCJzPWBJ67U
KJg1sJTf3cFWFyJWBjNY7DiBB+eM6H0GruhmvAunbPwLdQa+g/Hi+BMHeS3hfbUaQrepMT2yBrvC
MIypsU62hUoAc/WJYhwuRIQWklkpoXAS+t4HBoG9u7VxuFrD+Q6rgvY1SWaGST23mCbTFT5058wr
Tg96cC1fykAY7Y8st5WtuX2WRxcO+ImI7KHFIDhdL/W3R1LgMQ/MjfHAjVAipa9IQIn0UhM55n24
xJc1XgMn8vj9tLm5i1xlyRSgZqOJr4OUqWs7LAkPSdIY3OAGmWwrtb6dmKhr2RNNh+f4/y6xP/4W
+vx0Yd9nu5NkMXQiF0ve/QwxBdlM0DGu8cUT6NblD/RHafz27ARiKg90nWnbiQI5Hs7V/U+lKIe6
kRqZdWf8NAC0S8xM9H1YXyJzpsVClRB4gGRKs57y2p0AMJRhuo/VUYUr7ZsdzQDkQiLzM/M8gfP+
FFcdSVaet6JDYUrQfMWjnW7+18MTP2todAR0UxDz2Al7Mxsdrg7TFNM0ECHP/jBcr6Rvv7U8hmDg
lAF2ccJl4UQtxvhQ8uzK/hLL8mvlHrSOVWClhLJmEFG+tYMCgIlTDnC3xaljZ3bbM2yaCCvH+jVY
CDdx+yc52/gp94Uy2o6b8skXKAvo0Mo3dkpBS0Ni00hKDoBivemcatoOG5PalA6uNOSKxNo9xFU0
xILL/HBeIglhj1SaKD901qxPcStHPiUw2E7CdfsOCxcxBRaNW1EcTnyTeU2GDXqiowbquTZeDcIN
TlkK1mf9JvmUSRRxXpi7g8u1PiCI2GIOHs25Qul/uEGDnuW+SoAl3bUXBed+EB7rFy5l47O9+zmU
YaMNVphp97Ei75GbHKFaBq5No161dWQFqe5RoPQJiJggFPQ1KEWm3MyoMcw0sOzgFyhajAw/0WTs
Q1siFUT0tTsxR7HTA7WSsVavLdku+yXL+rYCuM5aRBxLCkPFoKMNi58TEnRmVSYIhv2nNRNZZgdi
Nw4ZMDdpwfSf42bGloDV0dEPWjo4WK08PuwHrzVkA5PmXbmxzhEUeT+e5FglnTojqaTncingnu4i
f60Gq9QI8RRMdI/GUWUpGsNhd/Pj8/vycNDDwFGy6hGUyMxCu+Cc/atJl1/q+0wMPj61BmJKuWEI
IRjDWG7qkH5qEmhNM9E/l3M+b1FaFBMJR/jQnjCKpqEhF3KL86u6kokcOFpk4RSRymW9tMjMkG/m
Ucl63Gn4kweTdy4Mowwm9PB7XSfdSPLWciNAKBED7DF06vdtTWTp+gaVPi3kPGCjY7GaaWAFlIrF
WGo7AyiUvHqsKT65DmriGWpDm+r/BI3LXv6ZBhnkJHtWIgw9h927nHsvie3eAS2BcNnXCsPqAyiv
HcsuhlZ9IF45C5peU5Vwayjfg0sxd/XlM3rdw/wQOOnckR6c5bH/Akgw99L9OH3fzzWVZEhXIXz1
eb6++5ILRywevGpRFiy+yUCc2yls3cut1e7OzuzGUzZwqyyA9s4DzKF4N2+F2rKnhUsZ8rYhpjmI
/DVf6a5DociHWHOE55qAqreq6DbzYIzdccygvLHXvfb6fRzxhLGW0cn9y5kOhGEyaaeJZnaOYLtz
QwxGWPk0FYdohsSUG9Xd9iQp2b3dHo6fYpxVFW3VW2OAT0Sc0poJ+UEHBDZlHNaMQ8dsutjkS26I
Jl7KZBJQbox+l+QJOUeYUOhbUHLd3hcAu7y7ISs1e04xX6IxiGWP0NBXEz3EB1eZAvlrOoBY05Tg
m9tWmfnT2LkhGWG3RRjBSyw3v/HNxzoUUgYpwDo922MxPXFMaUh/UcbOLasIvZYWLhnxezJzR1JP
Bgqq20oI/+KB3f6YKVURDjeZ/6ruGouz/et9Mx2NZx3sXUV560egMkFuz282KCqoSOq0GO/NYQm0
TqghqM0Cc+l+Of846uQ8N/TrmO20GjK5KWcdDDvNgtvWh6xEArq6lpL/HGa4QAmNzka7WBgJUllM
jxPJ1+LUpqUQwwLNxkwsDdnB699nHBiJS0kpoVNRpw/+iSufh0JLO23d0wXeqzPe17gdXXQ3UIn+
/qwNxXnLLnPwYGm5V0nqdrH1rWp8ENahb2GPCotbflrLEOwXv0S5sSI9NS4PZYh7bpOaASUAY4Gq
7+f4btHL6SHqGdw/oqCtD8Ml7VqC/X7JtOC+1VWyhmsJWfKp1+9Sn+RmamJRhSZl/eOQgNfWaagP
mR67byzX/INo2BhqbLrVvGVPUus1DLBsfmpHqyjZS+q31Os/MD/uRQME+KMEoVcN+kB0fcE5iAUo
rK/d38CtijyWTVZ9HH+P9dThcSpshT4LfG+NkXboYwXT06Ay2b1a32jmFPaUM28JqJouZG6jjsQh
rzIcgnBk5ruS2EwKu+7gx0VdggkfoRC57UnqJ52K8oaP9UqemNysjfnfoLGpB40tWLxPE+Jry1/H
VMYKOrbro+Zy1If8k2XZo88x5/b0q65dPT7G4wjB+KMnF3lHaVvpexldBaVzudtxIlWK1zs+7gi/
ZaQE7ryxAlWUPStya4lugaHLLVQLZbHj1IO642CNnt/fI+1cgSsRmt48cNMEBKl842tMNHV0IeWY
Ez0cOYsfhqDtF1l57kaZ7JBNRqTzuzLr2dKZtxQ5eLbyWNTs2pH0onNx31e7F4JujPLmZ8DYLSNB
0wtQRekyD7J3Zz++hTBcfCbk5Vzt7/8S9SeL23i50g3devSMq7U0TVsrTXZSvYd/H5oQcd1A7YEz
J/IHcb9aivbLs2TzDYSlcDfuL0SWk0HufbzLj8XMVa35ZLfR13wbt9Tt1HxT/jKeBNqcCxSMGqp2
NzRQI2w0SYBIGdDndAntUYSESQUbR8YiJelP54UDtm4IH7BQK/5DbAu3Yzt39tS3Q1uTqK2Mm/Kg
avIW+wRK4um2xqRr0h5L5qZDzXre/Pukk++SESYDM1RYGyBgq/gU4nPLPFBtZ1VDMzvhv/n+nhE9
6BHPSUZ4wgUMlobfuwl/N9PKDTEr/0LaZBXJJRxKkYQ3BwY6u+5vnkt8mvaYNByi+gl6aUUdWiW9
UlBKS6rLmFLo8v37SBUi7DgWcfoIE7TQeOH4t9L7nYd+zH+qnD+09qeYgZOGFmpyNXmtxdqGjTfj
ZgWEdv7pxAXSScvPVKoOsfAVuVYhJHCAIJHnx4VEkmTf0tminmWPnmD7qU0dFttqKDszhAieIpiH
LrVX+s0q0ONagBdHVH1IrmzpJllHoU8BdT4w9tnqy9wj3B6dtaK4e2kLqQmf6k424DEHCwXXBkU8
SmdCKJv9bdDSpcAPP4n5Q18PQjjo5o6EaqphztJ6YgPtbO1w9Ggf7ho8kLCH5uo6gMaBaVHPk3u8
J1cO4QbYrPVoG2vp9vZrUD/RjZzi4QIsy8xasRLjoWJMoA1BHDLYO7I4S/I9r1iBJTXksRfar0du
zz6zuEyDCIxWvK2Jq7W4jmHgTMwvDliniyM/cn8b8GY61wHbBJorNOSf6XkcJClqOCxLB3Z3dobc
iJwpIVcRRb3FrVan7wPEGFxpZcynQXmIOCPbTdnP/GmG27fulDPlTVV9WU7EHOUNAJK4zgCwFTdl
OuaNvehnFP7KP7Q4hhAiZvSgsfYDMUo9EzLDw9ltfTsg9PAoycm2LPa1xU7HVEphcPqgfNJHelFu
67c+rwLdUlb3Rdj0/lUFfbz/nkILpBOQect2P9R4jWViavqKMSuMm+/X8db6cFwr4vvKNh5KNcWz
HQlbAmiI/+Wu4wLjESnovjpUbALf9muib0XLPBoNEcBVqPVYW15CE0KjKdy8gUUxzG7r26f5iM5Q
IUHl0zbdvVbVIdsZD3mfq4nEZoWx7KlsEGPKhlq381V64UdxwvUlyl8ViXbbiyZZChx+InVN0Se6
yw6SH2v9UCvPXXOkD/h+s/Z7T4SSka2jp5iikHDxLDFituWmxhf0pFquxJeIja73kRV+cOMAtvf2
/hjMRVcYLTSzN0PqmDKtiRuPu65Rs1U0OcHRMkpQ6O8DSjkfFjMZVPgTTSs6Ssq+FyjVETWE6MWD
zGqp2d3FaRxvejtadPeWyUfPXm43J9WwGxAKVEe6u8WNPZf+tN8v+9y3YM/VgxrVRCUEUPXUHJ57
SrMa70NDSAQDjdw8Q/rE/mVGqAQEkOuS/AWVi6SncMIpzRTxZk5RghLTIJiP2jDMPtAT3HlFh68R
5ZwNzlSs7sjeUMQh9rfAXsGUpOoDJSLBC/zHMtaPqm2CaVFFaUggimfmuv3aZmgHQ6MKuR2t2dLZ
eES9P7dXVsmjPeXeGI24tKgW2DCNAn28h2ggBrsYIQYOM64ifcRfzUIkSGMRaqRU/sfWQBzvl9ZZ
vlbA79yrKEcXAL0Ilz2vzRXVqIHX03CsPiVCSB7i79MS7Yc9VGJTyZoh1NyN8GUlkFkEoORrd8KV
LIif4qX4PtrSj+Sxma7gpdm8pVahVFCWmL+vXXbBJh52/ywm7Y+83ImWePK7i4qEhBbFKlCsa7on
qfaQNyf5h1QjuN5vlS6/RENQD4sfrxEUA+cv9pUq3+YSbKU3UkVRqE3bUoGs79jeLyTYJHbJ61md
+XtrTyENQAFAp+xsPHrqJ1jABqPPfXGqiRDP0vEnOLoFqHjUBw/skCc9fzSkZWwxZ2ZVZ0A56q1u
sHuk/veoYXPoDorOkaHuE0vBPHWgBpStCYx8PI8Sa7d2p3pR8x8jJ9ZTlINbcBsYUaJ9CFDBNFnE
vOuJtiAi+cJYf5R/eNgRrEB6SQrCQe9KlN5qISFJ0wYy84UUUsGarIceyZvG3T8swWowqKE2KUCn
0m7oEsLTGSAm6MFakk7yShzkoI60Cu069NIrHNp+T0Ws1WnsukamcyIlgVecaOpNUz1D815dKFz9
bKe/hCryT2b4aUMDy9OydulG8BCMRXE5CRanxbAE1RJcIBbRhW20uLuGHqJf1sZGFuSilRu8zDwb
1KQ+b7uLzq6vrPfTSNOY3pbrTnH9RD3W2z42mnuJn0kSVuTULHFB9QA25rN/SsBI0L3dP2J+zE1E
Jws/HAVotY+qlJW1inPIwWvVFmV4pj2VQG5X0b7uQEEECsQ0L2gl7pTPE+H4bh677BftAE0o2JNp
HBE+pTusgqwEUiY38LILUA/hsqNFwuVBWaW2vVevwelaJOCiOmLSxGSzXcbLAPY7TZf1IR2NRy5I
rzBA9pk7f/oT1KknWeqyIS4ZqwbbKlfb5217a7BnjgmrXHDvDILTlLgq0Oy4dPIuSN5tgq82OmPB
JbHExPUC44MXWXx9mbPCI+CJaPCoAeQ3PpO8Rq6RctGTjqb6kelB35meanw3sWxJ1oUhlaLTQ1Cv
58g+td1ScLImtzic7g3TZfL7xHB9vwlC9ejnCghHCubtKoUJ6GTrN32Zptm0u4acczNqr80Q1Gn9
5c3e2WmycS/vPnfCqsInvH2Agu9HvZV6TubJyrvqD7LWeeDdyZ057LVtnHiAgV0da4SRfHpWmPwL
dUW/jl3kYub83VesdlCjFUTCXn4GfC/8cAKJZTOUcT/t5bchFBDBFnMyICn9m2mY8irhYXTGitOR
ClWGEOVaVz5HfsR9pk/p6Rt7ufEl6OH4lDDjs2xVhVjGTq8L8hCYkdoYI6gsOWgQ8HudYREZpv/i
5j3BNlgbF6OQX6SXf9ZAL4LCrfBpfU3dbiYaB93ovodE30etyPqGOGSOPee3pbJdT+Cb7r1FTqvC
YZZQ8licSkbcrFTCGzt/d/9iNi+i3xHgFrtnEA84QPirhtwjIbiQg0AK0faDZ4lXHdRiaZUH2s3q
T89SiagQ50w4J8JEwyT9yYCQyBkccwxH2baWogz/rOqEtzySwUvBkq7Iu+VcLuwY/HwVm2LY2VKb
/C9+0yYrh5ATSX9qBTtMC6QBU3dNA4pjiyDuAepcVT0p8ogedyGpRCEi48WhCnrpCrvs8qjxDR3G
aNGsZwbiQbTwUqgc0oolgIO/s+DKkm5FPNaFHD0D0mzOJ1TMGasvrG9PfxC9IclSUEWpABwIqR1V
hKUSiZVlNZOi40ITTCbNRCRGgTO7sVKIRav4XwSsebJ1r8lGTYrpmAySgN+DUgAXAXZNi7/nvibC
gZRBqk2prkeOGkjnX/EIt8w3C6NXychJNt78FSMpMr2QXxs1lad77dT91XNfRs1f9ZCH0v6n0KvQ
ilm3ACwAgSGLF5ildHApL7RuAieza/6Uf20itzEgnh6BaYZyEpNCXWrvrLAf0udaSnFj+8N9mA7o
iiQyKd1suqdIL4UyWipnhicXW5ZH8j/HxgpcP+87Q1FzxhsHuddOg0BN9upsrBjwylbAZJ2o3wxM
RF+nbqis1RcVQqTLylj7pIdJRIZKDMvVesCatAX19D1d73gOijNo4sLlzwBE5GykQSlYY48M5Wtz
/qY6nMhk0XWt4KG5HhudcKSXfAQIklDfzqtvwBEQZhVtjfkT9yFbyTcONJAAJosoxD1faSSt1lD2
2pD0ROfau0StFy58rD8UlUFms/83eQkz9VZhdb4AApCw5sc9TQWdaEbsHSpEJxB9L5i4ASEjozEK
CkwrVQpzuJQAH7a6NQoUHQFRpYTpK0T0ItKGW/ES4wqYhiJpsrcuP5/mGvJRYyVyyVHXE4GcI8nZ
uENEr8WNOT5RtNgYeLz1ju7CHFh0VIKLA7sRgtzg0GSz3WckCDNBJjk5+ttEHBm3Wzbz27bzlLOO
V7UYkH23p+NXrZ+866AerbQ2QRGHvpqvKnF06CvDkL0Z2W4otKKA/gErGhnm9PqDBwkvFYoMasHK
+MhPnK96QkVOC5cQ9bog8gxGCCmO9k5cFe6XfrsYcDkw8YUxnrvQeCm2BDNTyYvg32YPo1h13hEi
+yAQaBM0y6Afe5HMcfMONv8RnsVVhLFXeNn5Z7zQQr9zdZJdUVMVp4OVNXg8RbahrmBqcjEfyj8u
HWkSX0d67x9gy83WEOz0rZhqddpnAAQR70tGpMZki/IJDRa1c6h8TKhPHjzpyQKY96C78k/cwnUc
TKWay7Eb6wkDNG4T2gfcR0+a2dst2itE5z8b9053bK8YXzs2xqlkMzeTuptIYc9fgL/77tkg8zge
bC7I7+d6nmysfFZibKrJntXZU5tLKjnVoUdRxAL1V6eI9F98gzF6rFb5ThGxmdHXTBNYWv1wwch+
lcLD/nLUn2DIMczHsYD7He+8WXWhapNylefgiOC9Cn8bFEki3d52EbRXIXpvzraQ4XvYGpy5JeJC
723tHccb6VW/9Tmb8T288GkliGN2EYxj2GRFWPswrcV5Yc+Pe3DDGw0JagI4pFAcGhnh4H83nDT3
NABT8BTObwU9rqPY6FM2QaE2DWhhp5+6Ez9WbTNvxB6OptQkOxBu/ng9J/NvuqdNSYIr4bQzJR/N
4E57ttup2v0hmtPW+ieAzCAb2UX6z6y13JKTdIDs3HxVCN8iA2MmzV78UHi4R2GQB9Pl0/aeGX8Y
gT8vuNG03TaXM7Uk/jHYxuh4vfy7AnR3+NfNh6i5v9f0tHHX2k9OGCytxdQYxioTce2ADkcB28JB
3pVVEsBdiroVOIX6i00xDwEJRDbjAUGIy7Ubn0/iTcJlN8/7yqB4kqCWbmf4l0/OcsmcJVbBZtZV
S7LzNg/SB591FGihRdCl2iMzUtp3bvq1s0YHh8+WnjFRgEfyMNtt67dHPfhQsPAYSjaYZodDBNWl
jAYv3kd0kTBjBqiZgJHBz4Elp1lSTdlNPIvCgrYXy0CKQoknS1rBoNOMW+6msAwc+WjsTzT3m1Xz
h5atvtChOl+mLvDGBUpoVBrSpWS8BggFIWSRLfjfzLPTJUDcHgf9BmDa+yxL/c+KuVD0nQ55vWOW
tFxceDXE7IzaDZJNgRHzBVIy6JUJsNCrQBlT7LynIebanI13PB1V8S+jN67BtVlSimvoLZeAgIBu
SXQBvTacYvFVdrQ8W4wKNyzFzNY/NoZPUZuH4yFCIX6ZYLGQZgwPPWwryuCbJ8usE3iQbDFcuvRp
W6VTZmo244QFpS96P2KAiYcjSjLG0GHO4xFBkQWsKbHFYEI2UTzSXKum7QR6tNb6MdXk9rlVq8UZ
DiHLJGu5L0IU456HEmw19ww9i9nWz+3lHZTDp3cvKZeoS3hj6E+dnd+srf5S2xCLWCi7nLH/OviB
2QJiAapAaYVGIg9/P2Tmk3FYK3VGlUE2v9YH6MohKLN23p7EnLMuzExw4nwwAMaCMrh5kX6Yu+QT
iUk0r4f2Y+RQqWvhfveIaAC/+p1nIWwZq4xyrZE3zB54eXKvUVnhRjBVaE41XKjcGgag2Zs30UZz
/aXYwCei+N6yzQTUhvy4rNhlR0nQGlmqZ4CDSBKLiar+O1t9b2hACuudDtJB57ArkJhjRXBJ/imQ
b8vGykiA7d2d97l+R8k1Q+SSh0qH+0RCdM7IT1ZBFuFAkOKB6e//Hd7VoyYwHt6CXDtAhCK/JQd6
urpzFEeMnQ3G1XRKMu27HakaLl4VUfQkGuRf+Azy7UAro7ZIVdd8LCwc3CGqpi9gSzA9kofWKAcp
ToOmdbp2WPU0nWk204cTUXlQ7Dg3Ve9tJKEqMY9NM3qNBMOO+ybSCnKhhU6iaAtiJqkJfyl6XlzS
Qf3YqcJrtp/NrPn96o9FeXNDhiDAz6OG6XVNUpIt4WyHlb/acerAeu1+OZ2tDLnu/NYAEd01YjQh
dQwLgfN3HD938PXZoHpTn+keDgq+oYYYPOYno+d4/hbExxBj+ERlTgySoF2k7bVjuaCcPWYUGppc
VtTnC2fYAQ1T/IxEvX07u8HW4HABNoVIolczq8hLPdqXby5jnoH9BHGPrGGtF3LNf6lCcJxr8lgn
2/lWj1kR3tBNTH/sLWPTyZAt7gWN2N2Su36IVmW5bG4ZLy/Wi+DawT4ghSI8t9DfDSFBe1SL9Kpv
U25BlRBNCsd93ooWR8Vy1oU1L1R0apeiTEe+fi8lCpFOg2ILxqLClLIKiAKp0lUGrJXIbfoVwK6W
TkjTgIRttCg+HjjlJIyZCcNOPDcOGLrTZnHbBzEczHAVyYsOSrRFQRVoaxn9SsAqvfaWkOManT8z
P1uTLxQ4rpkXYT24gItD0STig3HzShCRKnyOme3B4qe+t1hl2mxPGwiIhYlnCKOEedqRJhxI4n1r
iS8ZUTsyeCssnmfsTxZiVjVvQKSUmSz36yxP8i71wyCaRiI1c3eKecJK9gcbLzDLzfpg0A1L3RLT
izJynz+8brXXxCU7c+CqARsyEvp81CifTwErctbLx1wU6spQUvDNvK6faVTSojRR6om9CiWx4IpV
agACW+Dnq0LN4PckX1BdC5meNHZRvXpSdcBAkmJ5AvIPc3hDrpbmoWVTODD0Se0HkkzU703QMady
hukIBfPKudAZABJBEb3MbPI1Z0lz749br1bnGps6Nhj9DyCVy/g6FnbLR8wMbwrHiIWcFuR4zBpN
9VvWla6EdZ6JNC8Wz6G2BKorSIN0HG4Bo/CYa6eY6sqR+9oidxCDGg1wqDYjaQzGmp1n5t30nneC
/rN0L8EXp0pcgT6k52K+LJqEAdLeRTadpCnvPxNbNvZB1CnypnwI3gNWNR8aQ6ECvV5/IcnR58pu
O36aewjBOb20yygEM95C0QjovPB5n5ILVuBWyDWoXOBnZZyYd0XIUrkhFaVxUMCS/6x49jKkWSub
bi35iumbuJ+ygBc5d2WVskVtrGHt37+NPpE+5zqC05h2AsDl1oma6a3dN5gfMLb5LxsMq5bFH8du
6bh+cB1mYXx0oiFmguseosoXleuqUmqdVpaRu3an8Kl0AUT02u48nyPxujJmEc79Vxp9W0iV8IYt
0/dsTnzR+Gn0Ay5lu7lzaw6lN4vwkXCzz078LOoFSlzeOYSvXkNkqgnDpfE0pbH04erE2gls937Z
qSWsgwQRWljuOCcqiCHs43vLliB46/LuPYBedDaQK4f6HVF5J8+pUc54U3uNrupc37ZqjHmoigpq
6fonfbvY6CLYNNtCqScXwIEp+ani9udCxraMfL8O4Ii1V+ilzxgrzP+k2XxAY5tFQ4rNLHpD5xuJ
Ho1JadAcLJKRQeGq+Xn52deYHuFWOBKor3xGKcKDrZu257d02MVwtHdfUHOsYY75A9UAmAXEL4lE
/YepZqXO5VRjwSwso7GrFNZpXcU2jL6vKzUVgPvlrSoOwWzb0pTYBGxPSCNL4M2GDevMNFBIjdcE
gGMb4t96Bci5I3pLgFdM38zduKp+vQbLSlXweBaPUq2j21q+RhiLZqsFbSJxnXw4DW7tDj2wpQCO
IpxLD5smadJRy+EgmvtCoHuTNtRatGSP+H55jbUAvRSOcTAHYmjh9k64n8ljKpGVt+sB+2u5IU7j
UupKTTimwcMaCHxCqckZHHVhUQ7SFmdAL0KFGpkUbzzcM7cEXwG2f+5+hZR+B/ZskgFCA1tBKwfO
IYONAlCHwaOFJhDg51JpEkJaq46PkEnKydNcOK5wruT7i0za4GmnLu9LtclA22Vb7nMO/YONMydE
8KBCstxqSbI3bLmJNQuZVzCAGwlQshcKjM5V2jGpx1efM+h+XFTkTpTiykZEZvv2az4goD8/2iuz
L3rBlvJa0mD7nA6wpta/AAuk/zGIS9BaGH5CW1Te53UUhRvtjdWVHM3Ik+wM/abPHwKvHz422t9C
yvoVjQOANekOsTmnZC3aGq2YCEjb2qjBcpUHdPsGLyS2QFsStezaZzs88o59EiNZgng2/6ODfQQU
jkaUWo8lX86l7kMu5tUzhLvGRnA2GTBCJXyLPGKidYldZqoLKC2gB+OuUWzYG2I9c2W1PLXNk5bG
PeHS9TMJ/KQ/wXhcflWNZz+yCvvv2cTLl2Q8OlEgfmAxE6PfQmV226jYItUcp2sHe8KfL7lEaUQo
/N0mDO1myPRhgwDz1Cm5KO2f58LMI7SpcJ3JHY/WkHy1biXlqc6AzsfBBihchXKrhH9mA7FRNGvl
d+6kzilLDGJhk4zruAQYwNYAPyjaVslAXIdEbfY8sB7Fwv/7cNw3WU04xt782N4pinJpNHlgMsfW
vBh6mxVCA8cDbOm9hViNOIn6QH3WxqN8ibJwgRCU5XXUH3WQLspcuH+Q1c/bw51ejQnXbHFpbcWw
xRc9KuN1F/I/cbfF0iAwEBtlZOWRpL3aEQUtqsHl7bVW0R3ABdV7U3nMp1CcFHOSdXMRSOAy+vvw
iMCk47z1S/6CyNtdYuIauwahUsFqd+Ta1gTzYjc9UISAz8CAgUc/lBq8S5ROCQO3DdsJltkjTr5V
9Q0rbLiOmDMJ7Ob1eZzWbo0LgHd9CVuqEYoRcnbAEGBBueieWCQSVKZvPJ8AZmUHivvtNppyT0Oa
8e4rCaWRaioqjaGC7UyK3dYGwD0Cu+jqyIX18HClvSZ8Ph6WeDhPAEnN/i3byV1oo7QAeaQg9dvm
+QAEzbl9gL8t5SxIO7cmEJAotbmwEkTaS8l1BXMTUaGfe0G9dZFY3v5B6dQTVj9KWfYBZcC1u/Ml
5EhDiMHC0O1JDHt/Pm5CYUppjuZ5tYzVI2LVlj9FVso5E3TKETwsd3q0iOagNFnNHrKGpfte+bfq
jyb1BaUWr3/oxjgA/yjdrtaKABdrP2cqoomu45AxlhW0lgkFm+Zcgl7bBCAt4wg3IkunvaoE68YN
+GleGX4l3epdyvmFD8jtIiqs8OMYGoo0gdj3Cl06byHWVyd1lzBtOs/rHdZu3y/0p9a3fJvIvSeP
Uf+ONU682KMiPZaTmTObho5qGD7iwJC357jL+923fdEEglcUrs83j1UNoBBlGvIi+2+8wx6mlUOI
mzK24ijC0y35gx5Ecf427pGCJIU+oxaEpwqJvXYdnT5y2YKFIhRCFrYcbb0Qi8qeuZ2BtRP1B5KA
4XCMZYH3jv2xJ6kOKu02sW5t2MAneX29+Rl2AC5cq1G1gSs+LCf+h2FeELzsEiCvZ1Yg43bDzHeh
yf5dQHDzZuR/PKzmJfjRGridEi43KVMEh4ysQ408GoLLXN1gJFWrJqtaSWbmBHV/KDoV5KHYR2nq
IhFX1UrIJBOLn/aGIHeZgmp+UnMOfs5Zba/NIFIrAxGHpU/7ij2YkPy5B0SaSyR3JR2MCHm9Nh1s
YYbaFcMHuY2ZnnrORU2+cUd4QPovmGiVjOI5jAKMAz0RAVD07f+3yeB5gM8Y8Uz167rMLhfV1KvH
SPaZaunAMEYrbyU6udETA5WikuDa4V20ABzibeMosaRksJMvTxVoupdtSKqRmjQLOih2f+UT3FTm
OBnZxHxg57bwvmfqB6N8OPVnqZXzigZytwsbuhujH6wkLs/D+S6x/+oT9/RzQhQ3MkQll/iujxqB
mgqsvsUfU+hEDJnDqvfB5AdvJwt6rFwaIshZSkyrD/un8vgOKaUNrFIPSn9en8DN2eK2w4QxuIjG
N0P4iVxVJfHGvleCmjFICgge8+cEGKgLYpQfszX5gPNrWnVJyaZ7Ez6UXLUzUp28al2oZkiVIvnO
VNEFQbJ8ksdqN3Hp8vGDZmaNecRHmG6+Pjt/XLU5EO5OimzICrHyo1VP96Vcz3zz8Uqh4hdAEmBm
xmdqbzezlvXebCQu52ruNerHcgHF90ykykav4am0gTy7e4Ye300mquouRm4am6IzcqZyPdpCKmnI
lCd1QYX4iZyI+q9MqfsklFsKm0yHdBjeYbvnuvhrlybvruxhiiI0BzYKn67AkZ/ffurToYR4ZKWO
elKBK9AsxKPLaBAmWiKEMel/sWh8mV5SwQyjcO9eaP0CCzPNPwzVbYwzm4hqFbfxqwF/YvRDo+sA
XFrHxcPsRkxIUx6UzpAT/5fhMXQZXuq7hcfXctipG5nyOsav8vFX8Hehh0tHBtm876z8kpYEiHPF
Y52pfp3gwlGTmawTSurNlRbTVDhivRPH6MuOzGFLFcKTO6DA6sxSGMZGsN5BaQhlsULGw4ShCyv1
E694k+0UThNJRjUxcdWDr+Zw57fQTQ0slhHw7hMY8eAQ3juRS6JDrkuHLeiZBMLFUljvOFPfcZz5
NdCCu+iIIpt0StLhVHTjQn1nO8nrbVGeV2xRY5/tdhqAxjGD9wfqxH9EjjIr1pZGNANO3kx/v0uV
c4SGC8LpvVNKj0UmK2EWUu9yrMztR1ilFUZpvfCRrdQNwC1R+d7uVphBSsEXgnJYn7Kx55Ai25f+
1CEvTkrpame0xF1vgE1deHaH4njkDVCyp0H9oPufOkk1/tcARpuxrTOLvYHSkjIWQerENN/gAjHp
FThG2jktQRol8Gt5+9gA0KqSqCNvAWaB6roK0GW+bYP58YtVJCSyzgRlX+RKBanUOGUmRT6euzcF
dH5S/KnuwAFZLj2FqoMYq15XfgYbVghd+TjUBhoK8rK7lNtsBC1LnReVcZ1MnCWqvi0d+XVboGbw
zRTz9fuyuUIrEPgmPlxA+lOr++zmP+/cHZ6ypnYOVMMX0lmJiCBQmVEQTNbCF1y+IWm1DcCs/6lw
2ujWSNwTStY9r+hoaKzLW1RaWMytsyuogzTFLFlSbTAxJyXux52+D9PRy1pRHuCReHEXFjB07ni2
/RcCSFDH+YR7B+a0GNRf8IgYnu4t05v2GebhggjmTemc8g/A0Z5IYXnVNN5XhEqcadhtLvjHKuh8
a6L0lPPkq7U2TgbPXUKvc45os2hxXX7MiAySaSUmliE+nppjpZ53oNd2uHtF/tJkdy4xfrekLfMS
8vcHWKa1BzJvhHgFh2MYGXL0w0CWqpN1dVAHm6Nhzoet0RsXalbWcAhqOwPMKX1IBorseEZpRMmQ
Nu6pJzo7EnW6oJSsu1QLbiNpBpTI6YAL9DCzwaC1Bmz8n1uh2PxpMTX6x8qCvqI5QFhGjIMbRcQv
ozg2HsSqZ4rYwEvo94BlWlRnWNWMyJqKq66L/8d4EEOrYEO99ZsmaA4UpUZcXdskKZ/DGHfZ90fe
/KyjOkGeMlvOLL0lshnCcS3g0tjMdbBMmW+UAEcrO1gJc0gbIIQPTCnbiRRsLFyt2R2q/MZaNiF3
/iEV4r2ZVyeA1dIeXYADvA0va73/pdsHD8jCE5xGN0RFsiCQtVl0DFdpWiqYoN45r0xFKPUQc0Qi
CwM/+gQ1ht2YJcfSft4AGS7Du7V0ka6R9nATxp5nf5TCZO24ZL7Ui0RUehNCM5hAqedZ52mJM5rB
5diepg6b91GEj0Vc7DKnj/1ZlmWRTfuLp1IjjyX1aw2vddV1oxjjNaXXEbObG20/yMaAOIxUTIzb
L1YW9ZkzyA8Vfc/9/8ndcds67LcC48UyfEHBm97HJNpIFBv5WWbou7RK5QBoDlhyU0+SVuG42eXc
rc037+gl/lMg/csMDVdW0fkVTutXwzwFrVDn2B3ORYJ+MR9+mn6MWmwgK8BFE+h2eFHfPNDkXikP
q2o3+Dgo8BoX/M52lzDpErSYcj2hAHdPF72Eb6uqXBEzwXvpLRp3MjUp0c/jEdU3HOqCZuR66oBP
fn9A1vdVnFAozL5X8I20XH816xL+RCGnhTbcvLW93FWgcjaj1NG2oLQmXAyaPYuXexlOWPGtJAPl
8sfUmzmFmSstBBFzvK6q7Eojnhx+YIOpMS31K4JXHlIEBp+TCoS+Wz9N68IZ8nkqsKDHI2gGcGPY
TxVisEblQn32opF+TEWHShTzahSEQii14VmKw+8YYeXoyx8jEyT0c8aOfeFao1hqJFM5sadASz+l
r+EY+h3xA74vMSfInrzD8LTN0OndENCElWxE5WrsjeE1p8WxWeaxXorcdvEUc0UzTX+OxRbHO8fk
p0H28DN0eSOAXQYB6kI3oPo0UoT00Tesd1YzXZI7kaLleMwpkd6JB6rVVN3aYVl7P2DlnUhrE07T
QBaNdw5tBfoK64YVs/cKAbVNBfRkRgXn9NGKqQJg8EAQsq+d4/uFIV2t4UbXcHmKqR1d2fQzVLIU
HYpXNjBhxAxQADJFNHRZ2QhHfKROzbZCsUgTEml6sUAcceO4R/dsycddDduU2lYpMgSjQCKRJ6bg
LddnHJuB8T8Q9syQgpFtXqCiWyyNzJZ+kCiMMAnyegl84BQKbtidteAhLrL6HeiEtcxUbaZj5Fbg
pN7Uyrk1YOogeC/GhphqSxgKRoIVTaFh9kQvpEFSOa/PZnwGYbLIDWr6rh3lRF2jAku8oCh4Cn2E
961mgPeJbkB5P8eHNzbPaJs+S2M49IIwVarDLLOzeIxBdIe0mxzASSF4x/+6xksEkGFRVX4fwz6b
YRcEWrNpXj3w2bxpGrvdueEePHnQ9CDRNWatA6/SOE9cooOUrKJDMXDSrJc3YIDiE4ncf5qAErTc
oAxWlgBsCHNxo5mMtK4zg2CiDVBX85FQYu4OAh0qvxCvfIaMRvuOebigGB9Bga5S+hpoOBXVNFlk
at5cJjGuikjNPLOK7Be4S73FrNABOTKXtmAOWnKn/H88PwT6OJeWEVwNE2IwsYl0xHcl2UwTZORo
Yvp1hd6bvpxtTFIaA/lbWmQLd8JlXGGcEk5Nsyc02m4VcuQTSz+AkPtba6ALxZVyhd1wEUJHQuen
d58N0qifoWMk03ukkVrqjIcuPiAG0mF0Dz3SbQGwNlECAr8MD1czjFHqUZ7h/jKyctFjWeKo7cRH
7rrP4Tu973EdSfgtQo+aoEP3TQP1H4EHXF8qeDDvSU+BHnrX2g6fPLI+MbyTSyjTPF4EVkioQ3lw
qjjJ3GRZXb7HYfh7f6ietCZwQL2qvbftAkNcLkpVx7NqhaX+wyEQIALJsfFs0f1NYA7mpUSvaHVK
qwxcLqf3GjFOGCJiYkYGkUNb0xa5KN+NduBKbuAwR2eqT+GlypII+E8vmEy/yXMriRzgKdxWxrji
6KVxaoItaXF3rFHrXpuWUHwTG11aInOvFQHQHmoXc2+E4ga2U+mieuJOUzkk+bm+dGSo7xZ2dQMU
9NDeS9bf0Q9BhhNGoAU7pW3NvJklzEa3u/AZl2SR8AYYpR219YDN8EJG9QQLJ0+JZIMoARQioN6w
5W2Q71ReKNueF1vC/Xao9qOlpRcNyFcQF8vTjw9EoueNmLfb+BtnB9UILhl71pr5W2Rv3os1JJ1h
ge3TkGU49LCsvM7FlooyAZxDFJarlXlmCoHlM0cg2W6ZR+WdnFpM0Yr23fJaGbRsendJvuNn8rm7
V8LxCMT7NX/xG+1UyZk3tRMSRCK/WAHBTfrJaL0xP+5b08hrDV72p03nerBxG8cMOO5p2AjhCloH
ew8Lseq8pLiiiaRbpUbpZfVBV+kG8HeQbpnnil+wxLp5OpoclK96lXy3mAPcfq7Q8ncqhff1t++n
RNd6nDvHO4yY0JixPJiV+4nRXsLkTv6n33TjeVU8hwrc2+ACvbP5b7LmWEYlLrdrN4iQ66A/Jj4G
TxIKe1IqSOkDP2TXK9lUoYSgPsG1cWKiYWH9XuWJbWB82EM1PsNzpREHcIxYsWKks3vWpnZd8Dpx
oL50+IfUH8mfyUqR7HxabLPbvXElBSTPOgA1urGBYId9zjdUcfdS7raSr3juFUJ+3x/02nMqeJua
eY47h9FFhKXl6dGx3tzba/0Ivlw1RL6vQJvBmsPt3nP/AxHYdXxMyHujjBoruB2gtEFcASxXbHzm
cTybvqNQxjOvjIFW2Y2qgp3VqdvD2joOnA9N1WVpPcR54oWc4cOfUbIAdLsLWgDD9FU7qdYo1Ryd
RqEkt2IeMMp7kro20OMtwfCxZ8buqf3EpWZETx2k+9+MdcTNWltRYzWnck0LINuqi2zM9Z7+CFUo
drOngABRCEoVr9g3vPfzZ9ukYD/Xu67p2CIH0e99eQEEU0w7ITojVGZMrS39NhglFS+Nj+Z4kROT
cLmK1u8744YbUpCXbFULMF5m3/3cgAHn06KdDtGaIuq3/zWh+jIb4cxfSutouIsL+UTGOIpyzdHq
uCwm6CrbCVaFWwqll8BY8txDuB21tQPUW95YXP/rAAJ24zL9aCieeNIo0shMoZOIhz3OfTpSmnVt
TcVxg4e6XWz7Ks1gWUVh91lby30GLXVqR0orlMDlZ3Qe3dMsmBwQD77Bt4KYs8qPtc5UXpBKZLL3
4FbEr4ylGBGJUUW/4BSNEJ/XQaRMt33/uCbq87bUR4eq8FuKN0sLwBkqBWgN3M//8GCXsMOFwMOj
ivA8ts8I+RQSkoMU/3jEyS3oCNTNudgg3Kw3njvsri8dGLlAP09561QmURCGY0iPuiFUW0Sga0tU
7ZP+TWIE+0fR1A+cIPzbP8YbClsJOq7TCMktN4TP2fCTC8I+Eju9cEbn9C+V0g3djNkubAy6fMpv
O4nPMMMnqQoaDlfZZk7fKVPrw7EWn0De8mMd4PkT5c0qXxhYE8OFeqDOvjDAA4bnAXdkdQjDgtp7
OkExfSRN8Dlukzfhe+SuML68zuJ01CK7qxiaeLYwnRe/yAb9y0Fj4o1nIf082OAGBCTvQGRsH/LF
yYCSz1nhgeMWgf5oV7V2yCHLHEJFiOtJHFAbfDE7LwW7B1HNFBXvP9kENuHkxaxH0lKjO6j85KIk
R91bnBR2KwVcqVZyADBqz9fgQXRL100vvxH0fCczNF5W43CWdr4j9OMa7WhLnFNUrnwCsWLEBrSk
IQgDGUiIWu+MTd+YICgt64AhwgdYgaSUDUPGsugWikR+OwjxskZ6Wpz1fN1LhrXr/9//qLA7D7gz
9R+S4NWx3AIUCw4BiAbz3hJm2yBMEC9y9JUwD6R19O/K50qyeDuhKi4zXEeBeYadhlhBCZhDbag2
qQ613wcHhJF7dnz788aIRthZfgfd1T1HlzLRrxJs6l0eQcxTBxxt9K2BBmg+6W8d9PVm2anrgvYd
GFmkSoKJKgjmGcpiOKJD4FxkD4U5bZGiexjlwlWHMSzfS5k2udLYplAu8BEHgyt5hhbO3Bn6BMjS
i++OJncwoUo5gk+W7/FIiL3aTjy0gn9AF1hT0LoVS/7DYKj5sGE09lBGdWk6E8X9+OKs6O4mYUEx
S2BXyokxJEC8fr5N47Gzbi3S5ys5Rx03rceeY4rjR/hKjepqqG7tjFxYiJtsIO/86cTLlQKBcr4I
fViAYDfh2mr7X7FnoYFqwLcvgalHtiN/rTZSs0lIdEMqgIhOm91vOezxO2KUgfGrYSRlKGuV5QEx
3d0MzpK0rMVtKh9pu1ztaoS5642up2/OVZXIGNWru62VeA5kcND7kJn9xQGk5JLlNQ7uXTiJmjOd
GGBH4z5MzrxKYcEf5a1UY9iQDpzsNkj8g45lENfAT7WQt7zK0uHQ9ZY8/okS71NvM8NE6rlts/k8
6N5njPfoogfcuBkvUz+gPSncBz1wbTrrt+bJa/YItS0yWSbsixaCPQG91iHdMVpFR/S7zFajkvqz
SzIuVQWnsc6R1PTejiJgqB1SKnCBaCrvhNrcZVtmXEHzQwtj5wIEUSt3vPguRSC0gpuyQHJYCZPN
YLrUmHPGDrX3q8KSlVlEFjLxXoqYOELRldC9BX6n3DsfR55lfUTvn/IZnj+S/wJOzMZHp47AV0MB
tvJhd5ier7qRUhxvgy562st4YwUcSj0hPJD+pHeKybD/1dpCQ/86X3g1iA+GX8Hz7GvwHPh7OpJz
agrb2OZbqT/7SoyVZclH+snFOHlqIXzsKUGi84Ux2iYxQFpARWt17bJQRLC24WVph0sEkGVmDWEJ
6ociwjmMnvPGczU/4BKSENWudDrCtDrSTiRITW6r6i/pXnpc+0lVC8pC1Meumvwg7R+KXdPd6gxP
SSLJxmDQ7Oe0XppgBbMJ2GvBqcAfvvZLqYt/hhDPszME6hHIVaYWLJcSHAaqE/+V3r0Rflnbm1Eu
2dLlKeoX+SOI+CnFp0OGzXCv5uAKeKt2dSZLlv9/aAsGnm1VMT7cxe67bZtBRVxNkTqDeeBjyv3z
GeCxwAbsZxiuouUwd4mij//2ipwbGDxrTwoz70RXfbDHEHJosI+XksVsKRz7YKmTlIjEswGw47S5
MMHkE3XGulqe4E7QzOxWNf3cdGIsmooAgczKb0gyvQpree2Wb6lYzJfChr9K1V1W+8D38HC0INpG
WgtyJ3J6H9LhC54B4VksgddOiWLT8Rr4GOja6pw/Mjycm0jLP2AeOC7MfFcRHVJmLKegqEpfB1GB
MQSbDD/93cuslACE+TlCl1kK+DdVhKdJjZU4SVOqTcELsA0yQ5GaTzEYZK1ZIcbEiUbRRhg512zl
k0n02weEPR+k1GqUZs/k3roq3knS7SOfS+aB47xPlbpCGZE6cAR4MPjOJStQx+EPK6P8AaZIoObD
Y4BKpXWUhBbMIGH7QJh1OK9v0cmMO0aAslh+TRGM3YGNL3YkAq/TXEvxRidzRGA2h8Wg7SqL/aAx
glwVvfRRF4BWt8kpgNzvh4QvaOuBktHj8AFldDsSHalvQzFebHG2jineBytN/fQldXdPyekzSZHA
8SWasZ+yDTRRuW/4F95oDIivb72KsH/jCDuWkagosLHPNcr9iRBTnz8VvK8dw7bi+MdElVP4gGOL
9dnZmp3eYiPk//t9z99sSE3k6sB7+TQa9sCFiEehf/mAsfOp9tV2PNlTaHpFE2RiTvYfaz3lksyy
5JgMn+5qaFYMpqx4F5oIaWvDB4twUEU7Vg3nmRe3e+3cmmek1DtZv3ubkdYtMULeiQ77bMwhU18L
KQscQad9aG141p0f19cHJKFs6l3VG1qjpkjuTBfpFFDA8J2Gp+6LUCCx/Z6xAGaoByDw1qho9jM4
adkDQHVKCgKJYu7KYBA7Xhwe1gCtzHicp5K9VnbigUYefumDRGPvDvNGn1RH/yd1N725iNBE/KHg
Cym5RIqrIC2CkxZloGORN3TqU1v55bemYBZ96Xa1+K55CBugkXd2Ybp7vYLmAAzDlQblwQNIe2Pb
iEfq1ZfK6AnedL1eXUK4FtOt0FJV35DnsbSPpL1xE7DqtOHLCYvt70nh/8JEeqS3OkErOXhQLuKz
GCya1vwY/l+u1OeIrZRyTX8vTE+ohfeiVlKZbDAU3SDNCGvhhMNECDCfXqfxDQq32WeO0JMea+6f
xHTFgIVNWMLAHAfZTlxyOPNLIXaw6005MOA0ODCsh3Qc8keSEUjNKaJCmjNtDCNOSlWH2Sm9VQzU
iXkBL5K1QXxRgcfPzWHpxOoqE66oGfk/nKswOhTczckrmYY/2JZ1fCbKEggR4zzwKlwC3x05Be1W
zTYbUgYyNm5tQe0pRqQZlcOPo6B3X6fHu34d2pfeUKgYMl6jAfhu402u0aiGtNzXI5iFQEjsJyOK
sdJseWxOk5EuR+5sERThTfIQJSiFwr87M90M6nYf+Xs2JMAbL2ig/lwT79d7wbcurTdJwKgNvSnp
O69dGngnT5HW1jgdvUrAzDfOpZGpBNnPDVsixU+zvz72yar9fs4l+J5hY/uHAq/dE6Tdn07uMEBM
AaeE+mfuPFL+DC9CI7N09WXYCPtctE2S3dGd4r3DG1PVKUgYTm6O/6a4YIgibtbpN4qdgA7VkX14
xuf9p5ZE8JJuMOd1hV1/cNwrcttKvaeu4vIh6gLwMOQ4hCk8DP+UgLiT2GCsX8NTb/38qmWzi66C
fstrnid1ui2RYGpU/FavjwTGC3U+OYaL6VhRmKJPK7Y/5pqK42jqqrlEC8L/bIEVL6d0kM6MboQ5
A6/jKIMwxpSpP+oA3cYXxUxNBKg6Rz05SurKF7fxFiLpOQD8ckKfzS6PzXezMBnxvqRGed2B1kRp
cp8YBsZFHzCxyqCQSNjw9WlPw9Lm9wkYE45A7vkBbyiNxQAgniMZ7ypXYLzI+iNVhSZ7r89XsKiV
/Dt0ePNR8qOPOHdOJEk3KsT7H0LhBIym8z1dl9F7AgI5tgQzhKRqNse1X4GDjpy93e8q4hHSw3z6
jmaoF7P7ZlzJGNumY2934uOPvkEAU+VZhI+fHsTMjW12+8Fk6ekqfiy59HUBzH/wwJ7/UZllxoIE
afqSLvBqODYhVfHiO37l8Mee2hCWEbkY3wxZzcPIqQB3l9E8kKpe7YJkzruXS1rRU+x4D3iKibki
jwcrtQqqfSJ21f8+9zQXvCVoyLguOwimjUL9czTrLpZOeOM5fpV/d7j9w7v5epFmhIsO3C6znm+y
G2Gj/9bcHBg17PP+/xWfqCFGhNYTgIsfQ/wNLtaB7tdRXOmmajrYEtcbfC6pL8UPFQWRg+dhKCIo
lkDvPiLhUPZAVFdVqoGBBj4BQUEPEeniNR8zts7bB2IiOUzpMvqFAJdt3UCrOg/qjvfwt4vpV8up
64uchZhefIAMkYH6naDIamJFotrJcf6W3NOKVMkcOgjVezsr8shUO1sNWK8F/0jRIacxdH3Pl+Jr
5/UfQuGcO6BzKPqAPTtGrf8Yxf5NdVretySugfB2Ny4q9/ln3Fbwg8Qnckl5MvGXVl2NOA9+urPw
qYoN3ZP8KdfY0pe3cd9cP1J9CTZFDvhQJzqpPVoWa+JoUh3n5QMyE/jYCwdg7pDoqwPXshZux2J1
tUdhJlgmmIajU2+WBD9dviu1oaHtUpAwzUdD6GPVwF7StAKTYx+e3ueqlxxXjiqh0rGEqJJf65fu
Y/lF5DM0Q1FqQ8gOpbL+ONicg3vhUQXLt83pc8wzmAHNjDR9eF0mueJ4ft0FnwKXaD6OggTFFhmb
xeJXkghxsJmfyYmiJCyGCgnDBMBvzkxhtBoEKtVOcp/8BNmmaN7nwV+nY1yzQMLvY5E60bRvFNnI
kDmB8GmIAALPTcLjjlKyBbtlDhq2zT8PGUGc4OJAGpEEqZ6PasbwUpF8JLWVQeho6hF767I0+VeM
1RpbBMq50YpOqZePQl9cCCqHIxDejuwsrgfMCW0rvFsjAKhkoSAg8grLVSg8Yc0/NWZUqCRTYuIO
GWcsSaHNENVkPvSRfZKjmgYgfaQ6wReoalO5xxKnLHMJy9yGFeptjM5ThyF6U7662f+vOmxK5i6V
KWidPEHkzt2+k0vY+D1saX8tP+AkIZImtCsa7wToNl9T0u5CpA3vsykr5cALXPFEs0OdKdT2qKzp
Kb9m3JjswnjWDD01eXyRI/LsgTrBrZFoqcE6LK7F2EJU2ZuRTmhgYn14RF79nap2YvyB1AsMAQWF
d2crMRaR5qghAgGqyDqCOS9qC/5z27soBr58AhEMz5rM77CLIVCEHJnAP4HlbUNXZWsL3vSjOAWv
vt/hvlL/b3BcgCH9WKkVRnppjjk4NxumVtpeEKGh1Yo+sFh1/Rh4zwK4SXYiokPL/zIgkmNFKlJc
M56q+odLNEncfrYjOmruRxmWvxKiWwnJ1zFJdqQqi3NEO7CZfUwWMKLU0Zzn3HTYi2T0VJUn5CfG
YtlFJ/QSroGaLbUV4q7tSSEHDcogfxs9RfmFTsIix3aCapJz4KZJ9WTQdbgBwSlaa4GlbLcZjRWr
Shmt3PyWyraTaVABJCTV2iwtN2UeBnaviqAco0tQSrqTw+dmm6K7C2+vYmzaQib7JK4md0k1ImP7
OG2kX6vj1n/HmHdCWOpDZedH9c8pT1r8KJkitMQqoz6zg/YMBdhvNqZ4av4WQjxaMETisYrjIcN4
sm2rDkfxSKd6hBvtHLixtmrcgKBzSyLM/FENAGttTk7sbkEzY9A5Bzue5MJjSsPkyAO75PnCM0Hd
kCDCkUNf5c2mck9wjx32a2Bu08FyOlWOQ3awRnTVih125ZvloOmsdEM2/SNY2Cuo7e/IpOmbcT9K
VB9bqqSoySi+1chjxZV2zR3EGeisGdcSBnx+eLG8RtY7Aqru4pQ5B8FHTDMC1t/ejkYWIBAlMXMg
j4nz5j/ggWATPWleBBpM1UII/vesRhOPlY/DcEGUHPzojHN3oaX1JEMtHuMXPs9rZFbIm8avJgpa
YcCl006ILrUkwBnqiDnTDbYA2igMZCY04Fr8zWKjGj1NQvD9XyF97cW3ir+fvGsdQszS1+G5U03b
h/ESDJtexuPqNBCxwHBOW2y1C6y/+03jG1K8C5ZIluL2DM2wncCT5yfJr6lakUHPrcH/M/paCmH6
h+fo4VuA/BFrpIJLQwOFMSSVqViU3ugB4vrSMlzOUT4wPYQM2gsChu69iyOU6NdikwPr6u8HXIB9
zf2FYJ5zfpSQjK3lx/jWzaeP2dTujCKqv88JJGCdwrqHmQWh5BNUgC8m7+jiL4ZuqJwFy/unIXeT
+NqixOmWzvv3ssYDEXYFH/BYlNx2PcuSR3TOd+vVFcjgGXNwT03UCPA0+5DwTZHByACq9XceTKcR
XxDq1ZPd5j1jjg8OGCRS+20rVIqTUuRXqtqwPjhwyKpQGOtZr8o0QJKSKB/WWb6qf+dHCM8+Jvg7
rfdIC83C6Ue7T33s+amaQ/L5lhCpL4Ca+LesmbXo0d9C5Qg0zW72HAwYvy2WrfBS3lqqure5BiLN
e8yAMsT2NWGULEQoT5dpl4siwZOUnhSYCaO0/mTlZU12lNGelY24cruqymSzxLYITCjBWQqsZdvu
qGUwLsUglYVIYqToBp8ptDn3CHc8sQB3L6nz6pEcsc6F26e+sDN47wloqMcZUsHQB08s+VsLuw8+
9blDfFgczbBqBlHrLzEvY2Zi9LOaxZ4afqiQh5Kv7aDJovyMhm9PBI6hI0cEnF5juZRY1XXmID6g
9U/P4CLlFATkPGDFSzM+Rqf9mkfCx2K0WhFUH6clCwpI3xsJpKdv8kuZrYvnjkZqYwrycxoJLxMx
XExpkU+tsOfhpfdQzmoiP/PRePUtX0ALMcQaq5QKqBje6TetRV4PdzaBgLItzRT+Y16mTesHtfmH
7G6YL60gkrZ2BDRGiZy+dqXyqqgwb36WGLSYKfoyYUgTVcQscNH/HmyF2dcnUsWYecKzs55xTnUe
ciKbdHLcFx/NQ7DeTHXBId4pcszFVOpVrjmftkfmNdqR1yMO86xSZq0YXLa+HkF1kknZjrXsLgwo
2a8B+lEjqmCQiHsENHy97c+dPWZbwl3e+G/J1Zavym2NiZFpbfY22ZtDvZyjYsY+l+al2LEc3MOi
5NPfh1P2OYbEhOJ2MHRH75KEOpKsPnhuJFkB0qk1U/TuxzaKFuSA689pzNpvZwP9FIMFoaF1VREP
iPz/If0lMZ6bGirtPUlqMinstI/yziYYsMhjgDFnoEPkfEKl/fSvnywEYP/TJaurh+q+6KuPkGzc
2itTIhAaiuU6o5+Ls3yxJfqz/gamZi9xr9dOP0xYr5vmppxrlu8bAxBR9dFcHsT0pRJy6XPE2F9T
KluunrUQin0aZdlyNGlXnHecVwy1dRH/ligNqEj18iWu/u4MsSZLJ1ld4Q6kgIfX3+LabTqz2KUo
MZhmllrGl43IgJj3XcR90R9WHDLCPGHL1pHRm3CkSPzgdgHNY47vjEh/tl0GJjV70pRpg9G7oYzV
7rAQcVwZT/sB7Yi+TQB8+eWKVwNbdwK4uHNS8m1g1pO949Rn29kmSwy83VC7OfF+y6dqvLyjSKzT
3SyRor6CIFFdqUrf+Va6XTR11/lz0QyxswVko9hZK/TSGc5T6Ypk7dP9lDlvcxxq8Ot55PPK0ZED
KgiLivHnbD/6luls+2DT8mdUp6G39PIu6XXRK3ZKVuyvEeZ0j98/Q+goCOwUVGg5PtBuJIyQjT6N
wwdoBj39GCJpQphSv1KPo+thm2bCtbOSoSrfpUb50DFPrNw0faVlwseHhsHeeuD7P8aiQFeItA7y
eJf5BDjL2wiMmJ5kUBUiKICQo20ZcnKI8J2PBpzLISXDHqiMezNE6MwK8HOB3uGPu/7HLMfyyYV7
pA3fux7ZInXlUB4KrGF6jlOENIR6cYOTzHVe4Cev4DrjMORia2hX3VnmwmcoYPc1wTgKzL+tqI1b
4rO41FAIBke4rkWb8SxtZcANzfQ7RPdKpNFyV/SX8d2ia2L6HIDJmGmjJaPUUHvnvSU90q9PifFo
JE7qXL24IMmIxfd+V1ojjz1JoRHEc3UCqw5GvI4Xn+0LSvS5YCa1WMzVGL/hB4gPn8YVIMPgALwo
TRfzgc6WKeNW2Q5Iz3ZcXa3WpnDieGGygU1QavG/rbmOXwX42Xa+lq6gYbCIimre98Wz4leEakB5
9SLCura4UJTlCeL4uZs5E8usLxQ6RgBy7U/fpNSKfAI2h4bZyQaOjkaec8wH9Pak4353gJ48it7B
VapCefTqJkxHt3XPgvjqjSZisRWbnBBl1+JO8DnXiRs/PSgPf80p++EAc93acz7pJHOW1NrYQbEX
dTlZLkBURmIveCuoik4ziHW71iGBdG5MfiXMx5rlDWNwaCQyETHqamaFdjbW67cF//rS4OZ6Oe57
t1aoD/TpDGe0AmN6mxeTsjPaVqguijkijjOECJUX4yYNg1PwH3a2bXk3HaqIcEO3FdWYuSMMiF6F
IY5NpzsSxdKF4irypNycX4v7oXtNoE0Ru/XtxJMUPArGyF0IohPW0g0NQtbCT3+F2JIizj8DRQm6
pHTv/TXSokZtEt3ZTAfCB3dKQvtnOTg/5MQxImBmljxpCeqHaiMEh90aLLqkJdxlagYFKGuEfDyb
1AIOKObPvwtfOr3eqrDciE5Mf0om467C/acN2WvjWVKJoZPl8wMv7En2BpP9gnC7b9YCDzdO7GIN
xkayg9tMVZrYuFlZOt24FFtqPcBDcDovP0rfYVkNlJDS1kjXJxj8ef9y5x9mi/3eBp+VMsmb/JD5
KxGBXSHwe1EIbXT8KcN+40kn/O45wv5uLmqeykFqle5eCNKQJADyEKJOIS2o0OT9eebRxuKLwqgv
RMX9lXe7va9hPEQN84hkk7TZ0bd5e7/kIYzou5qNAKDg+s/Ki3j0FiZcHwEljhP65PHomg+5ehE/
DHqerniDsEMDe6zm6o1r7TJlHpXgK76PdumGeThMBkmXYvyINSWfudlCh/+3RT0q1nmHJ31CK3lK
Gb0g6ohvhS0pXeBKtBPbZzlnvhTeiWh9QIsv7zoU1huyW3sKZ7zeKQR33XEVG5q38GX/n7Tx8mLZ
7ZvrfBqLCYSPb6B/AZmDjTgTqHWkogyJ5iz9EB9kHaBN4JFfFBz4TTf3n2vwjnihhSaViH2qAHpn
kH4X7a9DkJh1NhPKLJLXQRKEEr3UyiCOuQNVe56zw50WCsx2lo0ICDkuAXXeIE+fE05T4OYaIABG
Vm1uBqjQSHtnuIKRwv1P1aic8wmQyFeZJVtd071DNITJlCdFmXQntIUeQiDihnGTZjM70O4eD5/D
AxwXgGvnywjRXUk92aQGCNwP/zHOxExn9LJORH273TmqbLGyIkvXZYALjAiWuynLASzH7Ue2K+yF
TR+6HBdc3uHy0xcmVn95ADEgrYxTtcaohoQj5GaDWZBwzaisMpePlardmUIzPYDsASkzTmbP84U/
JFr61SlaxibN7R2ibZGqMwAMpBKcSP3TQ1Fr2WG4jHiAWKAKS7P2cCA/qV8cmQ3KP2EVagXgJ1m7
+hTJj6m8iINjlYNG11a7YCO0zroYEQNjMftUuQNmjwDS0NVrv1ZVt0LpBFZmj8lv5LQh9WFUOlOm
O7cNNjdbRbv+6RtnpUEMbWQmf2+cDtZLu4/7luNmNAdTu9RWgGXs0zUX9q9QpEk3LOFj5amOYupD
tK0TEcjaAezLGx7Zxc/ZorgfAIW7fQEVbfiYUlRcGftveFFCAv2500r28ZDOz983WosJinr9vWSw
jqbBCJeybJL3rNTeZMBbfxP+gDLDWGdALhDSd0Mi19wpPpDCdxCxeYdOybs1fUXTMLPELJDvJjpA
LXIQYFuNp0rLUmwIc66uDzbP9yCpz3A1+PfuqOxNxswFyEjjj8g/YbK/6jeFSrBuQ9/a45gl9Q8O
B1c5oQ/D7cTI9pz+YLVSzTms7gPhFXJ4GzPX4oAxSICzai7K69iyi+9HVvAZ1uXCzPBi4fVJ6PZs
uXDY+H3TtUBLnnQPnCLVoVT+X9tiOMfIGQHaP0gHzAv6RKnCVDKosqvbdR5Y0nujV5a8iSw083kB
OlBjZgJgsB1bbfra542RPc0uLXsYRdK0Yb14Wt77Ug0DKwj8AHJXumQQgHHPsF95jD8Jz/KaytBY
BR7Be+mftd/nwfSpO4JemrzI2aicD4kThWk1Fw0tYc77pxQFm6BtTFiq2S0ZJhH+USZ6D//kXnvx
GLUV2tol8ETwOIMQgxu2Tq1ZhR7vYdNc/mwRodYtgGJDtnPz2FoSCmeMddspveo412K4GE6nUvkO
HV/3VuUomXq7t3WtkA3X8In4TbcbyfQ+Z90ngkMhAb0NVGU+6Fhb+Pp2cRnN1rC9a20LWoGvXuS0
qYde3fF0WcyzN1aifu2WK4zDkfE6UT068Ebrv8oaWNdtcZs7B28Is6BKTeuujJd9w11WqBGy9eQw
Cqh8RdGMvaQvhOEzkgSpH9B0dPyN+PpJbpzC8kESdn/bkLXJS1JGWn+harBuFgehuSJQjoVG92KB
B1ZbTIDAwu9maUv+Hh/DlCN2i5y4rBloRclrD0YPg0HjJzNq7MHUQvq+2TgAinxkG/QqYDbRwJ6D
XEcTXGsOzOREEPDradZYMZ2eBzJC5Cjd+geDXt/Q1NAfr6a1EqAn2iYEAKixKZh5te18Vojf7huD
DXLGCZWUW1vsKIEa4Z0FmBATJvptcIDGoQy9myD41HN5ZlGfA0Oh2QI8+iegs3A/eHCpbCC8iLfF
S4gYRduJuYrBT/iGH74wt7Cj49+B6FnFrfF5es3RkKVh7K4+KQrnuprO5qs2wq45QnB/bUqt7fjD
7Fho3Oc/dsSul1U4m3nOKEvTAjOfFcAvynTI8Rkznq5YC1ouG9C/S1VBa3neBjWjiJqDSkLYg6da
+KlhyMnIFppEdLYQz4A7cUJ7S42Lkyl9ll8MS8f6+F2LFp0+AeZESA2SW9I3jGzfSwtNUMNc1zC9
RM0/k7aBncyXHWi/0D6kQhepRUzb469Ap1RDSxAwHDnASEJX+MvU3BNWyDs4mtT6aaF+0zWxEegV
SjTVLAv0RevIis4x+J4XPa4itb+golsOMike8ImIppOL50gFLBez2nMvb7SKdxJNzAwTV8j5iQwP
R5BUZ5b0ucEAV35veamUvE5tmrwR7hj81I3WYlgZENajXGAZHwMkuLGx+/y9clnQFZXK00kADo2E
+JovJTw2NLB/BYZ0uF3XhkHKMh0Gfqy0/LaPG0nN3zXMzak3DsGH9wSXlAYpO5ZnD4rt5vDcyQNd
Hc0EkgxiyXln1+v54xfN9j1HIbI11cWD+OI3Agayy1YMI7sTVP83VQkBlUfj9KmeGEjHQpkw9KpJ
ewYtm8nJoto8vQ0DQdDAQE+JHRyz7HWthC6Rivi6sfYUKppgC99gGlMGDdjgY5BALXgGqvTBb4+8
A31sEcjwjvmZMAC3W9CXrTdK4/EvrHE/CeLkuaxNQJhEF6xYPw0AWHK3vs+63NlvTp2nB6H8rEG8
9ad3XKqktPHRrSHc++lUIMvnMV0eKhbgaG2ElxMwPeBS24aPj4SP6kGp4ajubZMCYh5RoEOEBJmP
haLE1KTaHfJWxDv2585mseuRxeda3ehYk083tCu845DA7o+0jgBXwhgyK2OWsUwWbXt5gZejsh9/
7LhE1aNeYF4iMXlBEEhBnON0wgq/R9tj58brakMIs46jT2p2qY4eZMyT48vYx7p5IjMbHhWZnOLt
plwusNKzKYOge6N5PGTKSa6XUHJqQSwsR9dkNwxA159WMnD0v3G4/vSpbO51qJjqamgUYXqiBDvm
7Chk2hlUunQ0+Gu9zeV+KNStmhnRdzpXN5NJI8qcjcZA5hw9p92lsIEPhww6tprQf1pPjiwByftS
pXYn0bfuk2JZl6B/ym4iCf5cEu9LpoXgL6RadEX9LAA/opDQVnrP+b/1aa8lFzKIYAAZrQvKpojR
jsCbcnTaouvGClr9OtdqHGPGmloxNEvTsvYobCOeot0CKYEcqNBVIz6efg5k9zClOVCCcUSCwVeo
2j5MF3j/8E4wZIPmNGreGQhVHbmdEY5Krt1Aj6+Si/9l9+JWfjhkUg20DPErORBYE2k9Av1eXTwA
INZTJ7quxWFN1DI0qU0TcvbkynZeRKxwFP0LS91Db9xt/xLx0I8LD3LYS1UjYtDINhS8RLTh0/I0
Qn/KUUOfS7TgtgJbu0C2g/LaV+2Ken6OjvfhnCToEiZBtX1AAN9wkOCkK/zNipzpLn4JCk6B/QLl
DC19hUxUJPGsMWuBs290RL1kbysG123zpph1I648DXI5Lh0TYfbgGrYDC7PNYLnsyNafSfVC1uEd
cIEkQIBrNEuddxNRmNW1EIwEZaCtW6HjJ+LgBoBGbOB52W0ZJgFqQggOgTkrLJ0F5hPAKg+/RLCx
RFMXgfY8KACmYwagA3/PHnmvlHKW7Q5x+xr9v2JW//LhQ6VzH8SMbP3T2FF9FEqUi+5hhUWD0y2A
zQrgC9AjCFBYeYHioPw9JVlOmfuBGyr5X9qAVprEuAyD8KADT6CSs807mFEaYTEOQY7lresnNWLU
ATIULiUqu05d9fUFtHhSZHUb1D8zQFaV+MUgj+A8pKSyHruE2M+isSIrUQvbV1y81CfvIDvR+JOn
n0iFvGj5XkODCc2aAB4Ped7+DELLS8in2hU+8XTiFYc8k6N7wO/8o/9hK2+VgQBN9+rS6yD4/7kh
FmqbM86k3GxNQ/64F4gyhaA+cbozzMi+7sZXeBDfDuEgCNqj6Is7Rjhh2sNYB0XTbXBlI+lCfOoa
B5KIGErRbQCMb7mtSJgawoE6rB0Hy5Rb5syY7ZtGqUcstBVZrTYTkDqu3ahedBW+4737hYJGNDpI
3TLGZK49g8hPE6VpBOckqpLFMSrm+sJ8sZqM08r7937B/6+BsjeZmcIhgFsuXqhkBgmfeeceTXMn
ztDoyDfNUoPtAIlpRThrQvc048sQ+uMAXPts2GaF7ia/UvIymEt5QwmbfPmHWxepcuERu1WOOgyi
oELqjdhijy0yNwuaUvQfu3CMnvM9OFliF0eqZ+lFGnW1KCCr6tfod00Bioa37zOAirKENpGTGoam
UaECK+fwBHoPkYmVuh7ZwDlnWWnOMp8oeFwj+WxBRbQglhZNLqqCBa375ZzmxZm1OjTEo+9fqU8l
S4GKgCZnr7kGtiBpkZlFDHKZ8S6LDIQrcVKg6CBP7fiWPzd7DQS24H4rpeNshPF0kp14GN9FPKFx
u0EtQveIZ4I5TPnBdtsflQ9h4xP/vwbDt8lDk/dCdLLgxj5Dj/KMewBnZ5MRCtxdk4/yeNWVDKFc
++vGDbsjnbegGzillwmucSP4+rxutAn+Sg9XwjhVg5hIlD+kWrHsCRLkXQs/A5zWO/wKsNRB1gze
y0TQXSKQDGjPgZTALmvzf3clDXrS52Eoj/7pBYoQ7SKCiGqaDV46obj0KWlRPYFQ2JKlGL9FxUQC
OhbTSS5iPBYbDMuvuJ3KtObnQaua1yuj3A9z86TpcsEjOOaQrrhAOy2yEygVBPByvCS6x6C32qW+
RsAGp/5taxtP/dwyKIvKIFsw8V72A8xMV1lpqENBRjev6ysG8zu7zmitwN8xyxWDZ1nI4CJXPRnT
CoWves8w2/dJaStQCTCBuZECZsYeLoJx2NIV/jJ2RAKJezlSQjva00H7RNNqcL5FPhct3Cbku0HV
/uHAS01x5664r2DOn+EN52L/eZu8ltq2+H5vtW+kbBkRlZx0trubamwPB3QCoift7rW7Tftxrcin
2GHDABkQT0ZMjaAsd6Scb9h/oK+llmRPyhZoo+cEQJds3DHkHLyIA35L7CxMEnDtyOiQQiAlFLmO
h5v5t4Vrqvl1L+ipU978BB/8YSuAY68ZrnrGbsS72eH5rYNW/Z8r1j/ElYtyYtGTATQHvCQFNu9o
lqDLOf5WCriTVEQneAxrPoorp9DBE2Ud/T2WQaK7t//+L82aCthPh3jBcjP+wGW17WSkXwDF3A+b
Sw3mwW9e+Pe7C2AdTEyYyOqhn/X3UTWYi2e7bi/SSfY0XmDz3iiO8E6WD3J7SxvshMo8A+B/Axey
GDFx/CDr9zRuxJ/pgEc7i4EqkD1ehWZoZr81b0aV7lUhYmdJNnmpWEMqU+dcIhYldvAPBt7nt/Oj
c14cegxGRyErbEt/n7KCcxGiyoREeEdB8CbFH0l2kqliatYJ0GpnrD0bcmIBzLCoaeRypdFRwYOv
W3Z9ZL/N/cT5UFKc+oNRbsHM7op1W3qVMyb+4qmWYS8XC5VUOnxgU8X7s8LqPS3rWc7pSIvyKpi8
PyjJTpWaeuejWGmZPjqhPwTlgtr5Q+kN893XrwVT905vMuIXoofwf739lZH1/FzZxn16t6xXJDaw
39AJ5uxmN3PlT662z3KqjL7r9prFvbG5fvtBvyqg9OIMNspO63a/b9O6Teyq54Ujk4jhl0E2YaZM
IsALIvfZ8x/0YheOMMe4vitShiiQUBrmLdZGctMlEmEgLVyIb/lIu5a0yETMsTr/fv7JZraSK4tt
AwHSFJWqB0Fdd8RRRW5LFRdTLlL1z5H/SyHcsaCXXXFwBbAE7dF3qsY66GUrjXIFTi5bUyblX6bE
0I2it7LvJMCqxoEojKKK6KSV35VeS97AViDU3yBm3JbkM9I+EG2AcXbRIKkTMAfeXTSXKp62P6cY
qZ/Z0CmOOJ37u1t7nIqym18p657U6vHSDikTd53kNTOLSaW/jmYnCV1W/e/N+wb7x4enjALmxzrl
8SytA5XODRr4CAmLXwHr8x7KlCwoo5knTKKWEhqOVGAzGJgfedfHEojSIA2efeDyo6f4NbvxQEeI
ZxRdZ77Ohmq3hXCoW7LbJUV3juHFnT5eav5WDt7N1YErSSFA4u/Aaq/RxWIt1lplRVtfIiFvM/Sp
Cg0wxwNDCYjB+nT66TlfrhK5cHpkOLPBu+HHa0m17bxxn7n1qGtuKBiqvHDWbbN/pF6ly6x4LUzz
O8D3EZDNjeJL0qIhb/gGwRSksZJfPaAyfvLYsFmQgzeeWbZSgyCwge8SV06RbbbEvWiLKuaObhAU
7KRdFOAtgcoBCVqc6q4mC++UZiZ1BrBE4CA1BE/FEyaCA0vwSPPMazU9w0W0r2gtK/3jK9RNkyG6
akiH8G/if+WV55BzHCOHLtZuhodUmISpIw15smh+g/vdNSwfz317/9gf9b0dG1GDiqb8Gv/WdiH8
vH3e9AAaj0Kpim4UGTyg2dqWF9bvdGIVUGSki0oCTwZI8Uw9J4yCJcuXmdxEItuR/mXywG1GxGTA
U4Otfui34xZrhZ4vVR/SOoYDFN5A9uBe5rtmhJAsy5mFaoQy3LO1UnhjblEJ9RRxKPGYwFpYk1Be
7MRl8Ec4RMtgirlQG5h2tV+YuCX2La8fpL5lZAZeHyyGphnY+6u7Hb4zzPSoq2vNmMSdhxzwCrTT
1r7O+WVPs6fYdU/Fy2sIl0RWBNDW0wF9KVyZ5BcbfBxN/gEbHCScj1lcbXyJTQlrmYL3HSQ+0bfo
6JCY+4+Y/YCzW4f9mKLaaal6QR4icOS2AO+Uoz/UB93qbQYoQ1eDMH6s/cdeSqmpPYI6sOU3Qm2A
vNf4/5dCl/2GEEM29eieI6CUj4DjO+0a949/j+IRHgEN+O2rhRDc2Tkenbk0TjLI6HTnAm4pXdYI
0232hNEtiulO4ulACTOugBxW+wOtPzjRwX69jIRC/bc4VezEKHlbsfbMxi7Zoe57+Fe0pqNuZ77N
AYgD4zBpMuL+h29Xpnua1uFHHJmoi0yuPt64eDAH0QkCNgy5d5EDpTEjtW7xCaA1WocQP9V/o3rm
cnKceNg1OF9CoylP02FYThvI7q0Gd2wOngt203306O/q1c00wslHCa4ScE4MEaiWOfp+YdfSKw7Q
K6I1gKacXwklc7mAwgYqm03AFlpm2OHM9wRkLp3XHNFqei6YOV/76nyhyibWR63UDBRnVR9bVL6I
26Cw4p+t2tUiyjetd7QgbRogsAVh7tbzzh0X9Eiiy44o11hPk6T/xnbO1UWB31apU9qCmHhnbp4U
dUHX8s44TRl9hD/RAVXb6kMgS5hW3/sl1BcpcjbBrUzdF/GnDEA6aRiEiDTIJwp21K4tc16mDyGf
rcx+s/T4ZDtTfJQckeY3S1Gzdx7ZiygEHSh7E6oNmcjZ3SJR5Zb/lHhZza0O9CkFlr47d+mzGaSx
FaDPOjuGtRGoh4PkXC1PIWtZ0czxzZjMGrmbuHISujX8OemQWTrxePu2iKREEWecH2bD55X6t1pZ
cvOTr5k1wZgEdVGeU6qPD/QeTlBdJxILHkpsMMJveeOCkW31VMgwnRw8EFge9IUpMj/dvzse45QP
N5Zm/IPwUAdxRFfzI3mGVTeSSMvUiZptskeDSUeRql1h7oQERiX4YrXkj4obfk0udg2dKffrUN/z
AMnmTnBgThHMz7EShFki8XWstOyJ/CvZoky1ZPxWOSSA5jUgF2QQIZW8JUM5gsRAofP13glYIV52
QWuNUXxooJa+ARErbewy4oVD1yv1u7y9uPh8oMOQfwI2GBLdooLBE/iBinyz8uD9sH9wsEITOLbB
/9KOXhcewKmL22hETMlQbZyuVTfyQF9NZ3f2s6whZehrZigvcUPaVwdXURFHfz4uxofxdaSHAkai
BgQ1MhG/B8mPC5Ilyo4bUJpv9dV+rnoKkteQNEewAGYt4QggupL6A7btLj7mcvn8KE8jyKpjU2YX
q8ZFC+4VgvvXbw3qoqowLo+sdu+0Lat+K+krA8k8dqYIB4qF5qLAYhNNCwax2IwrYLnc9PO/f0Ul
kKSaQzZ/u4CLgXrjOytnMGz6hulVpvjH4OIWW3YIC7U7dNIUYeLgElUFi0dNgbaXwzTcIZWXLoWv
9mDyu08tgsgULcKpuzfzQOe9jzE48A4JULO0wV9+Yp3/52PVxI3mA9800bvUL3U5sfWY8VMlsroj
jZveUOxgmQWln2uFymlNj+obcBRZecfUXq8g6vQ9wYIU7cFqU/W3Kz+ltJoUtvnlB9Q17SZ613Cv
Y7SoEZ804nIshaIIlSrAYuUB14PbBvm9Qsgb4fRP3/gQ7JreUP6U9c0nyRXZct0ozeRrfa2FgcPX
9RRpzWVbFqndmoBOfP+ZPcSdn2elwuJmc9e2rSW4ufyRgVYpaqg5rR+nUdOYjWaa/VvUHsnkg3UD
+H6U/h0aymHZNBYCs3d2aLce4/Yn4ZOC9cwVzu7CMxH47s89ap/qiKg5+mqA/Jxm+6A700LcK4tY
Q1cscOjxuk+NvxraJXpi/fJ41Q/K6SEETzC242n2+4X6edguDLnapv4GvCYPEyr5dldDC9tiQJzO
iDrEbYPGVQGTbvHj1T3NDJsBjWiD7gERAJzjrW+exQwT7Vjb076pxyKGZ7D3cxwNx23T1sLCHLZM
XmVPqbQMeDAonyU8LWTXBXl+CQZKg+/YEtDv4QWF+rp3OuSIE8X5WgCc70jY8jxc9s/ugzBZYLGi
d7P5PkPf9QgiWQ8WcYn4hoUaaT1uwdGLvQnOhWG+k7GC0MmpZivwTjRxpcJPbD/WAxEsSc+bxibP
5/c4gi8r2bvsLELtdHzKP6rWioqT1nEgTGosiB9zDmH4Ept2aovhIIqChsIdjA/tYT0m+LssHpLh
kffUyJVOEVoPfEi7QavV8fnS5BiQxXz+Sz1CyeDfiQ8J5HBKGDtBZKqJjkJEVyyzyAAoFm1cI64G
yLlacTmG1YxDyZ7fvMEYJp6+ISiKwcnyfctY8vXOsEqsbz6XSP3ZI+C9d/T2a+EWQtNgmXyQewoZ
fupUpxdMEDSmea/PwCZkBOeUIdo8l1nP7JXIY8fiqAPXX5Ar7P0ePCI2cdI88dvE8SZCCAoM8QAt
RkiP7y02qlH8Lj0AeZm0esgYkWVqlo/JLmtYmmQjkm9iM89/T62YmfHwlRvocopIz8iZQlD5iBjk
jrFoBl6s67agVRCfJotthbcymHLqy5Y7Gf+DtxbZIFzmZP/vMxu/oiMVYFe9ndf2IswKukCpjUEk
tTlEwc3Tu3ShBaETNON3zpOPBobfZ12av1oAPkxDivs+llZs0N1FLLnIbH4RvkG4NR82QXeoASC9
EsxGQti/DnrRLJ8TdF71xHli5Qe3LlXQQrgBUV2zdn6hcgUlUy9owU1lQds21bZL5kKXUrnzIjqf
1lkcVGRm0SMcW+6JJzoqS+hQjCq3+jYjdodVplQ0hT8ruOgiflrtPpSa7kXsnWk8HYVZFTRkPoQj
HHYaTbi5LPhUKdQnTPLhs9aHB5/iE5p9LwzUfiWzBDf1cRasq4anpKbfgareMTDg0wlF9ZG0/Gij
jPEGICP0Lai8zP5OGpzs5HVGP3R1JMmlyiY3YiN3Xx6TT68v4xwaeGrDdPfOIlDFit4ntSBiIjrf
EiB+QpRnS1qlaDcDHPAG6jLqWfe755sConudQQcV5mUftufaegruKbv4HXF4SSQzbCOTz9jsc2op
wPAlol4EpYLf+1tlwufKtMSGtvJVMl6o05chwEpXIqbvWfNf1VdNBjW+hCeAwJOl9i97nTBhR4g2
1Wdp4pQ8ZrzWBmcBPhrCsIoQqRQmiTf9nyf2N7ZUM6KUmyfVLxrNAl9ge7PklKBcY3yVjJ2yvTSZ
qFj9c3aEHpGsuAwgp7v7Lg3zY81r0BlM3jFOOfqwl+A31eixqcfTE1wJWBvUFnoLpGRQBCUP2DzI
SwH9m6wMrgYiSop3yCWzRjkPtr6X//I+yhiDvwoZEaAeevLrpDXvEaM7qaM6/Odl9rOdpUQD5bBk
Apveo3Lxg3Op/W3o7Ygwhjx5ppTmN/L+4dG/2gON8fUsCqy/CTxi4gSPBaXVMd0Ek6BrrKuLgNOm
2IBBsEugZRm8JTlpKqKbDNgliAa7+qN2zxo2kyZodk2CClbjIRyXY/wh3fXIb+9QD1ZVuIDPj315
Ci5OvhTobIvU3YrXUeo0WeLQgyY2Qu+Nx0U2u/9AYAfYBdckvk+loHdbKj6Iw1aiVEsGRp/51LDc
nm1zTz82TNJEvOVcQk9v7N2wQrIdJHbmNkn7TZysmSxuN4glULsDWE6Mm+im77m+9COrKgYVQgaU
boRXC2vNBfs1vz8dq8CF1Dcj7SEXtCesNJhrI76Zah9EmST+rWZTLUn7MHxEvExXbS85G2XXcNSm
KXEuWAtQ7LLkFTQvr+QBkcCvEi4QMpEuuhUpuynU59GZhk3TEQRRXPb+rQ9nReeNpK/FAfeCb7zD
+8Hy1FdLq4ebIt+O2G90nvLqHwpyqIeqCW3++lDgqekuilyBMAhf2aQw3a9JO2hogH8KUHNLmxuZ
8tqMv9RRtNNup1rdHgXM5B83+PYFwu0hQb399y0iIORgAyxvgGcSqU/Wm4YvYtiq16bFr6tEo+9l
T0G1xaCbAh593j0hRraxz9CQM2niKQUt+yjah9F4m2zniLkijOHgRul229gM5LBnBxO62c0y2/od
Ln6qGc2PlPs4JL1ToWRF5yOhh+nLDwqOxd6apYgoyARuIRcmneI7ROtOTxbUo+qb/Np7tGsBgBDT
DNybOVJqUMfzpZ+kDR6lZRzcDkCjHZhyireUy6J0s5YIpPndv8NWBdBt5nd1w4TXMTRdYKGxrEyY
eZ5NNZRjBjrw/ylaak2EWMgJ90avzC6aMcdfFaAOJ+IPkTHEtr9pHl1TjnuEo7pKriymZkI5CibZ
OSJ1VmPeVtHPqCtFDpRIutEcllstg21nkxBw8IuGcJOC/UF7KXda2KLcLyLNHgxQWMszSmEE8bf5
fSz3B1yDs3J4W7mF04hdPw8Azi0FyUjEm7DAVjSW9DgY/Vrb1KG2Z/cUEzstElLXuBzO5FMYRXNY
v3tnbmSrltSwIOT6y3UQm68+jhc85gJYt6HkihYU1wVvI4RxKRmX9WfJezCucmaQOzQcFPoe1aNG
M+QbMjkCSLHxaz1uREznSgnEE/Vr2gNUUnGE36BWs19gSiVYMKyNh9JOzzK5CtjWnruU85HQio+v
sobEsQfD1DFXw+z/aJFowSlFLBZJbVusvToRIIsKeMV89NNBt0iStq87xUBg7KmOwBbCUNEbucSO
Fmb05thYLn4OSbp5DD5853mTk5wgdG/umX95PT2B/xRHKiurJMNuf3AfJ8M30nxoZ9jqpyKCj73S
Z1wHw9kWc2OTgMEoFB8xk/rEYqTQHWKr/G24N937HLD1Emq6SUlF8dBWkY4k3g3N6dSFGM+zq82M
eQr3Kxi/fnn0XBTOkaMLbwPFmPMF9TLcn7nR+n4XC6yqoNaRb1dEq5rbXEecEG0oELo62MeCAFhf
iCDj7Q1O7/E7t62BpvkBD4EKTO+593WbfC5yOi/K503a8EF2FtdTXkeuTsV+ceJsIdHOIFISJgy4
h/HmsExRLBSw/Ui/Zvdz14+CjjYEiSePVtKlsOxRJ5JJ/CivfF+p+BI3r/LPrEtcvU3SSMpN0qMG
C3OXbgO9LUQ99SHXlEsx6dxoJWtzrqpbyCYwiRTfUgR2/4h+JAN5fwFHcApqrTP7Mj+8sJtIf/CK
4DBtoNsQudo/geeAJ1XNYYgw+fBrCCjkkhDSnLXjoUmfsy+1i4GuAlFOthmtc/9AvWCABJWaJBP/
rItEs+281CkppIS7vQNhJWoDVR4VJlF8xZHiusB5CzWl6901IR63PR/X4l8wc0z/RG6nkRn8X82Y
aWtEJrkzAWXgGtBSAPBdQ0wkWB5TSJwJldHpSs9XXUvB0JeVH5mIXQ49ev5qUwBTnj4YoiVbVoCe
3TR/suFPA8sI8ieMFyqz9PDrV+Foe8eNrg01CQfJyJnXwX7l0NnXSLPUSkG9fM9+HpHtXObWf5vD
DjLEnbPhlSMNuh9eZQoR1BxLXSn56z58JYczD5Pjk/vTaxuNwmN0RUqyo7NCrJtwF/69aNNuIk3J
HG1CE6XmmJOG8U05ouV4hf3lS+0wk26FS1IkMfoWD3CDlasRCDHdPl0TBOxpDBxgKo8t8HpJq4I0
EM7PLOAKeQhnoLb+gU8k3sl7Fug/A5rMhaVyo6ST/KXStmlgwjsB8uywZI54clRnfV/OfwmUVDyW
6ZJsMkcwfePa45ZVmG/4Nl7lzyo6ISRem/erjepI9mG+9xyTEcxszNyUr/0vU0UjHwxye2DOriGk
EmvJZsvnbUnHQpR2TrnkfnBCSlToxvlKSawKAWIjLi/jlEG4fnYkXYbI+XvBEs7ePf0nDiwZZQKm
400oUzVcXTR0rPLInroY+mcpItqQI6qo7dLr2/dLDbLtdRNXcwUdbH+3ONGhCoSYL4BE2PqBjZe2
54Jcdu385ROwHSiI8FSwNoqzi8+KBCjzeJAICvBUHg7dq8o1jIqWsAduZ9Nc8TzpQGztSLMkhFkD
TWCZ3Gds9JQZPXbuwgfG/9zBeTQnqULhTxj2MLVOY+Ne1LWeacRLVUHtyZhLskbof9IsEWpOhYW/
AjnGg6SWFlcVResGQtrw6FyObD5vMZYskv5pd8v+Hy4VeylJHoMs9c1hxJPg9vbRBHiXdnLEcFfe
0YX3YhqjPWoJU+Hf+DiUo6lqcbyp5+JJ4mF+WKWzEsY51zvw5Sf7KCZzOwFfwA1Pb7NOi+5Wegx/
d4WIzZn8czkI39BXrTvS1bUBdpNEVm6vLC6V//zYuDf8vP1BceKHbYzAbWyLGMyL1uSviYcWc5p1
lRT0gUJOe6m1Pae28bRtOwl6T4STCI8Ao5mxYtRj4O/MfmvN6BCVJT6LxeoP0tS2dn5JLSXg3ghN
M5klfJu6hq1MZhkqz44y6q1cJdX/rpyfY6UAT5OyE/ofK+ZFNZaNVqKuPyi72ZIJqiCpzorJ2hk9
/dfID2SiwjZ3/+Esb3UTPyfEDMYw91GuYU1m2TW6q55awF2gA6vU5OFtxLkvQBEZADQE6GjijHHm
uWEEwYtYpj3RjEdXHaaRmHfm2RCtCQv3eHo6VGL5GjvC1SxYAwg1/1pqV5gSFgbW7/xBdmofAFsX
WdUrHNm0l95ejoNMXDfp4eTLxlU7IAU7DgC/DYkSmPnmDckN+prKUPFVT+9jXvFzbFwsDT9iddwu
ytFcUnhtk+Mx4UV3CTTaQRKBnNLKovS1Dq033iLUYFYVlBnAFpUxtqSroyoKHQiph87ZHSGuU7Jg
h19wliY+3rILDlYD7lcd53JWWLMhHuTjSG8DL7C6qUdkQC80G++zetcfOCbw8u9UzCeQt8NEvtXT
m6spcyG8vKZ+8moRmq2d+oBrmd3qvOk1A7L955V4NqEpaEiKi6EZlrLck8Fbaf7ZpPPOp2/459sj
LYz53VSO6mKz96xWAv/alh8r/eQeWzlQcXgX1gpMoyhq4gGk6ai7QJvhyQ/LInfOQYy9zStP2jPH
1JA7ca8a4fCoa5cEesIq09mVbJxfUCw5EWi6XCOHY/avUuveWzes7Xj9uC90M/BXS+/u6BP2MB7x
HhQemaF9zwHwSnIhx4DjqFvEepSc6L1qrCAwPbRWcl+dAuQuIUEE+D2bTPZGAGdNoX9Vr0yHagPi
eakRVQLZmYnhan9QVK6Na99h2SE7FsJxzal0WmaA0f202tn6iblqkiZSfWnoMqwKe+Y4Keowji+e
DjduYJm4s2lM+rNLVt0t+Kc+NwAtw7YdWY6Y1L7Dae0EfcoYcI8ADVsOMq7Fyne3r2W8LfoDc1ls
epgJ406IT/VbfRWOR///UfZZ67AeUvx7Mkcn82zWIfk9P+tcKq+/yDk4j5imqFFAQ4Uiin7e/B2Q
9v2uj1w3gfFee2ScBxX2jmntagwlMUoTUhJ9pl/cLY0/dYDGMlMk4JPE96ch7UAn/gRMc4+wG5XJ
80pT7qzJsxfn+jmX8r5g6xLY4O3fgOhcQRIM5cZ7gg/F9dwO5o0xrBRe9Qdj+tWdy0F2XJNpdB+Z
763trR0dhp0IP+60X2dJz/lRWXhcOWvTCdCcRPgggCEBWHtuJSTmjB1zLczYf52L6yhYoYQTqFgi
+5t4MzmNe4EzTzrICbbm12TemVnHl1ePjYmg1IW4d+5WDDLC9qzH/kGp6xz9mJSE2bHakEGZgp9i
dAykMpVGqFL9kaxhZa6VfE1IeEJ6VwkA5Bz97UxhIme/F5RDZslWblFXkWkSvJno1+rMWvtU7GCI
kUSg1OJU/j05x8DmePjGwopbmrfobWIkEUNp1lX9iIUcRiWHb8u9/v715IP2K902pbd7KwBXpASP
XB3/TlNxl2wQ53V8NFy6k/V4hOfTGIauC6uAKOZvP8W9UxkbaZ7tt6o3z7sT68h2a22eEsF44/He
ClrkUPr+DC91I7xfg7zSZ6M+4eL5JJjHe6GKQqu8vIIe9FxUn4liy+t2PNDXoUvU2egK3MvW6RaW
tfN05gZLvNCceKMUJlsR63PBNW0pYIYXjkWt1xDdSsexs+RSUupQrqNmwXaUOZ9uYjgHL4j3nLnI
aK5hVHB83f512kul0Dx+q8MKPPjW37WNG7kc8Ffuv1PLZKdK4U51xpEid4tQAYWKhLsL3bzya7Q0
dBkRW/OUmwKlc254GB+jJLlfOQ76HaFc5s0X63EiW4kxxTeNrFtZ+2APD/b69LKxOuu97bUAXCbd
XReOvnQMczWVoAnTzwbuVkP7OiFILIeHew9JyaGCK9kE3uBbHCIQntFKi458przNWjDRgwPNwPL0
I07y3PMpmsjBg16nCcYb7zbT7WeEKhcnuD3kMLnXow58R4eiqHiJNiz2a8qD9/7oaIBRsfSSh3oJ
ILswPSrdh5KTTgsjc8uYUhXzERd15+vmtplSlgX5SCRKmC7P27Eh6pQtixyZNbiWNrMC3HTYmCVi
WDy4ViPeHZxFvglF3KVnKMXyl1JkuVzgF8Fk68nt99txPpTRiKQXDGQ8xNIpyQE8a2XlO4NWZeDX
u1tJY5CNI/8OMLgiTMu2lc2pH+tdVFmocgQL5lvC1ZFz0uZC7EoE63KbttWnbR/Usjj39sPD3EqO
fkXIdoofLW0pHrSQj26zNdAYR8R5jQkT9rHTuoDUkOiV9YKD6I3c4GzUl+iyx+/9NXcRWOlvvggU
U5yGu8w2kPevi7IkFufMifWeR5Dys56HoygxzEH8BieQDR4oAo3GgM+Ui7/D/GFVOnGoyXmoQjIQ
EyyTXUWIqsfpEO4t8cq7fjhdqOOA8ov+g0+T2XOhFXn4SkEXr5Q4d+SoX7PUZnL8fajlqyhALH4N
d4JwCNsRMJxF4pYBcJ0RsufnANoPbq/ijHocqQxD9QmiIY8BKYLG9/J9NS+IMs7tyT2WbO5Y4y6I
xzE1rdOAaX+1K7x43QcR99EG7BuC9sgC+3JXlaOMPKn0NsS/lUrXjPkQGc4wGY6apNXBXPyUpElL
wuQ6a04BV3YJr9m5Q2PfBQBTmoPDjsuv3f1mIia3QrpT9JyLHEJZVcwT3X5S1qp5G+FILIAiiQaK
DhpURVWdzty3Y/jprLOeXpUsyDIuSIZhzJSHIdMzZQqclSZG4JnkC1/LODQ5dJna+iCq7BBEt4mA
HOcSgbCLClmoFf5OQlhaCw4GN9vZPlnK5rgUp2sps8JrmOUEJYze+rQTxu43zpjvaeFvcooK2J9C
vGdk6C9yWVKgear+Kb9lTetbiS4+B43QY5R8LfVJRB/slhV8hzq5LjTf09/ePoP8zR+T9yozC7A7
0mqCeUG6Fsk69Ix5L/F5NjR8ZybxTHtbPzj+A7lqQfoxDLcO0uN81RDTCz0bw0dROfGRgF/cuYGi
sZonxs7oMo/VwiO+ZthQy9ibHYlbm9VzLQBjZA+33ZE27Z0xJhHuK55Zn187Ft7lpqVRkXBCyV83
+jjLMCx6MIFkXEXCko3OsyRrfJnacUjZ7a6FnxAuRLUZUMJ71sDIYa+1ClR9q0QQP9xI0hXltNCM
lmBjZWTX00qd1DCtDm1o0X927LW4Y7xP/+paMZUBPdrPfraYM99j8+/n549pjmrSVr7SybfgtbTc
jdA9BDqwZYrSHnICpJvRL98BjOJ1U0TWskIPzyCcjDAbhnKiDW5B8+a1M9TQPTGP5lGPCR+/rx/9
GT+rogqazVlmnAb3qWHLUpftXR9/6KH/1uPBibWLUeBVBu8CZd/pmpeHYIVJvOUrq49y9iDpsYQo
D/MXA5xuxnXG01eEMIssOIN2Geka48EjidXyxlX/mdAPckFUbkaV7AtUZszMBVVbOvA6OuyZzi6p
y9BJviaZFrzchqV1ZUTBmauPDkAZzPO7y6hyta04hlQMWO86gfCLJvEw3dtlXlmYan5LbWtXx3tQ
Cb6TlOGI3YyJW0pwWl9wZ8ghZKGQrZS4pKnvZ423ZipCwzyXcTT3Yj9JPV1+9Y+eJ6H/BpTeOIhB
BYoKk/314nCh3BItUq0549ocYZJIJw4FIz0oXBM2ziDkdSrFO45A+Ane/ySu1/ii9Cb0EQIj6sY6
OPAOCmGrAQZ98ESyXSo2zeQxkTiodIVEG415SKqfva5VhkvC82WOmW6LmqGhnz+rHTEay5H+TxgD
SuEFlX4mFkAJA1k9zHTfNKpdmdDpWmlPWvp4cE2iDOfGBB5sNnfa5A63R2hRmwXpDn2gQ0STA0du
pAvrvpg0bKGNIAKukRilVgYPCU7+ACFlKlilc7VWyuzSwQO6Q2qaqDGJzNk4qODVi0PNWRkyU+Zy
lQJUxwp5588bmfWEBmxpqXJrbLjAmApW+i1CUoZTu3cy4/vx69OzIfW7qp6Q1tvdqeWGtqcpl4gJ
8BoBLqazqjQ8/jJ3oayVPZOX0neGXXwHm+yLgfLJ+Ccix/GwAR1KoUMi0++cboLcd6TyMEXnTDtl
1cVPrmZIvypz7cfBMatDkGbEL8ON3T6gR78DLfDA7rmcp+BX2e7VXM1RHDexeiF4SyAFXP84ZhU1
GcPVE7W2ENWeCJa0JhdRG5eNCWimfpipg6KnkjfUt1Iz41J80pdeWCtQ9sPI34GXuhQDR+a4yRi4
mG15Ch27/h6iyGK9dUgIYhRdQ8nKLy3eghUrhThe/dZ4KqfgSLlRCSMhMT2/6VtOjo96+OU15YNz
Lany5cR/wdLJKI3shW+nj9M9zpxzxCg6NvU/DBLWWZxCdwUi/eQ0bqC0kmsmB5KD8ellNe4rgG40
leceWYk9EiIdkfD7dL558ZVV12AyK7nshJ72t2mHf4DgN6s5GRqgQ9a5kbCy7QMYIp1i9+Dst6cX
dPhkRGz3qfqmxD+sFxFb+cDgPmzVVChcmt7B1Sx4wLzj8QF8mot3ttXuB45YqU3hfSnhkCfgFDdT
axpWcJx1ySSw9XpXzbSowsrrHFMsuX4Nr9VlnhzcKb0DVipSryNwH4UJiKzIR3WEz9eQtZgsumcO
1tiDQ8ynPtFPPGTC562PuqAC+DtH34vfN68VirrLo9Mf4FS6zmMkFI49mRn/uDlKNQUJWps25HFW
+2+CLdJ49/Th8F1oV4p/MxdZ8c/q8cNhqoafg+cJ8ur/Na9subluW8A7K46h0RGhEg9CvpVpsFMB
bpPFT8CgoQi4oVo+0XxgdGxBJaodFR7Y/s+7TgVHK7D0nGnE2K/WiJ4XO1aoJ12ZPbDxY6yfSwMA
3a/lK0tuihGSPuJoFNZykMKKJLy9lnHgIQ5IG02dtEgr3ltSFhsS6uouMDwgGSjeRGr/DrEa6e8t
IeAdmI0QRXTIFmHcawP5Y18mPq90bsat9Akchp168RYdlQZiugKcTuNRzmras3LypuLH4Ds1eoP+
kHUvDxrIXNgNmHYJPrr6rOhZJhuHE6b73RCc9LY2tZTLHRD+GnrfcOvq+up45+NfiNE5QHzslqCp
ZgqEQJgz33qviqmSXWwJnywMcXh9/fCbbhL4lq5pV8ksfvX+Wvul32WvYa3EIA7y0Oq/fQ+tsTXv
gaWgn9VIgrBSiZ5F6Qdwu9gBbL9c/V54OtQtToRuQdD72Mukz91VANWFHSpAOaQ1p1OQKq/hsv+s
b4kQvI/n3dymRjD5015bpYTNvE8PCjOcEjBTC2cdsr8aLLmvdJhVgKrhvJyOhJDJbaiDHmBhVipb
ku5A1/ubcDPLDqubt0tX5HSgjSEXxb/+PkY5vf19+5OjiU3SegpwLF+oQupSenzp4wOaTmq0BGvs
1qPP4O+QabHPJyiQ3RimsuAB454ullZ00u1pWl/HXGopQBoA1XY063UTuhG/l+rbxE0oWF9TVQ6O
EZMzHYOTdiSWUYSL6Mee4ZRLS9MUqdRRyViSWwtIj5TF6G9+EYmnVubTwkO9/cVFDyL55XFrNR9v
XiFv10n4+OduXjKp4lIs1KJtywkchf0fts8dxdDnj0YiOfMa8myiC+jcaMMi3xBZibxVVSMk1Ukh
H7uggH0ydA+IwEy217FQHOYOjQuMPTmkVKF7hpUpvlteuwdCvv5JV1R40BzGB01rEVbt/B4ntvW/
L8+c4is/7n9UWSPw2NefA96uIrNlnWeXRfbmekMuk667UEooVTUf7CGRdiiy4sjcsAqMNdDAKxsT
Gw4ryotqj7A5DFOrr+aSAUy0CQZtDXBH8li2cl8+UoJHHPHZvzuBBSGcyghlxElXgzTT38yileNY
i0qNU1CmAQf5PLqKtUIMKzVzi/J7noeKUVuntioQ6jC8xNVFS2h3FyALWZTMXz0a7UJCgBRKHm4B
4sWYJDYg2dn2t3SuxVL9KCCxLj6jtbnxszo1oKnvEWyqp7fncn6R89+ybGAs6znzvU/6JQmK43r/
+CF8jE9jYIBv870pcLVoQ8AbCI7/DMx56uOITn/179vUrM72WUtVia09uheLWqfasMSOfJjnbRi5
OZUY0/NKrSkgJFdyxWJm0jtggHJnkfYu11Ed/b3TQZjIganrxPgQn15WA+225h8lagu4l7Y6zXiQ
7WVv4qAm0v50rDUBrNYEY6FWxIDvreX8qfDvlpXLdgrwB6tYo2RqKpO+RaOKAAW1VIzMR5S4hlYi
FdPnmt1z8BHIV1NN+uEG1M9rNneDb7ciD/vIV3MtRvjQIFaR2CvMwZocHCw/Ddy/q8tW3J3zeYlY
w4PzyjtaonHX86hEqgSHd+P0O7VncmzpuPe1bcnaiRkPvJsqib3+4uj5rACMLzjoBo8MwmT7g5fJ
pbmtWqvbxFx4plDkyp2kx4WALyGrFIAKLVlDHTxTe+El7ivRCqeakn3MAGLGnzYXldqzXS1mS5+D
Ro6KyAQHE8pVjGVxTPIPofxeLvAs258sxs/Qgq0drbGr/GeYfrXiefKEAm1cy9jBP4KChWKs/4qF
aSBehSpbR+t2LZY9WjSDp6jjsjEKLo5+IpMz2Lzc1gTyajZB+4KfJR/abypKwa3AAy98oKM8cQOc
tfpvnQHN6xcMiRjDdIEMc+sDG5Gnhi5H/vBgugJmuXsi1qT+1X0p/6PhPBLa6LlyFrwBd3isHoDP
LIw0NrtDcAkBqd8MAE2/MxzcD+CnSqL4dapWzVBSco5524s0TLVovPU6GN1B0vzOc0OHVfM2Ksiz
6te1Vks5HMmQo4g+rqK1uoOOOOJ+Kdni4zptMtLzBBr+7r7A8XARpVe21zVjcR1qU8BuRqCcTYco
zqfNFQChCqG3a/fNKzN3EKO3IYPHtpcmgM5N3z4SrOS20totbNDuHEHhPS5gJdJIVgbVj73Qkp97
zoL6qUX+fZWYTsnqZRnfR6uxz6RjJKcNDUtGIjhuaEraXvv/YWqD6M8aF3lZvv30wKX9RwlPlK7f
1MZ6h3+yTI15uv1q5/2HuNh93DJQQ/KfFIs8pKhBA3w4rgdtNsffqr5JUtVuty0FizSVpf/K0S0H
3Uk4hFxL/c7t8FLcNCzeSCJQFSS5rpLFHwwGX9EZ2axA8gjV0aqMMw0hi2dJm47IIo0fIJtxsrAu
i/UHYdQYXE0TWu9oUVqhMlFDb1iXQRK1NdHKuYHC77QHeRlhuCAYZDwonI97LJgJ9KgOqZJUpH0i
sCA/Su69IMOcQDSCOkL4hY/oTYPhS2u7YNVmL9me9gqmkFcCwZPKrkrEroZVOr5vZNMhwh9pYf2r
8shP+3b/H9SqBth8i3WbfJIWggvlF/fRxuTpxnrhPfoV6P92DznO89q/c5jhfgDALXyS6+9aLYag
BuRrUxOjnbZN6RtK0T5JXjEvdJcKp5RAqqxSn/l2TGxUeVtAfLhBENBjKE8Bw7tNJvHLikDoUHdR
53cKu+9lJtVLoiNK8s7GB6AdKvvU8k3Z4VzsCdwRTQsIKpOmHt55ifI9HXaeqOwLElh6Fqib4rew
YPWobF2neZvAuxKgeuLP0CQKo5f3Y2a1P9yxsacJ5avPGuUCi6Q7YUBSCNB/CPfQsrbSlpqJqcHJ
Y7w0idssZaBhuaej/6Cpx2w29YGuErJAF+qx7G4wFA0cF9y1mSC5j8aQsU+wR+HyhX+Pb9EkblFB
8cREMesaUqFjZ3P03Ouk1IJhueYTQymXRuzj7Qg8H5qfELEkApeoyHrWiGKvmNA/tc6D+cIvCdnS
LvYA9maJBsL5jjQQ80QNBkntjjSn4jvUhmmh53NqZ0PSgI4Q92/rtMBQb+UhbBS/RV4SKM4kY1XE
bkJY0ZR0IaqK9i8Qtn2QBP/IlHLMq04vToYzpBfotntVLvWdyQQh/A7WNuxNLXQXFw4vKnVgSOTC
rGgNr8cFkfHgpF2SAFHjvTxdHKzKEuSk4nE6NaZpCKFBTjMd/2hG2RBXNEjKefrVHI3KvM6M/9rM
yuqA8D2dkzyi7wkZpXu11/DT6O750V3wEPnQwRckatZFyU/1SfsUg6A2Jx+OwG0cBnzE5hyH8Fhl
vtYKx6W/OEEjRtbCP+q8UoElXnVE4PZLBiz7HJPxtcq4URHYm19NwCT/h7031YSOG1IpuPPKTwbx
jipa2l/giFYGbkn+TW1NkDvaRttOdQ2PV6v9+KmARAleHFgUYg9ru5/ABjRHznSoFaegJ4kqPqv3
AjFsHlX7cemidrWnJQdq/nj3vwoTrgpbs9f7/9llTkYtEVEXz68d/0/CKiTI4SduGg2D2+1XhlOP
+NodaGUg/LNF7+508PcAgSGKX/17I8Yaf7Z5jJuTmKbasW8KCVBLu8QZcym0itRF3HSAwUsA5Uj9
vX/8OIQ6ZcxEx7IQGqzFD2bxhhBu2j9jfEWo64aeqBWFolCFna3LJyUXrBZEBLXm+5dppJdoMdsD
s/FdZTURzJOt9y0RQ31hEkfNedvAy33WjnpuD1toJx4QxSv75M3oGhjbJ+dwCpecIYlsDGuMpZF0
GPjrAOk3Ng49OEgb2UQKBuBLNpzEepzmQXeo9I4wpK+oKVKu+7d6j1s6s7Jx0X3tEG8oasbEJ2yZ
N5vhOGvRjkHTH+seSLnwUSN/1kJvlEVzr6/tKhK2IkIo1EBYpPrJZ8pxdqHiKG70lECZn4N3seY6
YhBleCzuZhZNVpJCoMe01+lwsmD5f3B8v35M9cpL6C0u4Sacc+BzPGdK406JBQu9aexTUX6L8BE0
MbNi/ERrYOgCxBl7QDIo8G84vsJimVXXw7feu9PYEXPMWrKOUj31VxUBv2pXrgk8yV1BQCFr0MbT
gNjiJ1FqKcEGfaq6AGQm64S/LoNBNP++9iYPoaUzM+13AU0ECeCvZskE6xRKEqgv3WuCw3rd7KVr
z6YLpmqQk9DJxoj4+6ey2HLUPg0ST8uGiJho2/JL46OvSf1ie6kFVkWCzLJsej6ZbCSSCZ5kqAlf
wZMQd+Ajz5h0djhJBGB3kuUGA+i5KnuqZK4o4TUUPUe2XLQkpcJ2eSA2NLZWdjDffKh+cXViVV7a
yWIal84hwWxCo6V+lNoUBlzQLRqSBMnhFLVecGXSOGbgIv9z3Tao35Frhf2iH2OfWbtzFCn4REMN
VVR5GRvecT0x01CrxGvoQpLVCSW/kjhErKRprpibut4jOPwC6yw6BfT5EjfIdIjlnoCMZm+TpHZG
BYl/LICHGyZlApyw4CHUH3owTu4hbs7y1Q79iNB6Pkrt/TI41cfEHipKcYJN24wa4GfUJLRo5J2I
Yb9p/Uo/PchZzndqmpD2sNpFtsmA2BOiFea6FxBOQoHY5CKypRFQzbr/PgqKSnMMKppCehRiEHys
HtSjp7QVDC+4yvgguc++AFDeHm3wmENVmcGwwqqSKBKBLt0zAqDlVodDwj/7RF6lan1KaS9QVqcn
0fY5v/C5vYgzHtLUpUg4d5mh9YP5pcPE4JGm5vD7R+Z0Jwr+fovJ3xeIRBmlK3PKKTWT24iIhgTg
pFmAV9ZxX8rpPyNAGPFBP7YpZHhKYSc/Gh3oGuWWOJUk/BdQzybRfyKO9SWVbeqogBPzaeuTv7Y7
rjaTSjN5N99sEkRPgweOauKnT4cQEk6qZQAAv/e7KEhGg4wEdjL5bYs/2B3B4bJFNrwlNW0rnutU
EoAy8s0KePbbONZQN7kaUDbaZsknoUOUW2tFl5xMmDxgNiErElL3BU4Txzn+6BBlwU7iIM3mvbJz
zwzsxR49aZ8FYiId+VvRlq7WWdFJdSXq7B7pTxjkG7irTBeTFXp80fPtwYZ5U8faId6x4tWxa2tl
fPVO9NDwfVaEIaLBm4ROA92lr03an5XJoOWTQm7/GTjSh68rqUu2c4/heEBkZTiUm7eS/WxoCsAE
JbkFyn7PyJ+osBSfo0nMJLV7s94a7eSkQvEo+tQI/TgyK66H46OtBp/XHnwDOz3klFEvshThOsU/
cTtHyqFwpXamT4RXGxMynLeuLoS9gIrSuV4cXMqSJR+zxQNNf4QJLqmrSLUZi/gVTweMwc5YFdg1
Rg06qoTOd9mMT5s0VDmVBcO5a3i5XKO4U3Uov9ysyUWgbEZuD4Daie6zIotbRuMXQmU+DCshw7tz
JtET3iMZlEwVMEXG0azbbS8qsQsrXByrGfTT3zzn/rlthY67qPyocTNcn79PQwoay4SyC47xbc4a
rxX1JAuvYSAPXwWsEfEeJ3x30TSS6kINhk9/9EukcMQOY0RikgD6xQqt4rDxQjXQhjyXUQSmSZB6
P9r9o1HoLMD8FTPIRC/Pd7BxOuNQWpbI9dqRF1EABplrBjTaZ653+IaU5mX0+qgytrmdev0Q3kdY
8fUGJPDdpeDwMsNcZgnuU2HCN9D4cVgtQ50JYYfvfMdamWwDC749wQqaQzW/f/Xymmo8n3VioesO
RtbpkCT6oXbfZQj/G+QBq+nTHiexq3IUBSdao+r5hWz4w1alRiZVla790UgVwBbqPHSzdv+ZHa2u
8SqEcZT2/1oZ5mWJDBUqENVQ4IuGJ+ZsvDIprllPWRyzw75MYXYvNzHKNPx/LdA0W/7LeN3gFpup
Fp58qRjBDIvJtuiznZWtcaJuxMIZyC7qLQ3jtb/8EElQIEh6Z+O4aUfPv2kV8vT2G5/9pZ1zVzAO
71DGIt0GwVdEy5gPyx7kMMv1pFYzvuNfDbuWDmsdlC0LtorlsASiltbORn1TQcKFL7Dil83f+CoB
RX1RRNYXWhW9zYJuGkFHWA9iK8lXkle5Lb4gtdse/arh394qI8jtSPHgfcNX+a/zI1DD/yALgAmm
6hlEv9kpjNdJw+iFxBb8muG73vKWXISxL95ykMn+6sBCG5EJ7kSM2PtIVIPkW0pSXDfKfqT30QZ9
VqYyY/uaUG/6xXgnhwk6EODW2Yju/S3MvRwPTdcjuKj0+7qDWRhd/hm2tgDUC4n4um0ZJLTbxDNO
J7aImajOb7fWVishZucUyfFe/mCUzoQPaCu9ol64I4gfbltXNFa+S1i3hfVv/KX1LiVuO+LNTLGm
alesctJN5/eiQJWpLaHDt+ylp8rdzGI2UD3/mVx1NNMFu0H0jZusSzZBbLA9WKTKfn9POGMEuRdN
xOoo6dTD+6/IvzenMj4diSxsw8KTPzlR5mhkEnHkpKqU8pkTHRYPGqKltc8yoImn61FJCLxrZP0g
rD8vSWHC7JnWModVF/Z77+b++24MjxtbGNo4tFXZbx+uyoLMRP8tjSOo9G7B4ISmFPOx8zszQ5mo
IQx1xdgEfCz4x3xkfz6wt7qbM6q0UQnzk6tJA5RN5kMJLHxphUYUBD9JDM59EhykXxXdebqku20n
xx8KIcS7ems8Sg8cHeRlKE/MKrtQHqinVj/qJFsSXErx9PCtWdPa9VrrTnl5ZVQTflzkSpOYagHC
XRehGG/lJmz+2E2fnIgHbOnOCjygQP6/YJh4iN+vhsXAfBEh0ndehltf8BJVbLItJj6uCAxYQj7t
Wi24zvkcpxJEWIj2sUlPQ5M083n4kTyX2J0PeoXacHj0PGhAxTS6hLDFy9DRKjuMKuytv3mNnTi9
df0hKC2jnTB+QSDGXZF8qoJOLgRgafa/+HudN2xdaYIDNhOa0gfYACRb0NaZ2CMPDKxDnNqzIOYg
RWHANdNBDBdMwXFZBG2xtZvN0h+BcoNeJssbCxbdCH7ERvsNokwYtTtYgmNINQngKlAdLZzK0wme
llEdEVB1LK8VYK1CJ2anS4tBUf2+zi47b6z6WbxMON5grU9lW3EiWLLe/5w19bsTLmsQFBuQc959
ktT/czryfdhrWfFOS3Ywck8xP1dgCzAp+038qTJ9j/yT2pcerdTnYjjJCYj6q2u/KmhGiUbzhrEP
0Ca14BOv5fxwQs7DOjzcwvKNxKIMh2cPrd8SSxDhWKLdaFdROIN34YZjLrTEPlH04ZL3MHBOSghd
o6YzCK0QeqHmoVn6hFDw5Fn38TtjFeXBeamd910GoHjYBE0ZxjWXfZ1uJB1ruUJYnY8rxx380iVG
SAvP0Fe5GkR5tLsBthGio2dmOY+gDh3Jp+8AdSnEN7dU41zBeahwNuoEqvr9trsfzHoUy3+0+bW6
7eNO+BD/+8uBEW83QDbCbxrQlzKntNCKN+487CvWdM+rhMrENF8iiI5J+jU29AQyx6KK2+QyA17L
vn0fDgRqlR0Vx8Y26+rSsuCe5Xhs2ly1G4nwJ0KPOlTgRoU2U2vBZx8K2wGVzdHkl6RekiAdckmF
TkU/eB/xVPvbgj9Ma7ERBuG/W3S9gxi5GIjLOlYoEc7syrNbZoTINdts6KeLCNCtss0IRbV8sPUw
DVGmrVbhgbYUFoOXwTQPi7AUN49kk2yG0ZH19XXDXnbTuwVE689WOjk6bQQVECBpS9BIJcVRTmEq
Z9R8xPFntc940FRezC7SK98fQ7T9lVMCXdCmNttiXSICXeEOH1I+U1LclBEFWCQhqX6sN+W7Sa62
DpnUx0N8WdpXkE23dsawMktUUeRpKx6V2dzr/w530Vn50dCJ+1nqpSU7Suhfavn0iuJmF5dc9mgB
uNB7vuhYYb0q3W0Blkqj0RFox5kY8uMbwnJx3ImgZp6TWxbCl60+0EIQvXQgdPiu5AhQSo2UJ96U
SRU5ENEC+S9yDfZv7lHLuKOQLejfB+a0YxBcE0pQLQiXo03PSF2wcfHvBEzrIb/aZ5mYogbgwaGW
kAY40A4TXHMHW11Ph8AaNZJqr6fUlbHqFYuUaeLmi6AnzsAHd/Bd18okP2xm++UJTl4Epd7r3+OL
aeOdZSHKWm3fbLe1wDodgscAr50dHK62facACQjJUc5ZBWNt6ItUEpBFi09JBfHF1JYNspe6thw7
4nGsUFfyCstFqQdfZMJOAQPgSsZeX/vHeOWsH5A/5MijFeRUcBopl9sG9rG0YAFBPFhr3KlEntHw
0iM6HmrywBSX7ZjUVVbzCLxLvxMRluCV+blcfP0dWFj0nTPBRBOyHZ/i3zpdQpfxF3veM1SXf2iZ
kTeZFAQu+X/in+9DkFb5pC7m6qJnyrlP/K4U4WjOaZlpS5i/dDs6q0qrLguxdYRwkM2d608ocd49
HFMKVJJNrqSp7yE0POhvr/dyQ/sz/oTK5wuBCqqP0geHX8E+Sls9OkCnjbjFwwmIcdr/BJp5021H
uXlF1SitZI4jb2Bd0POlj//1FPXL14sIGGrii4r1x55t36cLT1mt2ZeW+UM2v3Wd8j5MuASOV/dk
ulTzOhxn21YjvgPSOWYuqdudvAepES1ztEar3QH17Ca7q1twE1B+F/Hh8XRI2BtJLpshKoNUASOd
+/Wd5NoaodP0Et/W+rfcrMki94dgfWGFgBR7hPCbdJH3pU6SBuH3II5Db4e7TyUHEppYshsZ7hjh
edt5MWxumWLmyK1c2pqvUI906C+Tubqq25ngSduK47CT6EVRxGWq7PPL3OpsytBgOwF2+BgXCE0R
a+cdwyB71GeIPdY+RvThMipYkkC+7IMGT7qGOm8oKkXem9+A2v54s2B4pWCYyGC1dChRG1Ld7wG2
77ba38CHrlDckmFYiut7yWdCiuOQdUBsAUVgkjOz1g79V0DBvfW9UFkDCpP2ngFJUIq/Cfz4w5Hs
TkC1a0KT5RYPfhLg9DOg+dZdmmxtCqLQwV8C5/cOiRyICAl/cpXCsSzfGT9MWTQXR1Kf4Z8kGwO3
kRdrrio/rQ7FzyzUo5U4MV/dHzXIQVuxjrWjiq31AUvnE7dNlFFeA5gpR0ZBKcSaG+k92GA5KSVZ
an/DpdchS++nvIe1SM2Qni6FDrUL3MLUKftBOyYD4oFuu1yO33c+qP+ugH2L6leO4azo27tPj5Wd
v5j4JuPlEkkX3YejjoibtHhgo1fXsrD5bWev50Vdy4/hWvI2HqvHLXbb2lWiAWN5o+6q4cOQMu8u
V5nt2KJa5ttQXyB6RsIO9HhkGdnUhuCu1Y23Jb0mmZ2YkXhKtFJ0AIknDABoWzSMrSQKHaafaVZa
UdxYaFBaw98YnuA7B1iC8+t0+/tyePJV2khZUpryaEI7M7Xga2b6/B2a48e30FDen9WWYb/wGlVb
lGOk5pUXCz5djicUlp7YPHVV22B8P26xqeF14UsZc51OSEnNADVgfLhITnfzq4IoLacUIDEjhQjd
jdiFi7jNWc26eFdW2gkdqrsVSscrvtBkoH+xSY8iPu06F6et1sfJPy8Jmc+ILN5AQoort0fPf1+b
A6metV5eEy4KBBoPSj6/XNNIvhNflvvdf0SpUulfDEglmyhvK9EAON5uZiRpHXsgjxxRWUjRWasI
pGFddFIvDN4mVX1aS2LYvdZRXAbX8cXo0/5YIVQE6plMwZfPFzNwFsi344TZiA2cAl6gonqfhams
V03EnP5RNGSByN/i+OJJg8XRxc8ALUCoQQyBbTXRYcfPG8eoQmoDL24YGYRWNLAJtzVsF2g3RzQI
SRhH467r+iwMd7+Hs1ss6MD+cXgk0pp/sISEWkWj3sMfOTG7rQKPqY7E1wRfeO4W6plv076/1qX/
lsO6LD/e0Ysy743eYAKGE3AHH3T7oQyiqT1tmZ8wyscXDRhOjbKhbATfXQqT9dVeyjffchYq1g0j
Zxl+AqSxkJeWJr8vCnf1O+1049vIiw7qEsJHvimzvV5NXPrgofEa354902GHyGjRKKHzSfaDihDl
IoXalzQdOE8E9UFDC4DzIX6KUQZ6rx1ft1IQQTV+vH0FkZP0gyHbSNsdj+vhbhaau5OUXAb93FFG
ofizsfaWoPrTSGoNQ9/zHZX8yzzAqgXWIW8yJPH6ftJ5WThzFDWVqGhtdBFubSzHKrpBIexa0cN0
f5hwPhSwP6VHKONlLwvJh+OCi0pN3In8Sl5jWZEmugKl64gudg5zRB90NpjSDyCgXCYGia+dXens
qcS5rE0I5/LM8J2Y8FEjJ79SaECbalJ8gaPyqAIRqR1XPaFxqvUsEMbOXKKHn8C9VopilcthJldA
i5wRpDpMbr+5mHc3FTvLK+Oswf0vGJxHG2LevLyRSW1P9/qhwr2fpLSTqT8qRIsMrF9HaB7bTmJ5
mUI8wEZ5jcyNJfPfr5k5CoBvzsicKMS3WFk91La9PsGEP/1azfLR4KlsCLr4u/gUGFAVlwTbtPga
3MFgRk06jS/cbr0rsmuYuKiQAzcw7KDxK27MeXMuBNjUtBDxDV7b5cM/eWuWYbIcE8UOKdBZZyMQ
mdoHuYwG1Y/DNz38CfV/AmlVZ02RS2yyNXRokltj99iJc2vm9Re60NWmdl0h3fh9Y7Xjen1l2qfd
0XBUqb+qvuFL2kOrVSa9zaI/ZaGQlYxN59ok9JvwcQ2ZMIdGsm5u/Pwt4WQMu/ycqFTdIpiiohDZ
iyCDMLVPU49RELuxp04d6sByJcBCO7Scx8i7/3mlR/sBRmXdRtwGEPfjIqDTc/WExLbSM/MY24ya
8o8bs0C26u9SnOXvCpTKnbsZllkufOZR7vzVEgekovAQiWX9Oe6cJN87uS7+X5bmoE258BnztB0j
PDLpzHCoa2Tw6BHVHsBpgAZjnqm6MJ6vj7/skLcMPj76dRScydcjOe5kx5DKKtNpDVgeAgeRMC4m
sKOR/rzZWXhRuwlSc8EkvRwVCL/oe+XYxrS6zjR1OCMDCU2QMkJkJxCR8eqqjxQRgY7YVJkc2I6l
zV4A4p+Ofv4wSKJ53sPGjx6NGd4yoWffjY3aTy1I7Z36mKktSPAD+vu/O1JNjku9XlZ4xnM8CwOC
WrKDRLpMPVwWOPKS/WTrke9l9LfSIPcS8Ecbl0kU2HERDElERzkIy04ovyl+HtGxyNHt3IR9P6Qg
znz2aR353zS61On7hVeuHdndRaMYP0v4KHRKy+9fR8z+0mMnv7PdbzGO04ALDwd1UP80CA6EFXWJ
CqdYRvE6l16OywoJ2GyaQ+culfEsdRemr1Zs0Gj6ykDxMK4DjomvIdl0GwmQXBXzvoOjd9oxl+F7
DRemHF9HAp1WYg5i1BNIxoKv9ns5DHfRU09Y51iRObfVKYVWKPbZzr72HTvJkn/3K8CBuVooloEp
Gm6OwsbOe5EtQfw3Eo93ano6k5QoCt6Pa1f5SRCY0dI30NOVv9GBLmnLq4JEpmEfEoHBZLRpL5CZ
aRDrFnMs5t2inpZRtYWnpOi1pW7jr00qP1sJGxduGnLDdQp1AwDRUSMJoOXB9P0S62eg1ZMTYa5g
GdjDCNSwr/5+aqzJX6hEQ+AaSebEfnLyBwP7hq4mGpcTAYyvj4oe2FVFdc0C/5vqxbTQ6ZDwh2wX
O9CnJ6u3Sxx8S4yvvJeq2dFW2rhA+idSPJv0NNnC4ibVt7Lzy/yotrCuUC1Qekidnijc4g2OeJ9y
2dMjsEcn8R9iI9fH7SZCsGPgrSzMtz4dgEotyLBfa9C1suoeXnCxKaYpcgrlDyoT0uM9COd3H932
cQdTpS9j40tHEyY4R83sdUww36tS6XmjqdWZROHH/M+vJ+CwE69DKuEFhkKjGfbuioUsPoU2Fg1Z
s0a49IMlGz3b0sN+RHFJ3ZtS5s5qiNd1JWWj5Ckvo9LRhd3jHPI93q6zVlU3Gy8OGuwIzXBGTAzd
CLSNcjsqUSXP2HWYvttHHJTrzi7DW5hRVjfk8xugqE4IW1RgFS8X4+Br40Neq82/CVtHMLHyU8H3
OT3PqvDxMj//EywjdIopM0kIy/R6cEPyzkGRRD5PVNgwto2l2zsW5DSQluOnNOgzUkMpayy9wSfp
MdIy5CucwL2gU3ER+FjPqQ3yzi8pnmQyyvHDLJx28/tU3EyqkoidiZwUe48RG7RRFIJuBxEuZuuf
0oP292Rxi1HtuY4yWs43T87xCZeBekPkornpRPCIuk99THwQEuRGPtdMbUXym8pR0gO6AWFHMaEQ
gXbApztdkSsG1qXzedOrU+x6ZIDyrS7l8PrBcuPap0fNYhHoGcDsNY8KEzrR9Mj6z/wDDbmMfmQO
IwhMLapNNsJ2/L9G4XBXiYXqYxmZxpXyQL/Br0KjpGfXnJVd8IRXvuS2faT65Utmtbs7LRmp0LpS
sZi34hlnxJziEDLDybd+06duRk8dWJWn4tBQWf5zaakcEqMCneAfdUqRQH2XxZDJBlPyAkaj65Re
8X0QVJUd9hmHvzIdyf+Dxti0jobuoliVP5hzWciHWmNqmE554/mKcDAYjFM2vq0ISaGoN9WdwIu6
O6f8ZSgU2U3KqaDwwvTIigrsJ+D4cLvlT1wp9kcrmw1K0IGv9H/TIyZlfJW5U6V4xNaz25aYRNWK
DlCKToM8i4r+2ngtFBHoDRb6+lXwyMKrqLlG0JRojMSmP1lFsrDKx0RO5EU/dtitydWAOfNaKZDn
bTFZ90x/S84iXDagrDqdWQibDeN5mJmgMfGbJe+YQTCm6Yy2qwIi7OPi0AyvoeJ6NUmW13FiuoRn
XeiK2K5nHNKAYdEK2PB8Ax2x8OZWdobwKAhi3Q3ep96uf4DpSTtqE3NuEwFlbttRq0+8nGqWEXJK
apFbPqJSPWw7lO+QbTU2bpCr62CBwm60tX1R9c157AslVfH4DCYtQxY24K44nvaBcgosZezGltC0
48PQFg72gOGcmlakMIimgXEgpBrrEmVdZltgtz9KyhEP80QcOdKYoOp5yYZxGX8HqcIdl2VMMxV5
JV4mK8uo8HY5+i4n0spWxWX/h0d3iZKDfxnO22tc4AYMl1wcROmk48aQETr8LZUAXGnx8aJCysWE
7SPw/ijBw+Fa1x+ArUMfaVCFTueIxXSEVH5XIaY1Bk1zocdWL8O3m0szctlZaQZUmlplSRbbVO1T
Rxk3KdtQGCX6Hgo6tNFc1bzeSHM/Z+YUpQKitxbKexjVjEDPio8tcDXgzfY3ZszFevbmx5LrbhHD
yItPJX5yBqyRQu42V5RR31omCdc38hRm8TUTLnFj/JvyZGuLx4waYemTjhsoJVIrhMAratewo02m
+LnkNcteJHZLPzZA3B03K2ZvBKY/4jPcZi3fF1E8TUiot/dqHqgIegZ/BPM15ZiIV3aEMEykEJgH
npDC40PrMpuNKbFB9zex+32FhGb8wb5Uo5tmNKuV/bORyDYlHTrZcCK+Wr8BnxS4/0da30L5X0DN
6tbqX/ChsKRCewbHBI4sJwRNo6CQ/mEHafF7hteWBHenw7e8Pcxi9GB5oxNxtjUrEbLOpFfpJgLy
eXqWKj/tw/ATsWo7igWadzgSp25aeBpG+ZkhAUFW9z05WY0mTuH2bLc/TAzIJFANTdO/hKkkI2uD
RY3FoMI9Te1NJsfxSw4GznKGvNyFD2O1RTFyhxqcgqvaw1uxjSQn8H+9La5BVYwWDhjBnwQRuPqF
WNQLb9aJdCQeVSkkb55pvW97lKvjxQcC31ke6zl1bQTt4bijOmC4wxMPc5PdOPQyFSfl9XurbSq4
r7r9aSgpIMvaSgqWZ9XpUPpWQymd8OvJGFikTi0u/RTzYXnLH/mBUANoMiSPUc7GCDWCXy6tFYYr
XZW0TLEzosDV7tHXFVaaAvwUp1sMsZFQ4z+ism8l3+LoNtaQ7j6ySocgOqLL+voyWOID39uTY5Vc
zhlYSh/kWY27fUGv7V2VPdnNsNjp/qDTdrG1bUFXwNk259vew3NVphDOnFZxmZxCxdSCfM4HHWmP
M+6btfFdeJiHEnGUdMaJJtqhrTdh0fRbfXKXSKfnqqT8FA3uEVV/nw1UagWA+b/3+K33K47kKECW
558XgHqm/w4jgMRHnfc2BDWuNmYESSIJoTbJj+bCTT/12uoFtxmEEqa5kjl8rpmHolwLOnbHUU8d
F+xpO7MrgKpLrGNk0tjFPCoxlDrAq0MIf9lXvxd4YXtL6LoSkeerVJbQc2sws2DqvAVVitA+KqzV
tt4Yt1cBD+9LEv1EWk1+jly8fZ6lG/G5r4lWb4VprEP9tTVHV8fcmw2Jpzijt4S5zydnvLxzV7DM
S7fiJW2t5BBawfXM3qKFEHyAypD1eb4FzCljmz+QzprsuP+xodZfNAeWu+QZZHsE+0pZ6pabE8oL
vOtcqy7nJ9olM8IHriiJWVM9a9DSBzeSyhz15RzsgQNMCwS1X/kqPHzSKBeIgvWDeUVb3ONj1NIo
tY8jX0HfTHpmkjT5V8BOvr/ChOsra4iJlqPpGN5vIJi4n7UmuGMg51F9Qbptdb7HJD+cQH+Dc8NQ
VGpT+Wop5IC24plGvEapPf58F023Q4lGwkVBAUQcbAVQtGzGBnATdcuCetkBrolZg4NqyF8kVm5S
drIUv9LpYNGe2KA5qR7m99wrJuzkcDns0LXaDRtdDg0kYu6FaSenoL9z5lRxKCYjzjTpwOdrhMpQ
+i9OeaSZ+vS2KFHT3MdZdQdU8iBMzpSc+27YGPQuCgJaguR1uDeW/uhJnrnXRAyZvmj9iFjhstd3
Xk9LGl97KLDcP90t2mam015CmkK1BCW97Qdgvckk8dFCBy4ynOe8tXTzbMt7hDkBgRJn11/4Qm6q
r72JAVTBYVhhouJgd/eKdB4krDbHJtlH8c7EnwSXe+YQ8VOaivugpJDKC0AugetpnoGEkQe8+i63
zXVeNAVFFeLJ3cUnmnwb3zVHUMxprYaI5paafi9vqWen6qbk7GPu6OXzlALbFmSiEUKeAhlh+8uc
x8U3enNj9EHEV9EGiN3fRCVs4Ed1WQGvXi3KqXa3S6GdcO+IGWfuf1dk2rrVAw3uPSOlLeJmrgkI
p4PITx/J/MQm4Gna/utR49zKyoNuoY7IHmZVB+owqRg9rP53IaybD6q813uAf1/f63oEzPhLr23M
6VROO3uqLr1fPXmsgpJ6XOP/OXIKNv0QxJ8+/jfKu1Q71rxRm+cycfqPXKVWu2hs/1/B2jzQ548X
ip3Kkkrx1g7eM70Pw8uWmMGCieicXoth1OTDNSgi2RwqKoCNLeVl9rovTpLADhdiMhxMWTL8bKAM
ICei9iEreOu5Fy+60g0vD9hcyY+H/olcdT7nEfoWiyEpu+BWrnQM33E6zK2MbEITwy2kbjONPLhP
WQheplAyYjn0JqD9pSs6R7qqOkdFI/vifHB4W0RvEtfUUpiq9cPkDueOSvDwmm+L6Wz2mtzJP9NK
4DF0ObmfV3TqiAQnAjUsYHmvPKyCHKjBQczoT/A0JTcU595R6q5L2esWmZQR2axxTw2p0/lH/xiR
p7O0MDJ7NG1WT9f23PNhn/RnQsNLU+6jFxTAoXhL7Lz88vxHDvw4+Tcy8ps0ZmPNnQIIj+tDn9oR
XhFy5JHWIgddrTqPkMahcBH1xKwPgXkQCpNgA8i1526mUosXE1uBInbdmOTm9ad7FBrM5uYFOEcn
muyX4guk2oAZJMg/WOJE+5hQ8grBcI7GK0YkaznMrr3rp9xTqblWCAsS9MNTAAtlJAtheTBBt4Zb
yrCrHTSmnUUFoQ+oGgDZtFKgKutVeFycGEpmF7O1z1imsbnS4tAL5OGaAxe8bg49kIbwUm4K1o5i
WADvGy8yO3jPROW7t4QGU5j/NQv7VJ1FBSKu3HyJiHxF3Bvq0Ykis3/jnRlbyQIf/6u98WnGbHvD
VeHBwDw4ah9pFRlvSAkkUj9CyTMtA52oNY4Sn79knsiJpRwbXhWxM9JC24Sjw/FvdRQn8lOX9KVO
ewuE9PZ0M0v2aalFHszNu6h5JQdzUsXyovcupa5YUGK44RlCLPWRPVJkOIAtGEuMGAdS+yZuluVA
rj/UzuUDSfTPwuciGnQBCSY0kB85Ha9mdKttmB8u7g9xdR0EkqAAhTw/wUTb/byIwfaVFBGxRfVb
oqP1sgaLNQ5xG2OBdVIrxmq4D+k05Aqs/lwkgD7oS+5QvTzTyS78ZGOEVGvf6cJg+qjJMI0vzC8b
hm+SZEyeRSJlwaaH5X05piXeB6zhMIEBkuPAk4XzLDk1JiygazjFvdkZ0YiTepnWG+yA1gzJZ9s5
KTRlfGHVBrFDjF76nNfMsc6J5isjYSTgczmAR0sf3rjPLCi0BctbBqRmRdfggmuiDs6FO6sjh70C
TxDbe0wBlsoek4gL+oEvHXhYgLzit6hJPSVjuB4E+UmTx0XGFl6XDngsvad8nC9T/sqE7LBluFc6
E6cu8y3PYp62Gxd7K8u9kgtkIAX8gonuNFQQZxMU7giXD4m5w0HYcN24KappPFWFoeQ4fr1YsKjO
t1Lx9Rq/s1Hhpldvsv3ohzcycWo15nLc+8qiB1dbNzmgtVAV/Qi45aUpU2dGorpCvuaBZfxxHUY2
jckC3G9JYXlW+bvnP/d+QlnaLcLiAwkXLgmfz6PahHoFVnKALU370Zdz1qnq3eU5DrF6Fd9iOlxH
Cwgh4JHy18K7Nl+P40T/0tNelwzFelRLlRHpCQO7w76UDKYNIoLGUsAqWWOPB7uStr8ot7F8ZJsd
jAjNZBDpYcCbsA508Dw/b2fId0cEUqfi1n9GyvONKP2vK2umXB9pz5YkyMmOzbLz9qjBsMRG5Qab
V/K1DHnSQFeTdJx3JPG8GX8aNmOd84y3czOlxgfzqO/laC/R00c7YiBxto4XRW1M3Mg2dEUIk3Jo
EA5VIweemNx2uwDF6K/VDVOKNa9+Lin67vGKtRb4KHgL5P/Otqpn8/iSApmtv4rnNa19xCRBLnrf
i6LDe1MiHEITWRCihHvwgfecbaNXoSaag0JqZzi0Er3UiEed23pG6J4aVneg4NUCceTgHX3XbH4S
QkDf7u5GIERw3D76F57vVUBNJtE05YQQz1RE0vOEZ0ZAYMLdWcFP1HzgzInnrNC4X69ZbuCht8I1
xsuifNcT8RUY24x6PisTqLhC010AedpsTcv5VoGt5JhR660Pj+VYWs4fTkXHAuBEFd+mGSPcRv0d
b05nMW4a4l3GO18rC/Qn+hEr8HwrUU/qPdoZPouuuKXx+MyFUJhiZEvhXLaf9836fDoQJhOboqcs
uNnt4MGylx+6OrO0cv91L8c+ic3s9oKGEwjdiSsvOxkKXnwrKDeYq4uYp3P/Pt6B7dGFcR5uM54j
dI85Yu0QuT/b0iZOXjWveoPcLwYg3LbmNMW/bFiqoljO33BeF3i4AYwYZKU4F0NiOe+7cMQWD1f4
3QAAsOiKsTjKcvtkK7HDxmn842bzEboSqiiaaOyG2LzfZxWcmjdfxb94NWL/Frajp5wT6c2p87F+
BH3SRwCd3pGJKUgjs7NqMRXfMx6po3DASuNxXHhf1kiyMCplCeu20a8P4BOooq0DBDBEs+edjBDJ
xIxmqpF7sIavI1Frpjpd/wyjlFjHF6Z5ipWayx7fU3mnOxcFkXNfc5LmjhpWWsxW2kHgUh4MJybZ
89KYPNID2F1uO2F4w3lvW9EaSBLzCpx1LlBpqRkaI+p9DgepNSDiEv1pwqq0LT/ABRDPLxVPf/zR
juVgnsyvHS3z/cwR6iueqnTA96MYe9gqq1w1aZLbycv2jfCNSjrFuVno43XuK3PDsxSPBJ7xrMVu
GtVjtEZ5we3yTDUiFRVKCiQ4fHsevRUzrBjpXEpE01gHxAl6VwKMnBMnph+HAJewXyjHZMSFxxJc
LKKCxkF73sQbpICzroPevpS/33on8xJx4LeyaBO0j67pFfWG0nsPfBXXNavhKuLbMRH/dq+TKF56
HKPFXQPkjCS8HgZtgH2uigmgf3QqR5bKD3Pqy3bYbMsowYP679+c4cD1Gtf3uEPiFhsUJ6weesyL
9QPFuv6SKDx4Muw2ScXYAhO9nIGRhYzxdyC5GAGPMv+guUjgNHj4PNQVEhLKZ9H+n1rvetzf/XKd
1nzVxhBz1V6mPivu/o9xRzZ+HcvsbezJDTBcTjecOGlsjaTevOr4hpDV952sUeKvFiUtSpugVIHl
FfAQtZTt/2rB1riPPBFNSlo5UtLOcwUo5mAuoSwHF1phIMiJj3sHkMAcgOA+U+mCPFXqptsPlelD
935ZqKDSPmQBnt0GNJdaHEAq4O29NJFg5QPi00ThloPNAEHyNbJ92jD204AUu/fWQi5o6pEtyA1e
kbvUMBceSHHuYlLAVAzgOMLu7GQWGM0b00TYlWDPaiEbJ8MAK6LjdfzEDlPNYBEbXrNrkRZjsgjR
yjPfpuVpgx0xNlbeLsMuXUzT/Msh3bO3aaZfj2926H+Cko037E6a+GqjuCk3hmav1f9OHDaxMkEQ
V870KWFrPg76mD2XsYTQtRhPMI3I7GHp+BXxAgYJiNw9WEGcIul9o9Cc0bxS2sKR01AtpRs0c0GK
VEB1X9eSZZpxqfLJocfmHQ8+o62kad+8CLURuLsdcxDt+kBm5RX/i2q0yTHMKDNrXj9HElvRMKWb
9x0HU/otR5UgEow3zsp+fDCaKtT2leRqLkaXZoYAWa4Ef2sT4HOjxZKZcw9ITjp9bhOiDQJBoKF1
JOv375hB2Ar5sd/oPR4wGgjyOqrvpwIPEwvZpFiOBCpQoo22ZlRO0p+l2jb5NEprS/tfYtVViobB
MPN+KuAFfI849sJUyLY53X6Cs4sX4li2Ql+obLDqWPxB/rBRP6tbclfcSDmVVWHGpfmkKNZO7i7b
M2s631bh4w2DDLYgVBu+BAKca9zjvPoQXbbvrKAr+VU7TW2yEeymVzVaCigkPEmTXZy0IOcAakmp
21ggQa3tIus6QRVgdGsYKsDzk/OY2x+1GvfEUK2Wj8QHrrNt4roqeTQ6K1kQPdJy9axnUrFcO0PC
zi59w22+ICFmqxUu/4NbPuIKITsWM+gC4d2FvRaIuejSKHVIrE0/OLAmtwhBiB44jAzM7fyCdljc
VhP0fAWybSKGFgNBopzb+MpohgGpqrX/8CCkfwXbW6pMtVp/nXrvX2fvFIqQXY7gBeYzCUEz6b6i
8BvOGjoRiht6VPWIdFv5GLer99eHooBRVtDusL5mLyv+2GWohagRmmYQZcyXj2Fq8dkSvwOdEgSJ
4PjEyqq7MJ/Huair2ndPVja8Ikr9wKR93Zo8VfytmJMC8KOuQvydnYUDzEUXFrlkP79jV1h6l2Al
9dwTbOADEimVBYHHRnh4bio1pt79PFZGVQ2KVKrcK40qO0AzWgX28zUE2yaiRrPXj6hw1IDhhGoy
Wxb+2Lb/KwCuLUzJp2tIomqdGkgoYwyyaG2sAUIWxOVRb07sTZk83Bowc/oOr5/U8sdXRwV5is9H
j87Y4OOkrBNOPg9II31KrKU1jL1Pc4r/QJyMmM9DSZPhbYAMJUdQhbMPl0VOZT+I0sISem0PBcR0
BUDy1G3XQFSL5hdnsWvrnS9pgxpqshqe0RHa+J3jYhIH5iSOPfkv/j4mtWEX9S2Ni/31oDup2fA/
+ptYFlVsqn3O7gkY1gTd/jtMnUjioKyRHPPRk+Bhn7hxQOskFRhZT6ugNCxtpsiuexyNLjm28JXq
ZvOrx2RwScC+OHMU5PJ2t8KoF015RSJRj7nmrdIj8n9tiklb0oY5ISsr7lt62hroNnFYFOHaloRG
GwRvScSZgeA2hzRAAZR4t2Jde+gGpQhxCOBYcBZEKKuaMXCPxVno/gw8ERxAoIJ+DPNyqI80Kukh
nW+NnPcKtiidiAQux9JZw3bRyPjY3ROmLdO0AkJWF+G7AsOAxCMY0uZerbLAXg98QfH4Hpa4Ov5F
b2phSe07yvuzOv7JrcxJlbgGomTt3VoQ+kpG72RUCrzhdsZtWKAxCYvEabYh25rMyrPvBZkoq3AJ
z7WrX3+W/r7uQRzbeq3rAiuxDhSw5F5oqP1vwTcspMLVPtI6JendYTmjO1was3xDOzSCB2Tvsj/r
JSEtL4F84U2AkrkHE2N3lH8W+VHtz6RxmZGVUfHo5ojBEjxfoVmtd0IhqJ3RSYImRaM0JGrYEcLS
MDFnFI0bqriegehqVDxC2N+q1RU3js0iQ1XIhjfOnTtY5V/X2NzMDKJbniKy6UjWQmA1xwhwSlxk
KkyekYgdOwT44ylOUEXpXROTMyyG5wz5UUYtrwr76PSIlZkdhQJlXtaVBtejrqmcd/OaqQT5pebq
IPl5rAu6uoq40KioN/ltsiv50y3VDFoEFOv/XPT9YfzZLGlAG3fb26a1q1+N0GB5CM2uyIglYMux
Vbt0veFTXIuX6nzQc28pGRpGYjggw9bhnRaiAToLS4UGPcBSe5q1ulP144HdJjGY04j7hxfJeOW4
+AwZySQ0qMY4DhvOc16gXyPR4nhL4f8yxHGIgWoMK/c3D+2E9x2dZLBK6l/VF2xnIIWzY0uw9KeV
kU2e60apc/dBPt5Q5x6/Te5ZyOYAizFBAfGS0VYM9xd6ugp9y+oixB2m8ulDQGcaECzXcqzm8WJa
qR0OMeS91AJ8Io6YbX9VzHw/Yzm2Ol9y4oVb+x2BKS9gCkO+pRSSI/wK7aenwwZ5dl344NwA5c/s
k8NgeOtDdnpJ0jxWarx6IJj5hAHg2Fj/3zLN3MJ51BD2nOQqdS2e0Bl+Ext73V8BH2KGFUv39tlu
IYnpUMv287aUKRtRzt+wUMSYrZzfLLTVfzqnOXfxbmRQzqwdkq/gyWj4UKAFkLY6wrjaZXKlgIwI
2L1NcO2iz1Xk0XFEOMFjPVgLWFV90d7p61Nf/Q0st5L+KoTyUH3qV+71MSTc/953eLL2ffWEJukI
2wammGlGaoiFwmWoreXd6QrTZnx629LFCatCboFESlf+P2rtpcfAq4fwyNeizqx8/X1EfjrP3E5C
KTtXhzZapVk+lBmSilXFwnSLXGLwiitncTZ+QDYPv0U3pg5snqOG5wxdqAetn0yU9FZKuZE1LcM2
pTFwoxXpTu02bYXeg3LWDw6VUCwTSzcfYtbSP53+64bb5uqRdaCtJsWG6Zw7+N0udkoukkeQsvnN
GXbH5ghJdGL2zUQCJ4bxXJTpRyAUgELYNnI8eoOvsMJgB6H7J1K6TOt2fzedm8FIC5bW1GI+0ePQ
FQ1wQvp8NaG/gXR+/HBTmW12r8U7Z7jamOFa9/XxJPww01uWXl61SY/XGbuJanfiYGoER/oOBSFn
A3S8ApjHsPxpGg9N/d7QeBKJl3h/t/WoNKmvVCIYCdMicntWzc79aPBoJYydRrEsjbhv5axAXEsK
6QMUkPxxeQQy8TeJfgD/khO4+hKWCMe9GanzGFHxFnc88yOvvIlimA+APyjyhQkT55RyEYUNfV/U
WbHRE1o/uKblI03Wo6RHuNkxk2+6rLHhqV2wm5FeD/INWeLzOlcNwRrIJEvbYWXlHSaN1Yc5EzVG
P8nTxqmVFGLIGoVh6LxwkyOvkXiGTbzAYXfeI4AhL0qzAuU/IJDg90X9+VRvDzKvnS7ucd6TOkhR
IE1L1LwxqN4dq/aRyIIESgHUN+WRhego3BxUy7EysPFvKymS17lREgT8OJwmCFRu8hoCG+r8N+oh
1QDcCmL3ZmxauXczPSFAF1bq04qI/QTBKzgN3g6RjN6iv4B+b2KQcckappDIISGIAC+3rQR3L5UW
3+G3eh18PF9Przhgz/RipU+qb9VxfO3XrHkPBo/SJbMJPct7uvSR2s5uO+LvLeyXDLQgW80nrohn
97kOVydUFEi+Dc7ECgnTQuDUjRtKn4WoFi4ba3zyLYDModuvkDN36Hm3wMWcA+JshgsQNo8akWuu
As9j/0RXhrQG1X4wuSeesKyd6y+JpCTreCgqVFNPPU2tqpFbvOr4LSoLR+CW3Xphuj7UQNmd0/n0
LVufJ1Pwtk6f3twkuDK/aFbP6U/gkxhfq+OK7UcYBKRmE51ONq6a8Ft1RWsQ1+FCUf8IBFxuVxGr
VTDjh74opk/GkQijJiwG2h4ssxElpuQJ9afr7kq8OteFvy0SyVfiR9XcYWKtSF9daM3V0EKLv8GC
toLLKpaDiIzNJ2dNV+sDzo/dfgsOxEmK9nZmAQ8jc0xHCB6KdjlklQw1LcCYAVnR8zKBIMTHKP0w
0gPPw4mMo+SXCahwT/waXe/Dipqn+c90nlAIFQu9q1QWFLMEc2dcRFu/O6ZLzPHF0dVqYkblwN9o
BNNYhkXOeCZ6ChpV/4MrB2I8+yEbizt/Uo6mgT2Xly20BMTZtgsT/IZmK2MTJl59cNaHNPmcAqR3
zdzgguH6dur1d9FE8Vlu78efoGpyRQFy0I6C/fRBCIBvpBo1kb/GSrLiqUQ/K5jJpgLLCAbJstwk
4xGH1RLgMJyQLgis+yJSRqb4qpWb96nqumWP8oc75ZoYcsix7LfzBvGa7t1Kx9gtIkYBgQ1KS/fs
vpISXNzog24KLJiL5bZXHNxzviVUJDpBC7DOghPyyMShtxYUadeL1XvlmPPJ8yoPEBll+zxDXM5Y
8aHkJVcT2RiMUES6SjYl77v75KPoAjCgP0e3eRhOmWdS+1WnGywfafKEe3RKPAbx5GkwRAjrLCUm
fTjXGQ1zplt2PYhY3r6Ju+SNUPrHCKFiUFdFpyo/0ZECT97BdOE0mm8H1Op5B+KAh+v3ATmC8584
C1dCjVpz1GgmdMrPkWDIAY2PTUgvfFzPF7OJGNBvVx7R08uD6x5F+DIXupNopt9ttoRjYCypzXO7
C+N/PJgAr+qoFsXaTjtgmfqDxqyf0UBnuKF++TXi2e36F6PQ4sQkzPwMUwsHpKfQXsM8ScCmZddL
C2dQWnuUjRfb6fuXHqZcY1U94EYwGqxuS6db8lBPphrOILikofd1S9Rv8DZixfqUZdWjNPAS439A
fqVgx/rVhAn7jiTVFRtrYCOL72IXRkVm07O+GwaYrDOdUQnNs2iX/W3sfCHUFrMI4d5b/DagpBub
RDitajJRRJ6ltc/4+Y+RyyFJ/CwzJfoQAKXQ7rhY5Wly+HxSAJaf0Fg0r8r6X/ZCfTlRZFPxTcYA
h7415qlLRUmz4ijzLIUjqS78DEcYohahVeT82cnrDqvJwgV14cm84kyMP4ljcH+7e3r4CUd7GtRN
TvzRMI/JwaYenaMxy4N4lXQSrRarphD7cXjFe1kUsEsreXCCOJgJ4FcmjT5EL60QjIh9Rvv64HsR
ICFg87uZEjN00RoI5sJjBUAxHhj0YsSiL8R3yGIjNL4Z+FyuV9RHn9M2EQXj6iQC7pOPsdXxGE+B
T0W5hKGUsGasaNt5JBkhBznSQ7fA8Ie5viHlgNGgBwudM15hdPVejSvHqMfC29QXKEjeDzikytei
3FweNqwxAyn1w50XU+QvrS1iX4C9kFh70peUl8KBROnmrNp7QUNJgOhgFoMlQXlNxzOT0WnTYzxt
1a0cN5b1xwXDsh3OKGF+YGaszHoOyeMmRE/b724OE5yjT3i+71jWvhFZZPpY9kJVECRRjHDzulP0
kigwTM6CHgZCtVmEWYHBNu8fIZzT8+z/8Cp7d9Q0RM++bEVKtqdaIg7XvBqrGHy63PtwEULnWWEl
daTS8nlEvCOvRQs/R3osmannqdEQ/Nm60NmfEGZi11WVJ6QU0VWrgRcwO5JBH8M2n6VLVy/Oyb1+
w70pQbVy/jd75RDEEBsDKjCcqPaQuSAqGCXk7IHucEnZA1PlZcK21kKW5hJssdkRLt3siP8p2czm
ZdRDx6ysBx6RuaGEtqSX1CyyOc0MZZTxYFNPah9T59ey8/8fmlSSvnNsDGNz8O6Tq5aJkv33S+L9
6ra4u3KGMQPOdiMMIimsRkeaKT9zcV/Q9rq2HdTT/oi5feQce17aSuv6wNnWSoIDt+AchovORrQ7
ogatP+qWTSroJ32gKE0IasylPxXkS0xzC6q66I9qtEII+tbIOBEIew0U/KnvuJQ6lTRYSl59jIEw
PYsO8/LWzXxwrs6Qib7RzKl/qCV3ieSvP9u1r8JpQ7nlUbsGZy/LlXJs1zDa8u6Rj6RSqfm9dlbs
H9rzvDU2yi7+sc42Fqquq/Xx0VL+YkMd2Sc0dP0BQDwDhgei7KsZXhPJXyWP04T1e0oI2Lu62hNQ
U++72Dd/ZRUi8EVsxMr/Oyj7er6VRTS5XaOPU8SC3LQVm9eoUpjD/AqG3e//IrN310HyITUkPHMG
Ze7UGbApeQqleKBaKXYEdXp16HQ/NYM864268Q+WD778zsAEgmA9huOTHXDM//pb+LhHQGQEMIdD
aM/CjAY2bEb68WJc6FCOwtr1ZoHtOvfyUCsux/BEPKvjCb4FLZJVu7biVevsXClQhEF6L5Q+TRs9
n/0lp4HDXtyFHkLq8dWijOubmI1pxNaDjuMU8hygMKnMu0NSfxzFx/zZeZBbpLCJGTfjJjggv7UR
aNWTz1EuYhotIR80LT4LlwAp5VFAM60dHpkE4SrIpNs5VnYD28V3p/ns9OVafD89SbC/yvNQLNgA
Qm7nCQe9ld+842HsgjP8+XgQuBSFKDMbN024rLuW2GbCZMmTPZWIdjiUoiv1a3f6XxO5OwOaG+1u
jSYxR6IOfPTY3myGYyHN1bDtgU33a+MLy3Xn5CD9LjbCArAqWeE0O2Crpeg3ebQbTjzTbw2UEej6
4eB70GRZf2g+o6RVqSYWr6Qmu5pG7l7vcIs4Z8CrEJVTd0zsdC+nmLX0sslmzZVXpF1HMvGLlv8+
ACSNoMiNQvisfOrD0Icaa8RHboFqP8JqO347fJWkRDV3QBQ2FddjJjgNKsmVA1ry0BvcoFvp5dc6
Q22rpaTJ7oBQuYKkQ6wJugxJRx4L8Zcfu9paD9yNQdcKa6ZdI53CVKSXdeQmQgu+4Rzv4cYmqwoZ
F6IEM5rV6HfDHqoIJlik7l40h/Na7C1jRHbVaXQKKtlN8Is76bAM1BzfUp0OOhoGWGvnnf8RB/61
AL/flR/DYrjpTyyge5PlMzM06g2FnZSJbe4IsRRRXr/w29Zw60e2QpjlVd6kNkMLi3b9ez5OcZLP
gAbCF1yYSoHAaqmDmRGsCBodUfN0sBlmiOtKPffEDFkob609QZjlwVLe07PAQdr8+mGE1QGVqQDa
0DowEbyrmG+xzHYkmJtnDGEuttjBkJDPX82mA9X+/3mlD27XqcmE2XYuecEVTDYEieB2ytyVzNl2
zjM/PcBnSJqMWcPPD5TpMPnkI3JcD9WcxChmyfSzuL73xD8sqB08aHmKckw9eacKXiTgcq9hzkwr
tGUpkRc9KP2T1r6cCzcq3OJQTAdsDy2er3XHA/2ha/ps3BnRsyYrrWtNuTKxd+Ckq6kAscm4zDaG
Wwo03qBRc0eHni8R5s7WZnSpHJsJVJBgPmf7Rnoo1EmTb9GVyzwuEldRJBRAmKvAJTxZY+dyqQKW
Od4L5cxfvOlwt1rltW1mzhaw9fdWe2eKCtw0j8t050l3Ew8mK1ptYYD84e4IN3PhGZUxq8PSQwRO
mg20u7luJXW0vdHeKcSLTdtPNA44TAb00tjNCKcnLf5jkfSlMCT2U3OcqOi3mDnXribJ9bmpnsev
5sQQRsyD/TB2Voo4JC+6/KaMlDTkh+PsYgvFsYEWtf3LlLIY3lBG8HdD9yxUCDWV5pw2JRPuBVGO
Tap62cp6DPEz7+SVwLAS5TvOeW7+EolCXSmydMqiS/yBfv7ffXT11fsGtzorm6T9v27BK4fMJn3S
yAGmkXcRLPN7x3+HRYVCOYgwYKsC1zrjR7DRxegGqxbJMsP0EUalkerGG7OtYa3QB0c3arNYIVme
uv4kiHhDCNDY5RQbblW3HSEJEfYZo6x2PFAMpcCCDvPWhLUhPQoRRu6O3O81z5YURARs8yXBOOtQ
s7hsm0AKkhJIZ83q3nonrtsHtVC3po+0gzK832hIE2zwLKywnS1nsM8PHFwkSuXnNpULQYEV3IQe
DrEtZgq9mHRN6Wvr5YOPZBRfr5cgCPPBA7QJakZIVSpNGp8N/SgX8ldBhd66bY1cidiBd8Yjziw8
FiyaGxkSKPjQYS/ypQxYdP5ZvYrFe4OWp6arpdiGqLmbG/BZhE6YlKX3tyRJLwF79IgPuF/uiPf3
6+BsYWYZfSmz65dw6c3oYOBQaHYg0tucz0h+MmWlHkfSfSBMmQAz8/joTuy0/PSL5SASy0Lb4c4F
S1P1E7I40AN0zt97Cc4gTFGIm+uGSNmBfy/z78YcY02FGh1t96waUiL1yVldxRWIEa+DtPcEf+G+
bxtWjuQSPRvVZQM3G6Y0Z1GAwZcB2pYydvpwyrhXM9W+ii02M/PzQOVBM1PA4TV2Bw9bNhOVCeuW
GH+otz6dn5QjSEsRZ+crgWTSPBAjUSe8defkdku9b1+a5ozATsRXSoW0Sa0aaItb2MTBKoNPNBpU
71Ze9SKzV7XO7/xI5PL1894a06G8eASjaQnkkWxSrW/b5sE8fv9SNneOb+g4yrOa5KU9E3Cq+Dq8
qDrt2U62mebF7EY4fa2kdYLCFgUj5QvaXWeYWhJC8euJNECCCtBsBRvF//tG88r5B/4QicKkIYUe
d/DZeAjYQcz+S66ScHILM8sM98iU+6F8no6+cAwcZtEd5RqXleeLZzTLh9PNMDz5a1W/gLpTp1tE
GwsbJDLFFd668YM4OCNP7UCvvMQAgtyYEMLWIrr++D9TeMqPHLdlGi5MCeJrOL5JLVDxHQBQ3AZk
LE3hCvs8m2vqAYv6f1hlXxmNlXdiPAYhY3OWX3smLbUDBLH2Wx1I7OiWx8ASl4rdM6Ixzz3W/3/u
f7iAOFmIY/U33wHqt7RqOp6J3oGi0xFrnj11I88RNqWfdhR5yX2Q9BZvKBgX52IOjes9hcLCfG0V
YKezmgRxGlMJB87SsVV6Cz3RST8qKFxRsbzX7q7pWokj1uboxqKQ5Vd3H1WHDlscgszlLRKKL2fQ
xizXJIOO1yKiCr0Yap/Z/cBdxHd5B7vAnNYZfhkh6FgS7dnis+6b8hJ+GRIClm/lzDHKNwRBG0qc
BKLzxksferRKkYP1HBvPD6LpKQwcesqsgMfXSMNajXvEkeIyRAS2/PvrwfbbNcDp5ZtA7xbzzQaX
afAqOWiEMvUS16MgRPbIAQx8QL7Bs0pDMIeGcJWgGAXYntsjlQHJWVnIyvPEB52DaJD4E7YQR+3R
yl3OyBWqX5fLRzE7SAn+mufCYdwFLdcKWi3NhBathKdi5b6BXSRJmHl3MbK+ox1HZ0vLWvYN6z27
euSks0nxwWBzlFZ2d2uNwU4V2E0zpVuNXNvcvaBTjR9/UWjG8L1dZV1sZs1JiNf4usMqC3nElJ7D
ws6jfYtZeRFWT1JCCHMfKmej1ROv6sjyXJBGk3zxIr+0sMOy3ylt3hkQP+2DBHvsw+05o4+R8UUX
bDwFjL2cvk6d+7nkbDuVCSyJP/W/zrRsa+8Osp3r49Tnwer18dj+rwBGhmd5KFmQfEkw9LGex7PK
AW4rYKu+27yi/NKuwakesiCRVTqwDMxfpXrHk/lMAt9+Q7wZ3tCgDA6HQzbNJ28grBFP0LGisqfG
OftuCUcde2VNrbnqWwj0WM+2TTONwssNJ6Uay+mabb2e9uQIe81ehdAwIX3fByyOM1wdm6ICAEyD
crVn9X/rT7GHVbORmSnA4MmlrHk2Rz6JKRhyG8KjZKR/fBV5h80slDxOUsgnnwm5koNH9CPRXfPU
WNSSNGB50PyIGeq7rLZTMilC6TwDq/F0cXV5GUwGQgXi74v+gLFYM0DTnRFF5JAlrcbxFrFTtk+d
9Wz8cRwtvNXjRoB1FvGzNld0/2I32JrWvLYJF2601LpAB647X00wyRr0wsZRiCT2ETwQlPlafwy1
XAD2qaqFeZ5ELm45OZxytHce9gdk/+HiaGbwfrm2/RqzHk9M9mXQRNJ6rXJFZlrUbczC5DHNfl+R
uA/jOblssc7EQrX7kaIlfktmctADIhsm+kCQhwPPAA+MINccDIIiAqWcxmRm6ru/LIcb0yiqveNw
rCzkf+s+bnox5A4/2wrqoEwQ6K3u2jmVC36o2kYq/BzXwDQM8shoFHV/pYFTnap/Sht/7tHXjpn5
8YYf6ruEjKaQlXuh9IRE054SqSUIAlzAFpjfvqYSFGDGibSLw/79cIbY8zBoeWGHyfBcG0WhDYJx
VGbDDchrx96lG6e4FnNwsOyri1EFyFCeJYeFjtdKTLhycPhCgmVu7ODPPnjGthJiuutX2OJLIX4G
Yd/tCVzn/sxollLq+EF0DLnksA3mf48ytLBL9ZkkNZinrKJoLjane+qDb98/q2jRPXYGgAIBBmQO
eiMfjfemQZvhL6AoGhk675sGW81FPY2zMdd3nyi7npAqd/cd0dMjCagpPK7+sNyJqAA2oh8JgPvB
xvBjVKPSiYiQWatM3XKYfmtO6bIHriS10yYtgb2YiQAnV4P6yyjaQ+/s79F1evHYJ1XGD8cbwTWN
84DbhgGS/Z9fdh1q8JgE+an+rauAoGjIc61y+mHPUP48jX6MXE2K1OUD5DtOTusK9JwBmjM7XL0o
dPOQAzDwFkdafV0QmxuxX30cwxlJIfAAk2x2+Oxd7lseVX4jF8hsczJtQO7QRHSvN6gqmmNiQybp
YZB/DVLbeV7M6s6gbbHUksgFLotD/XdxUojTBrlC9DnYiqvQVcfGT+Pz+zyzV0v3gXPy6p6pFaGi
c2O0ZV1SiSwVFK9ML1lv7UtaOKP07tesHodkax+WABT20ebF5iND0sMWPAVD5NcVtDyIclrMGPWC
gS/NmXIlitb6EQatN/vtscyqauAIgKolzRj2Gu5rQKmVx/9Ql8WwCe5YaDYk9PojwEd4TN1NHfxQ
fXfifvi+b871TAfeKh2ZwkjPrZGxXDcmKlcSo4N1U8eLP7PmYXYlj7Mzgour8jgZV8tYbYCXeFFc
M8hz3ymp8sqhZOWS5Dj9vP6E0zSzphlrlGe1IsR7VmruAb/HYmLMbFjQVuSh8NjJ3CyPL0tcIKKN
66DLoZkp+Kl1sHIgBmeZiN1ARCr9kSYEgDh9RIykCLba9j2HJ+COCxkG1BEj8P21J666Jy9KSYmV
Xl/ZfvsD3FzTqT6rS4JBZxH7Num6wWJHs6A/mfjnoaf4URH6BKAoNG0GXk8siJnx+MTUapQ1Ojea
BLZ772mD3UDZrJHv5/K9gVcs6LiQGBfJ8ZlkRRsPOd3vXVD+9BH5RhvJw7/TuMLUfTkyuYrU+6ga
u4c6dXV9+yvr6F+u3ltrsbW2mg1z6QNI7L3jUbXSdBCU+NJyi2P8T+VxkAHhjbH+uEtbSOIHC6F8
/2fEXRbHHVJjRRSRGwKVJJnp9WvNDyJjrul3F11e0wBuxiEpRM5O0EqY7nd+c+p8mImgCOK5Q5xq
FOxMejnSWREhKL8QbFptxdJnGNl0gEJz+/B5P0lsnQOCa21cH8JjGo7fjz0j6S/UlQ5FM7OJe6Yy
ceURTOdhDgsLaCHYYQqYB6jlTyd0ik/cWZQMha06dpBeWkue6GKiz2/zyP0aqypOCT4XhVZMiK71
BfquwnPOOJBxwSKW5vvyPk6JIqK/4YrLUvI3JlM9tQ8MI4q1nPwQZhuCH7+i45o/rpaeFdpb9W8U
H3tA5rrjezQuYXbA2UV7I2AKfMNeJCGR83R/ld2gg+rMNsYBQTEHBqo1wI7YLHRB+XqWPAPj1l3g
hmTpgWYdP+w1dagfLIHfXFRZu4JOC0TBDrZYMc+91221oTqhtppRyoso8vFUIIfHHvF6oPWKp4Bo
c3GQonjhCAdTzeOvhiwaMcN8z1GrJtEkARm8qDeKGZYN9pw968hIXJ5WYE9c3IO2aP17S8ShPP2S
nAuhdS/3szp/frmLd7M1HSZSvmizurd1Y9QI699oJkPGIpGV9jeRAM1Q+EyyXl06A7xi/BAY0R/u
dvJ34EGddd1vjtVuQQ9zAJJZKpdLHBNzAtKvLM4+iiuB24/yvjcEtCAHOb63oCdVdQIknxJh+Ip6
FRayAdRFZnxPxmKOCsY6E1jDHmYPBjo+MbrGuMcLsEoaclbrW9d85yyYhpG2MnV2hH1Pd543jZY7
bYDMI10lvwB47KTjYneSZgjOd4sC3fsHV09q5N/U9nJEqrr1g767JOnkr/KMP3UTiNhrBXGc9n8T
UZ9sf5kD4jyiBaVksZpTpnXFD4RPo0yVIXvB86v6NI7md5ycbuUfSfvHBz6goG51ezB3oKGl/Wly
cKziiSxNLuroxv1rUdjCgZQRwcPJc5XARIJPxthVAWXP20HpDJyK1hGMjKY2obMg6fPXucrbpk4Q
qK2MgKMj1b1397RurfFPCMAlk3aQr6kmL1OwGlM6lJ0gd5ibudSKaksAL4Ct60XCkQ6lvai6FVYJ
pA1W5Y3Rh1ku3dAe80GSpFwaF9iUgZ+Q1ddPC12HvXETypL2ztYeVpdvR7ObcUYtVzyDsjxt6K/S
TxHVBf1dXDd+X/nJiMiEb/3nBMvPZq8PErL7m+eiNu3uxJd+VCCVWKfnbwbQ//0KSCTlJ9vHhBmg
eXEdsp3TOUgPDVLW7heJWJTP9w6MuGBxeJUcWuxw//9q6YyB4aqaPhvCKoKW75BvZ1xbpcLd6skZ
UF+sF1Bb0M6x6siforI6c29aW3gIEU/MXxPuxr0rnYzHdUCXrZXPtbGb9udkLd7MDX5c0hkwWbek
phQEOAlI9xMVITCL8LTdE8qtAbLUzL3Wq4Ffr/Q6JXWJh27Ro6RM8qXPRkfR5bYDKGMp7CG4SCZW
hYIIjdeIP98SokSo9GRcBUjz9ZJMTZXK5QQsgJ2UdLT3Oj0ORdqhveqUcwsFze/U4skZGLpbzJGP
hdfYPCdPSOzGehe2J23EuWhf7ezAGLyXJW8Gh3qPKwChNCnbAwvYmjx0Vyb+C4yeUCaO1dh0vDbF
ENKwIRfpb4Ikwzfqzxt+nUrl1VHTKm1q9pwD2ReRd5m4D4aP2VtQDwYOOb5v+UhZTD70NX8R0Lk8
iq2exEm23rxWdejRVai2HX+fLPWyirYoxwfVueSWaOJrxYo2dXJs1ht/MAzxOr5edPwMvr4khtQV
jiedFVWCA6UZl5vZQiNfPpL3eDar+Y9BLTdtXGCqTdjss9xCfsWu+L/H4X49ZEoZJey3LwGzTaTt
2GYAOOlKW5RoY2In2Rq8u7f/9TkBOKVo97azeDyTpqrahOuYrGF6B+9F+G6ZmHlVbjp6Ts7eQb94
qpOmnK80b9Y5AOJh0O4koCqv0AtPXFMCTG3CtPobcvZN+Z88sCHR66/DkF4K7/oephPwMoTdC0kZ
tbqES8XZySCMXiYn++Rxum5ry3netcuN3sNvqD7wmyYheGe3Ujm2wWIc+lmJ/DBAgWBzXRlZKRfG
t1R3fAcDmyMRY8SW0pfI3cW0BzT7uxQYylMJhhP0GhQDGJb1GBGeOX83Sxs9aKe3X6QHRo8NCimr
6Rj2CIv43LC4x97rdlQ/woQsfwQmk6fwde4Ux92HQhl54prN2AwJhoY5RKWVi5YfqhF4nSDdeOzw
JHeMWh6eoQC7/PClJODiRTi2U3bD3LaeYYUaRIADMNg4j+1MVBZQeMuHfzozx1JXn5xXuy7kGJI/
/ogrYqSt9XGVzDFclrjAWyyjtKxhM0t2R/jyKVPU56vv20U+0xo5HaV4RNtk3stvcLzK28gBH7AY
1oZsdHBFyK7cZp1u8Xywvm10rH9qZsOxDYMdHl562+z2F56FnaG4LWFHSQwr0Uh5W2uSYyYz+KBF
iNI32vdO/FsrLYChle/Dad+Bgg1Z0Uje1st4eu3wz78o9Wkuez4yfMrnlp5Sju3riF/2KUjuwx+m
9reTLJFwVahinVdwp4W8nqZb8X1mqI3sycMRApJDI9G9fZ/BW1ewlSA0PamivOD8krQJiVba+P6A
iOaAc+8cDh7vL9YKckzYzHDn9KFcrtXoJLLzfE/e+A+9zmFsxoFAb39XvwGPc36zez6In0+tJnVq
CVdzxYsVDe3xVXAP8Bi0KRkLNELox34A3ZQw6JQb2x0o7QQAEk1ecmBkNhBSvBCxd2Mqs2g7R5yW
2jjtmozQPfICBXKgYe3YALwujZE9364qR+VT/Uk7OoJsdNba5lhplyPJBlhGk8DszymSewm+Hpsc
OmzdGYCFUBOr3yHxrhtj/8iOO11Tou4CQTDHoVkd/h827zN0xXtz94Bnd9Plgwff+kLWN89KBJQu
GRb5DxGpGvRdprR+hWwbxGUXd2L1AzcEGOssTFrYfuWWjZY4tBbhFt5pfCrbVExin9GlE3rAyd8C
hlC5ssIJJeavf3xiOCD++Ya7tsTgMcri+NX2u1Lw0ppKRCeIJMAH//0x82PjTa6GVmi/X+BSi+mc
yEGX0WBFmItnmB1XvrymenoaVQ6ghFQWX9X3gypAZe9jmUA9iLo5/lgQmZROmZg260zuV4j8dwxH
hspWO/vnHKNsRmRZzYNy5WIv2+qjSFUwAkIPTv4oxO+QPSFZyyivTbYxw18FyJFNW8U1uyznb26p
p6v5BTB0yreDkPTvZCNcnzaN9IRHhR7vGdinbC24a5JKoqT9+Vu/SOmwOzmAJR6qAR3MF+MEH9/Z
PTgfxhJti23ccv7ieAhvgQp/oacnuDw4xA56w0i9HBHiOKGlWb162QzMXxc5yedmsAePARYrakme
UHzfCBm5HwrZg4fSymXbvmApOnkJlK8oynkTCd1ygG3OE/urpvna8itXaDsKDXcp+yVv2imAcE4W
asw33LNCLl7ED6aHkOhVsD2t7J8R+e91pmpb7vI3GjYBBI7gPD1oI0H/D7mTKe/jnPjjirc18UXP
0+GeXJcDUSs/oYZvkLI5hrg30jJ91x3soHiIOwrMp63Co2NJFq71D9Jtu0lr9AkxWWhgG+7xhXkh
S8VOx1pN7LRQtCEZBTvBSVODUWvSvqftYaTyXDf7vuKmCN7Nb0TtGbYimHQZxm/9MT3wJsMwihdy
F6TErY9NAFurxk5Yv7zifc3JEhe+cNRq4wYXMKaGxrh8zfk3qalHdZ2m+cc9fbwhNYSQ/57ajePU
QrRPwdNaFxhkGPj42sgbmF9itc3EcXb69gEw0gHak6MxHcqz1dlqRvz84KeHTnyUE1CuMSlBh0wD
taxSh2zCEXOVNcrgIkIyuwA+woLPC2ryY6SotHzUrI5f81oyWmbwuNS5HC2E+GRqbWj6G9aoRWyu
HwS2DQRVoog14cPLaksquKOGNxRMIxSyN3AC1JLF1eiIwHmSDY8MI/mPYMznU6oG94jmSOp6GO+S
8y5DXGIQrrOMJPS9wbstwGX4RvTxIA7dtmhHmzJu8W3NYIxF4m0QUE5UEO+QP0aUbV4Lxo9CGUfK
LT8/2jJuxqNgtMG6/zfWOf4fbu0Bi7d0ozWiNeWNk2NYPxdVgLuiOanEpD2MqySBchSjIpyTdNct
9wkqrxBqyQucJHOMLwcgm6lHyNBi3Q3LjIbrmppYA1UBjK9yfLTU5XtX5aeafoauaLVVQFoK8eWt
NlwLBUorf0S5fbEobNOleZKXBuapmnhT4yTjWMM2o8jp2oD/iGHbezPlXSD8ZUmNkGFJR0d7kAAp
0h8iXC8q9X79Cr1z0O8dhCUqhqsEqUWvNAJt2y5MGP11nIT3Gp350iL8ERuUD7qQ20ul5kZ4EPRW
Puz9j9vQdu3rAvkN2jU/vMk533MeEwTBsaHnGF59o6CXrYf82DeRkgWUAH56wTzYEnshL5qCsHne
6txssjriob/YfKtC240owSgq8r3458VMxFEch/tB3rgG1P8HkENg2wjCsXAlGn4/6g4WkkIQN0wg
5CL3gGASrAaf9GN6Vc094egFTm3Z0MbMHjtzZp+r51mIrf7udTxmxkLuK1rTLBoj3juHYZm9olOk
wL/RRG22G/64Raph2ULXsdK2nvZ++azz2SFmMIsjAC8bxOUw3B6sjbAZyVSs4zp0/Ajmo/725Ldd
FsgIPoTzvLyHcM5mRPY1c5Qq04Rn6QKbt5ATE7GbbD2k0uwaK19SFmnnNY9vYV0whLOAhGIz7N4n
6UWo4Opz3+ZiauulhP3PYArgDtGPuHFDT+rFIwDmjYVuid/3n3llNQ3EVeLb4apTGEldkUoe9Zwn
twU7v58BBs5wkm6yNZBxs/CgO/D9C9hWqvhAmBRvsBL742X0lpgFVW8Or8mz2sMSfQHqmM/R2FV7
Xerqm/N1idxqRyR1TvEaPaBwZmEmBTTQ3qBi78z77IMdb4rx3D5kvcxb1QkXmB0NfH24zobeCHES
4nddWPVQ5LhSi9OTvSDxU/ZSWeDAmoHGovssUWZiB1wjJQ/YNmEYHIT/vhdFj//Q0qQMm+28kQBr
U8n0PKH0aR5Ezrp4SUvTPi8sf3ixkHJGtoB1mXb+nDNBrmi53lniAL7KJvebKpFDB0/KzFz5h9CL
qjcSGfBHS6ROVsE7pJk/hhNAGEcpnqnbcsk74MuEuvHEfJJXZ5v5GCaTnJZFSOoRGKJAfU9a6djX
9ixFtCTntLkxxkCUbXmWn42OA2kxMt0d57dQwowIBfF0BvvHKTGLS0z4PVC1r5U6H0MrAaUlMcL8
6Z0XznMkhqpC6XdqRxzMjijDO4ug6LpjJPkaET++8tIvFRH8XJojZvxBL12RJXabmAMfXzCTLiCC
zaNUcO1dnmW1W5tYnMSlxxUJtbuGq7BNI02epz2gvZYM5lUM/ffa9FhKXZFWjLs62p9ZwNVhm18f
kWtoWtx9QeM1YRd4rWj4C1IOhoWCqWa542qwJW+ouVcKglAYrRfA31H3YRWV4xH1ih/dCkD4WowK
gi47QZPOFmKzzvuLMoE8KQAmcFdAXid3nJdl7AbVCDxZKl8A3Acy582XDma2UPN7VZCLtc/2IauA
jIZOrWG5RyU4YNCwJFcBr1tsc2ajwK+7iZE11pnZU4ld8zJY7bCqbeHKFcWFKL9VsIzXaFdSM4tr
3zeJyoGSntRk5YLmXJSpLcQP+zZaRNbL9slEBUFEcuehNPxuA32GoO3sCQN9kRvbqfDm4HJyN4Rf
+5IvsipgO0Nf1iufolMD9cWy12pwxxbEsCTbNXqZVHkmQURBfoyAsx9DAY14VD0kONyw2zDnBQhX
fzVfhEoBk/O5734aazmvHmYkRXo/ojxCcrbeQ9O51Nk9tIjIfftTO2CVEtw0gSyrOtzijl2UUkM9
48hzeMAO+EZbgnU6cUYrzgLrSi32vdr7uLD4XIfhjZeojRitXxi7WlO8Ee96hLeEoe4u/MtLpIU/
uAzm4TP3Mrj4bJdrDoh/EHfZN45DyTbA8kzSu4airWyLx7jopawi9E+o3QVrtE9q87+TGzXRqZ3A
cwUD6C4zOlBOPw2+3lwbd2tqBoKjjZukXKR7dgixHB14NWcYVEzKEba/PbIXN3i2/SJfcOgpgj9S
EJSThXmzmpNvx1qAkHq8PvHtgZC6Co3ADhckD7/KNw7DbHPzC8PRwZfGrn4H4B+/Fc3nMZEpRtyF
bLVTpwpRVcz1nVwRI1uKfVsGEft8PhNFxBrrJCJj90qPreGivuo0wLA3JTF2vGmYGh//wTAftssD
0rOVkYEQPOFQrxPvSqQ4CcAzBLWp8GjxrFZh6MCJvAaDvz4pmqReNYHPkZ41PuPMD2cd3NuluYoL
VFymMCmZJhXl7QJlzaG7Vj5dfrrR7mKqWCmEsk0OcgxfMMn1CgMfCCTvUF5GonlF3C0t0SpBH5mk
K3JCaIdb4LFNMbDF5BUpmWVAH6PMY+bbUtNE1McCmiWhwhqeiwhSQyQpavh8nMaja/+OErGPqLLD
HPLIC8jNP4IjAbsM7Fwn411JiI4RbnSn6PG38tyqKiH0lXhh0KSoMbeTzG2lVMZnHwPlw3wu2TVx
SfDMljDrNkt5eOagruZFsi4vB66r9Mk7OouQTmKhMlFlt6+fBLNVjajLHYwbXbx6rxsr4sSxXBrK
CTvYjf/iULRpZpIvQdm7rWGvHjwGWvDS+JSw4rW/rMR2PEcR1Z+H4G70moR7n8MeIeYfIPPpYBh6
yEMd54lGrxzPIkSSUqcqnkJzMYetzpBgYxiDNNv0ZOsEO8lHg5R2TC6KDVnILdcPi9MmEy+en+CD
O13uRhVfgTvkL00nDY6kPupLoUAmTjqad54xg1xmfNQvLIkthm2/9jbSiGAyA6wajjcjTpaPVtTm
waw9EBkf6aZgw5RBBTpInlNGRDHq2L7KDmtynOmnV0VPlEmbectk5tfThiegWOyKhfezTz17o5TA
yY5aVxyq7MumB6qjbf5IoiZpW/5rPfmR8O7B/rbYs6n/PMlHf3tjylC5rb3vBwXK3R1TRuku8AXY
NOPfn4Zdgv2F5sBRLQQapy9VB8uf9yKeZXTsXfmH2GmUDkbrCW6FTlhyvbVZP8PjYlIOCDb+TKFG
E1ywZIKHW4DXQWg+VV4+Yi18GmGyHDF7zxJZ37bklVzod80RFMI9kyJlmc53CEZN8lJr1IBL5bo+
5G7drjFjnYpejYBYZsTQLGNx+HehwFKE69xofra4pKvjG3kVuWVVOZ75IyGDlq64ni3JXpVw1mnu
nr3txRR9CN9300EyUOW+ok8jYKuAQbqV4BZ51ydEITNaIO1QG5vv7v9oLnBBm7fznpVi1xxhYYZn
pA+kaK5U329xddpFCnJUuodT4Vskj4mB2CF6GvAIc/7zswpS0UGnBnY01kBZljT+AF03DUcTP8vu
sE83HHmFQYptwuQz+U5dPMWuw/PMzWYVcTm8MXPdOu+XagNnn9F55lMVamAkAOVtRY0n5OGqpJPj
zLY3RYaiP/JkCvoaKysBkw7Iqi8vfwt9kyvqDsXL3XecDID6wn/OXlEfDO7CPoY9BMEBKQ62luqZ
gY+SBy50usBqersGZV29e/NxGQFO2cggHQYVjdnyCuH0ndIfbuZirvNO9F+/v0aJdFPth5QlQ3W3
14+/R0iletwcEqTfrHsKi+AZSiJN/ZtRj1hhsNJHQMgmgYwpEDSWNX40+YRHNoP0zBRXLurmlLLR
/RI01v9nIx2/ZK0Hv1ASh8KiGCxQ+mZHpSJ4ayvD9FxAW09Zap+IZgN3fnCtQNc4x2EoBbekSVWZ
gvXzlFaa2iU3vj5OjRSNApIvbZSJtBfOc6k2eWJ30BNjjwgyArAlwfkQxWzemI9buQTrIMZX6134
rEAmH7Q3fae13t7NKKxoXLZd3sHcuClrINp41tM7CD14w9+mAdiXu3mdOodcn4PbnGf8oPq2QmR6
cvJFDxd8zVvXBpRj9T7Ejoe/71m533trh1DU/7aD9lLH7hT5r1DQ5a1DZLV88YjFUN4PaxJ8UV8A
iOQ3lMSZnkfr2YRWoWjW3YZzQA/MXFMYoqSKI5vACjVFIV2mSbIcl/k+YXEUd7HgjO9LOFrbwhXn
R7BTYGDmwGAwrV9JseTzAxSGTp6b03/3WGaOOZtKw5TnxZ7+LyLt93eK8unXYi7PwgQcZ6bIwPhq
4VZos6ELWUrEDcVmRsLejTRcCBOdM5gE0dj3qv5mV3MzvylsHvxvfIRIEMSsBtMx+oP/eRgNHTA8
vqC2SrHiW/As1RypPc5+98bmMpunNoB08ng82Is5AvjR1/hYIVjcLqLBCExoSmqJkvkrBCbvhu2H
ecmNGlRcJeRfG40BRyIGktUwERUG3jIccAJ6qWHyr47re3m9obagQoBPzY10tG1UIcbU3xOMmELa
7OBqGbCl/rEmz/9kbA6FelWMvMb3NmYLylnPIGXQTNrTvd9YQqY32allQGc+ishbyfAJOm54rEs3
QiIxVwa6Zc6SGGhz9Jk6Zp6PFUmuEkYGMGZf7gkv4xFWoLjnkPR28S1kCPLt1+6lIVjyYAELsb1x
QzLxFvy3l5kT5OfkwI71v3596Ls6qrZrZNfeKLSKIQ5zIL7aLzPKKsSpTdIsvdk1Qh+F1XQNRymX
bCtS/wrj5dcEkMr4OZU8mOD5vont34n52J1UKT5NAziN/F0fDFg6BmEuoehRB2cHz3VaS1S2w0Zx
lHlXV6MJfGvMBTXceU7MnB/cs2TjCyeuKv1EfBZIUzkuL+35+G6WWkdAPnUHMPoTPnip21yxPi7j
39hiIyaRA/3S9M0Q7UzVJ6/voJ0eIpQTY1T1wos4MQbYjfwFVl9VcWJdL3Jvq+o2bk2trDKdAM/1
J0y+IvnSPeeg51r7Dj8nCmlcCKBRnP1sKUbTsgX63OcBU3ARiG8/KWOZiFIhk23KtoA3LIfDhxIP
eYqp8ZhrCkxVZbls+VCeeiktMQZ+vXvtz/1zobQ4gLYQ/ZQTidXGGY4xi9WnR8K513SAhbGZ9KJd
6P0HRB1AOqXdWP3Z58yeHT6t0E/Q+WbRaiYiJlx7Nf8WkL5xCJwnIt2Do5q4DeQooQauvWfrZbwg
7shtu1mmuSq6f9Acp+yWNq7/jm4kXOYRyUDTT420a57ibAtTxvIM/Y2D0yfkq+dgnx2KEwA0H9z4
wlKN7bOBA0th/u3B+FWpTbABj6NLUIOcvRewVHmLHwMaKPQJKR3ShNEnvPm9gtHmx3iMNk7qKMbV
VWrEJhXdsnay6ItnysZGtodEZovPmp31lXlWfae9aYBgFhvRUYdyX1N58EfSdn0gBVGdkKetIOPm
19guxC533A4d7hKnYs+1ru6A3d1HtoRgYMrvahHo4PDQAwVvwsRXa5xQYjSV3w4dmNAIKCEBvxxo
TeckkymWBReIOq1mEY0pkwJRh3HKaiUFir7SxfJq+ABT/rvCnFtIH+iAStZ03GyI3cmqf5yHgkJi
xgAJdQfFbCjsQCbPhPm22YeQhG1VKO230J+JIYCOtDsBHzKrEqSiHVFeGRbnc1oqXv52AUmEM7Jx
zEudSvvZqueIphh88eW3M9QODAdp6brroAfRwtQbJgRVcpsuEX+z4rTMVKeTCPlztE3T4lvvttTj
qPIQ46BFMUhsHNVHPRzZ/tefntE46c7tQWn4oRWPPfB9ZToQqA+HYWGVFNy/RHpdQGHd43VXpYm7
dshWm5JM/tI9BweCjgJ9GKyMOPRKa+e6WJuUJKG74d7h72t3kfHi4IpM0ptmkJ51si/M23vwhQFV
natlt8SOGLPiHyOEP8GzTe5EEdivu0LDM8rxAiMHn7adqXYJGYX4IpgXCME7jMP5JfoS7Bj5ueoN
K0Ujl/FHNvsrqPXOkGyzgKOierSxh25cI0gU2OrksnmO4pIFJPrQJfprTaqmgLNH4EXqymzlE5OQ
dFqVFvCTeWMQen10McjKDqlKWV0WxX1sRnQ0WpYov/0k7vshXtZyjWS9MF/1T1U5N8vaCM6De1/T
f7Icdr+cl05kDC/c5dzKblRFiZ1cr5AC6dG7inS8uSXdiJdfITpv/GUPyYS06bdEhWLpFj+ViGa+
hn1+Njb2O7jRlRgIB0wyj5umIRIgm0U8Zi+8CFztShB5QAb5aAn0OyXruH4mcpp4/H8VBGapgqyg
IJE6OcNXAI55fUqGJRqXT3JtM2YUxCtga+uwJQ9xmQ+CC3XPNF3D/UTxtks9sxoljvsz/+YuDLM9
mfvp5M0Db+m5TKYcGGxHjI8OVWxW/CmeCqQUGTb/p9T8+2HU9TOmiRBGj2XX/ZsSv5FZMzjBVazS
+p+oWIBoPAWLV6ayO41T2BlRlOz8zMwcMqWCbnxq3rStpZUdoh+U5XoN6onRwwoqsdnvWmKXPkMg
LnjXZKgdlgNFwhb6e2jtck04NdArxQ49is4CocxoyQI2lg8rvOeTvGU8TWLHTfxAg4gYMRCvzYcz
uOAyuZxWiA3aRJ8wq2tFXA5QvMuijJ7fKhPFHCO1VBjYv+n8Py0HrnaPlRdIZOZFJyGwRu8qNYyy
M+HdVkKZvEb5xmQYB3dzNFHCMuM0LjZjYUT2agssrqpXEqBLC6Nb3FkoAYJfZiMJuAjKcoL3fNWv
97PQneS1h/iwrf4HzX7uqATh7qzfeaWyO70mSXA27A/ytkHX9jm7BuzPaeKukn/imzw/ldBrnCWO
fzTFhe9F6FbUteLjKTxaQ3v1jbN+dL1f9uj/qMHadKF0kpQSlMv4t+k3WEZHJayJrzKu3BVmkkLR
6MiznTCU71XPwv35H9BiEW463UbBuKwoDM09ZHxMqV9gSFe6LtNrRHzqWYRzbzHkvezIXB7m6ut6
FdmIsi0rT9JX+7OI1ZFzcoAhHkO8X2gQ/j2+8meI72VMeVcnOOpcoCFFQemE9JdjlVCQopfzVMmh
oI/ADSsDX44nPoZxL0D/HGKIHwB26qNJJzkCl99hT9BzB75vRULqJw0V7ZzV75YtM3QViwKWjNaZ
kPiI2X8D7BR8EI8uzjBNMFpa5h88gm1Gtp44M0h/JJIjOwMKjJLHxJWA+sDb5dmTyJkJR0kPZkfn
pOEYg1Igvvhvnj+BtqAlE9F0pB75ol1JQ970wkSP6uR0gX6W2x0erFp2hJxDD0ezvwd4LcHixMLx
gfyi3/ndONuzedEISOgqsnWvx2zxfH4wY+1AbkbOyh+PSrENH2TqlGGXljmG1o1DoRTWz+g0c1vi
5QZ2dh5a6MZJNOPysWMLJ/YhohqgCP+Y0cLJMarLmrqatTSOASj27VAa/CctDDGCDq1JGHCrh29b
ouVBw/76jZbygQz1VcNg4DlDeaLTKFKx5JK6tT607CPaZ0xAtd/SJfCgRcLvJSDEI5GnvEELgINc
78hBKP6ea7Doa1THMPjoBlqE6ihrRbf4e9XZIoLwRkPt0XMl4qIlP7inpRdT0zHnVgFaAS7OgQt7
ZFU6Met0No7jyQl4qbVl3Wp/067gTTOJGnM2EBedQq3LT3a4GUviGZlbQ6DkEVLn9IsNTxWLDzPo
EhvHhkyFaS+OdBoRzmDjZzdI8VIz23w3sEEaQmJW1NEVtOTwr726eSUughQ+MX7EWvcf10W+QR0s
jStFmbZPOPXmY2Zk2RmAABCkK1DKPXQxDS2OLCXjpzZyyNh6oOPrUWnypAF/G8TkAVQJTvM4j6xm
i4JCuPoT3y6BHIjW+AtaYwm7sGJJPuKjqe+3N0AtM4Z0odIm92jXXWdo4Fn2cQnWY02dnBDu36uE
bxadNXnSKWKl5P2zoZ++QeS0qi7+RV4+z0BE/fmFwtnW8htG2SwsysQvJCI5HEBVpFVCw/XszHT7
mYb3HJokdfFbutsXkQrbv2SvWjbyfbiFo9oCIu2tC/7gaOtKfXQ6aXbX8epioCF2aR5piJU0EEDE
sByxt5D6Qm/Fd0nXg/iq9+ZpW6hHIzqTruC0f+UybnOvy+kZdcBAU9cgHu1nk3bQOD5FGhZdEhDf
LzBHHcUIovewEFhlYpI5amKSuBrAQ+obZdPw803PPwWnQVU/sZnlFmphpXVsGZsuuaxLxJXxd4hT
o318H/BKs0ltcIAPpRKXMyaDErcN4CjUlaCfUViL8wI+1QakpPFLvURvJiTkH03LZTRsijboBq4a
Qu0jaLBiZyfA4qlzs7rc22XrtjvYgSyciS7aqndmER3w0/sW6I94tGYv841mHOD//bQwJgeeSB1a
UgPFIdzkFz4pokq/SXFg206ZebfuLPb4/d6z+y+Uww0Z2xlhsyx4harO4hRIzbmEofAaqlFc3nkn
LORemf2HDBep2qdJqEu9DQl/BPsiK8TyCpNqLt9hqHBA7vjK/j3428A8gC8SPE5I6qAGuLrWJM0A
XFbhe5OyOn0KntosxaofrM9d2pm1wXS387sptyzMusuw8uK884NRhivcN9jWUgEEUPtNwh8ChCTC
zH5wegiCJ+6ve4E7moBM8q7TSqwR3ZVPW2BUSjzU+GEpah+4JTq2rKjsaBiabGDShVHBVYs2g6XD
Ey2MYJ+dLVivudHQsaE3aoCxagU0sAw57qeO0g2HMhFSjUMuY+lNNeSN1+YHIM5fGlcpAW6Bkom1
4qJEBd7LCNaFyj3GBTrk93wNY07tTL+nqOgj8FAKWn79UV/Byx9HyxyHM8Aa6Cbbmyx52I+bg6yH
H9NHM8itfuYb0NxlHLKH8R0O99KWOiPYVQXojOnewy348LEHzBIORfFgIOr4A6I9MeQzVxVfBYLC
2SLzvxh7SGsOSJfwTNUqnZzL1x/DgKxkhkZ8qJEnjUS/MpOHSmxL425BdaojQ602SrAURb3gUtVR
YJzFxIRFY6KgnfNI9daEnXwqiIK69Gbl7jF2lWps7tCNDZWZI5bnw31LxITMB0UYJ92hetkdiTC4
4mzVTSsSqTKGvBHf19QfSs1EjC5qRqqeE+aCXvHKWEmijdBClJenC6vvwpJkL9h6R17IoGW0vZ+o
ITpVyQcvaeFUi0hxs5llQ0JwcXDsLuXnti+yEnd6wcp9aVVqGeToiosADruOI5zdAOQfPeU/8LFp
W6uSbVOwC2kqfGspsn6Gt4ACMzLLEa/OcNdnbgnIeHE+bGCTdwAdgyYSSTp3EL3DnfcJFZ1nCCO7
GC6BZDwIXXeh2O/dgiPEJoOczS6OJ+6z579jhUtqTjbdFodVaRi4bHWNlWf913cJTj548R7XlOeU
sSBgJZZ8S2/BIhS6mIK2l374UpbbVLJHSSyx6GVZK0WtVzPM/yCy1UPA0NAgUCpqd7ysR/5qJSJz
vWh091AMcG7W+A9NyfSmm6i3oTyqLi3OYb+u2lO+qTqpRNqWW4v2T+KBoYypXYDD1o28B1UFlSkU
sQJsezn9AdHRAILiaABRk5zq+zhguI5fUwpqKtWZve5v6keaRet4AGoqXR/OB601b7ERIpueF/9R
i4/ULMn6bI64wmc+5gVBNVpLWWpWmmS+pxUn98IdzrNV3+AA9m+hPL+pJmtNG127TMP3cDQvBZwX
ZEV2xs5nBcWvrAsnpfpuRuru09TTbZEcCsueN7e0kGyFoC2K5JtxkQiYK7dpPhiTrat0pIc4+iVy
2/VmO9DrkAV8NfCa60/DPGxp78YRRWmbrEDsBHmQQQYPMhln8Sh7p5QWu3XrcPABfKFFQxR/pfe+
U/pzA/GB3M1V/069YHuPrBNHWVU9/rjibc1SV+1y8OfCvTqqQsWcKfM6Wqd8B5RujeDu1vBIPcKv
/zpnyakG2hUpope5A7J5SK80Shc/7hPU+fB7sZZW22kXGLo/fBcUyOJBX6CuzapE88++UqnqrGj9
BXlLxmjxBkoLeC9xX7CHSC0+IZWhfgFByszhT4z3rw1NU1B8xWW8AKDFNnAnSLUtWT2X5OTtovJM
O0QBo8H8iDgYaZUAVng7rxchyqfKvXCZa3KujvP0MVI74POjM2a+pvSo5amOOYjdDwxkvBg5a5MR
ML25ROvWMHKtts5WtxT6Q3DG/vmcCUKJgcEKBwrJUIBIEm70HRrtzsiHYDrDvLO7Q/7/2q0WQtEe
WCxgS5HdDyeWKEluvUBNBq2D0Vf1ll6GJclAWfyzEUxvVJ82BPBhRwiYep+QTkIsstfDHJMzzlVQ
Q0FItK4fak1OBmxkNt4n3jL4bpW1iJfVCL089/j6nqaCy46zpRHYKq0tXc2DRNG3X9+1fU7hEJqB
5XMn0xY5DFAvRtk/3yuGlC23yHGDzBdngfGMnp5OBljneal9G7ncuIW3NmcEvH6RG2q6SgIFx7jj
MlbfR+KNxhmNc0aH+FxlYytgY6L3LtTQ4iPi0uqPPGD42Qcxpqv9j6R2SkZP0UZzRQxx+KRBzNnr
bAlsrhc3khjMs+SVlgrbcwnugzKlx+jyIzHXhSFhWhpDbgmsAlb0+APKhmSeaSsqXRUG5eHqO2EZ
gRLWzo+cj+9oVaK8YJvVS6RCJW1JZ4k4oSOZOnn9dYzI3BXEdKne0xtbqUbg7TP4JbjVBZpysRBq
afzIc27Zu/wcMWeBoP6/aHuor7jqzK8DeOsg2YRNGAStk5uCb/PaLEyPUkV0+i/6LeS4sB0wHLro
26AIUF+TKwqw9+sf96L9Fyp2lheHuSRDYQibktohFe9YZdDNI2WlI11ONNAsH7U8CoGMymQ0UCa0
wOPgxbj4BZeUb8XXJiYVhOGZcrGVpIusA+l/meXnTS3Co1zlArUVxIQZD/QuncSIYNR1Iik65s2S
FHFA1EAF57aMZ/Tra8WqM5sIJw6Em7gt+ViW1BHBs6gonhfEwrEpRRX/LRqJEZMjpz2FX8q6YMet
E6BfL+GVYvN010wWMEcwCrhreedftEKajEQkffeYn5ATEmg82ysNIWRB0RaJ9grQhWx43SVOvJBp
11r3pfIpejHX+8Fm8okJtvYQDGy6Vk/ZS+8OSqzMZAF6TLZiip8bi4CpmykVuDbtAc0XWXG/uk5k
RQVPRTO3MaH8clwJf63ZHx/kUCT+IsHFshq+tg2QzM9lboqFKbhG4qHASL5i7xN5/Eh7rwCmv52I
Cj56dFSrAa2aYRqnyUMnD/1gt+yX6caRT2b8byKFttqhNZRbxJHsuWHD09+MecClB+36k+aK6AZ2
rpUl3NgwxQwaebZl4tk82yR6aX/pA2V2PCYRofUBt0fgktpQ/xCQM2irrauiR5iVLSQ6VLDwBuHu
XrXHQF4rObC8rmCbAg62SfH3GSgn0XhbxkP7gXaHhTAWqG0a/XYU3wsapQf6LynTHI+hVUkFL/dg
N3oWm9aWXU6v9fHOfTOxO8xgj1nGXbJ8kdmj80pKma2xLjVqXH6GuZh/sOfiloIYGDotDoIM2MHI
vAehMiQsgupo4kZynbIf7VXFlohJC/bUwL1/9anpgykS7orbqoGNDS7IQg9+7DDCmbUYUspf6ECP
5pVlO7+R9RvYDrhxx/7xxjumK4nfU87WtMGRGIdleGDw29cTiI0WE2PwDiNXKpvb+EjUqdmwcLdL
/buHGVcaQtwLMsDW89bjZcEOU7oMtQRkXN6Obc5wnbpZjpEdPliI6epw9J68nF8R6XkTIzT8Gtq7
RZSt3gphflwsJ5dOn/y8YqNCsnC5KmEVzlc6VZXciLGwtfZCBLJA1HXsT3F48VHxhk3Wses6GQ2g
cKiDY/OXXrb9xmgDIasAkM/62EV1gifXFzze6yFtjVmh0ud2t7TFQe/aBjogOXwzMInkKTL1wm31
gKQR6F5Owjw9EHNCcql/4eAjOo2z2wnkNF+W/iIgLI+1UmP3WJgYxdfXPSzmfo31Ny0W4VYFCNXo
D1J2pQFSfyOKGFVCCMJS1fdHthmru0PaJwQumyfkzFN1lq0CbzIY7S+4G16WAlPAoedM1W54e5OC
QqXnDBzcbsDj3e/HkLlxtzACdf46zmyso3RBjRuHrxnozJCkO9micvyHCP0ILip/3B+LyCJ+YJuw
lFqdKaMy9y2t1rwUePNcTaxhGo05bqvULBZUWCi01O7/8l7SssAM5QfrIyzjUnV/lJCkIYueTxSg
hCXyx5TXbv3IRDEa74tjY3g8BRs49jAih7wkrLoy8YiYzRguEnlyiSr/zDv++pig3r0Z9frjNYEQ
6kd44TeeGpwLr34ZZeoiL/EhuSOwh+Vu2DkkJr+JBeyEsFxYnXxQCgtwOnDzAJfEO8wBd8Zjqjaw
rz+O9Ehmqdnr7bKlDkFVguhvkA+3Klmy8CJwL0HEloKm+bcUxQHjJFqXcIMZoq9+ZzyP/v+jtOTA
HJQuGISqG2jMtCyM5+DwKVj102vcVAPa394da1J7QdvBI7Wc6CsjKxZlcrKw8KJ4UWnYkhOvktKN
PSal3aUpI8qSL4CdT8vRs0wY78vVOKy03znvdgZRAcyaKdmc1aOcNqzFDLa8Vr0EAxn+uZvgdxw1
LcD59asnjyiAd23Vvj7DOcBErRxZukd6G3G+Saq8sPpW9Z9CQGntu9NmqWjaEfkgPo9ANgJxMcl/
792M8w4BSn9d/LRLIqwFvprksPMpAAyLKafcqJBotAT+dCQkCH01z42A5h74yelDb1PSPve0UIQn
x9OqB7hnMSnTOAU1kXwJqxPd1Z86+YCl1aIFKTCswAyE6J9EpBTwVdTNJzJMgbld/ff70M2FwAu8
HrPU9giknphSJpAzNuUkPagTjFFfigS2IBDCNJWSQzs1FvTHzCeSz/JbGVq2UCng9J2e59Y9sTal
vHInxacLz9LDjLzcMGd/jvKGdW5I/CiR0GfVCI+ElS5+GhfhSnAFc0NO5gKmoNMimyhmmOcO+8bN
0F56HFRhah/NLPtPizC73pediUmkwwnkgeGulORxFXQkU+67Rc4UxVvXVlNgHAIflkVitYdbq1v8
nGQh0bns9tRWOnxSJPtdAqRwGur1bIATqJHHhRI8AuvTiUeFFHVHfdvBmlIQQ6VVP5aHAhV7pnhR
3a8+GJIL0hIP2odlBt7+oaPNKqPf3fAtjJRF3FAPxCHrM+ZiJ7V77BiqflCLq17MWOKaeoQAu+cq
EL86HJTp9P/aUKCJKLTX/B7xpjMav4nGhkMSDNNiqsRWnKTNlbe2+3m6QTaDx10vMyQC67MgGOpa
Oq+CtM+8Z9rJtyMtgHChKxXOTPxyrUV3TU3Zd20BAMpwfVDJZ75ZhBnL05e3ussMkGD2e1MXO5U8
yWFS2LlGr5nr51EVz6/Fjl+MVx1HiL5HGZiWrXXTtco09Y6IcouJKuspkFMw1MxUyeL9D/MmZl9B
xAcamNDCqygY33sZB1BWtjFJSUjkS3RBcO3WUQpdI8881Ep54bKvfBXDB9EE+RUHT6pBHdjUI/J8
wWlhm/NErAr51bIo1sG7kXjiL02ZMa7X5Ad2b1XMUvhDKVlv0qZwytCDVU6cWguArDke1OpT+dJx
ze3s1AyHTBR0V9q0vUCak0N5McGh2qXj1gd2h+9D1Dy+8Y5FoJYqFofCjLD0EkSv+Wnq5Uy5ULXo
TLHxULMHkb9/MIENCUNq22qxjNo34c66vDrDWPiPMmuLFQO0dRUSRtkAIi+Bu6weDV+tJUq2kJ+J
ITByi92mOAtL1MeXOhahpbHLjdy/ONV7zkK7FO6QfW6aObPGZ/Yty2kMYlN/Hdm+BolDGUKdxAI4
SV12QHrpSoqKPKbmeqk+kl7RGtOXveDBKZEGeIYUugDh3KfUc0c9Z0FQTJ905Ynt/YptYlTvxJH/
QghJ6jHLww5Bdlpm9XSTtTraXpu8vrdIuVMvVlvT/XL/IwEq944aSR1T51PGh9ZVprNeMzQeptaT
hmCUcnyagNDi9m2qAF3aJsIG05t7GXFSXe9JKO5+PvCAOnTRRBDbZicRm/2svsU+Yy5D0XyvxFLi
kI1BzLumG7wDJZC6ByxSAjwvlh5SoKXSJjMzh/wIDLmSgu9+k6owhT7b+Be93pH9eO4lAldSfJ17
9l+5vncoYgVw8R1f63t5iryBaSv12qts+M0TTY15xNJNqtWtwu4A7PZiEgTfyzo/IgSgFQgfCWPu
quyqdFM+FTM7Jt/+wXnCIIY4PoT/Pyl0O+OEpAChmSe2pa8Iic+n45m+NNKNokXSdv9xXkcfr/Bg
IRQnBu7xCtbsMLl6Isc6iivQZVNbcvsvsdUc0rGQM5sbfYJVi/+nD/FLYW4lISNM6nc8HkY5Bb94
jR6KmCphnwUJsVewym8D4XTnTgdkjUN7VDOWRiafWSyjnyvAXTRXPkLWnQeYGEkbwVAFUcqy8jMr
TrvNhVP2Rc9vu7M1sbvsmyIniwRWZ4zq0bRhLXAloVmBwb92iTLYBjwtxto+2qd1YX3Ndtb7FvHx
9e0dEq+Xgb4k/zxeVfhZm+PPoyA+95B9Ml4ElDnw6o+hs+EiKznVg7DbF4ZlbF5id5DsqtfHVtO4
+4DGgwVkEf8Kgu2yr8HVP7tE9HcGwtCk7DsbYJHRZ7hERsmZs+NyFubtV4DRoNipd+TXlSQGirNw
69mZe7koETLNv4hUQIVjlrjLeFX1kPyyZ+yHS99O9lLqdq3t7TqVechmwJjTVfhsOsYNM8IIXm+Q
x0dkEUhv81Y2AsLuw8BDhS5y72niS466s7yb9+5iW/Tk6O7E4CSgchvP3nS86zdscajNWPQ8/lxg
mmVSpSuVMNLp36LtRLr4taslGScc1YFMJXg8+txWd4aMQROorJ4T8s9rYS6zQ3aCATp+npY0d533
emLe+qB54sp8Hb+4Dit3jaBObPWOkQYZqp/iozbUSx4PJWsCfQdJMxox/c2Z0CfgSR3A/+gDmhcG
sku1bbK7jMyI6VMiFlMDoNiNTXTIS92+EGWIHIx1JuraJTP6rN8K0VBeXO7+Fe0DcQE5k9LRh8OT
ZXJ1HrgtlRyVgjlElLspjuol/ljfRYiyqjyhs63w4xDzZEn/9nrhWpaX6PbLQfuSpYVfW4Jqupxb
JApXGG7qAm9ZyEXBbOT8crqDpeUVpPsLfuCDPJawm9aWdA+M8QyMH81gq14umDJfHZ2Rnqy4/dzg
eikqQcXRcSeuyfYMVgyejIeOursoKlBTaswUKbUoLu9x2gEN06WKluyEckgHxZjHvV5zMocgPXDn
/oYugaQCuyjBG9XLZ45RjNheBpZdxa62+sYGe6Xl3k8lwd8BLxBkH74lyVf37m1vdn+gO3yKi7jD
i1IPUN7R4EDsKOX3q+PXD4ew/0RPBsQ5Vt2qC9q02Ir4sxBx6ySUU3fk6wMW4NunlTy3KV+WPFVp
ypG9Dxpm3ajygtupJ3no7L86rXkz74Hyxci57GUAAdBKHAXuuC2Mt47r4zLVnR+0gyPoDipLaVRs
wOh3gW3akXHciZObRhNRoubM193aEKYiWOXJS8VMFqy8peWG3fNVpv3gxGskEI0MGafA6Y1yrPbt
dbgDcG6hUySwZaNFZCjEw0pHegYWN9YAb+N6yW+UVb8cHCN4dHYhaIp1Q5VG/tENuPBfYAJQ2eE3
5K3iNC6TztZ8NBKKjwmRFFk3ykvUOeJrQmhqHC+hPSrG+ThAFAn9GUx/J3aP2dRHqdiryAm0PaFW
SC4zf3nDrlgqo1nX92JM3aDnVyoTNKslgD0ydAi79S5n/OsdEYuctfwAr4uFSmNxGHNwvOeKMOha
Zedu/JAaWVbefWWvpKzYpGW4vXQAXUvDT9PDToz9zYEyXSSstF2s7/DCaxM5XasZVaqjVwbymeLv
QijuHgDF7Nux6CowAelDWdJBfIg+kOHqpqfo+oNnILWnIjMzvyjXMCUmvP/j4nRRZSZaQsPNYrta
x3tzVjvDjhmGIff2meF6DBLI6nCGDa2pqBhQLGTbbRQocqonXcYx3qDiycxorTUtTiyJtxBKJGOh
PcqAOCF65lGMVy9UwLeXbFHfYUbIeZaMR8jUVdKWGaefcNuybGumqDzgvrSmkuAGw824RTvWfQ9B
tH2E3UQN6eSQo1xc+aPL7sGm8FW9OQFVarQGYrxA0xrCzJYwB5MpXouux+DFcMBcrVxxWZKx5bF9
t0T+9jX6oBf8HERZbeEptIGhLccKtRo8hWnbOcCqisd/7tYrgo4jArjQqq43AsL2eBvNj9Wh+Jth
IoXtv+yRICKx/q7lpcTyifaAERZU4QPszRAPMSSj0yqZoCTj7/kEF3+23hDMtRUcn9I5W5+0F1Zo
kZp1GPSozcZ0ybbiZQj+8Z+/MxrV8x7fxVcDyFYuk/eYNDXUlxPI+URDWfokEkHdfpo5yaZrA8BL
fgB/iG+lRqy89V4X6FqhMyK6ggqQ2TG5Fpcme12RaF0Y/1SsEQFQ2mEIYBU0duNP12PRWs3SyVs+
W6j4yve8lh6vFoVii9TGldxw7dDWZxemPUXr9o1Oe+KqpwqVE6JufJQ/WFzwcC7CjmkmcvbSBeua
tDkjz0hIgruGiqejKL2Ww12yLkxvQZgsw9I058PTxUehFzr0VYNr718Ey9aLDpuNVqOF0n6t0BGn
Jlq2ef2CzUQiFR/pvTQQMggXQHvKALXxC2SwbY7dd98L/pGcD/y28bXEx8FmUz2TzUf+z+UO81sp
paorn7Ez3rMjzHn1CnvvXDoPqDXK1Nobr1oOMHB9/RUfh7N95QoCr16FA1sVrPHgAJzNUNgyApFn
xw3TTRCtmrMs8TedpLAUuibds86OkPn1YoyNe12qKsdCL/exW2CeUgHRDjTcRyeYjzsm7GWvTUD/
TMwYxGFVbukeZK3jJlELovd6kMPNQgd6GrRRyMktO8pbv0C5hvSz5Zfx+3mUU+txV2P6Lm+bo5j0
amkjAfeUzLY3rM8D474t6zWrS+VX3XNuyqs9OC7niQwlvSULS8AtlptIH8zi9zrpYXOpU+9q+hvn
aDl1Xx26d26TNGxflmSdbej3ZHRHLw/Whlsvro/kKu3CqGYcWmrDpK/xDo/tvWHc2zTpaqpCTBXy
fhClhlYeHnmlMB1mRMpHEVYWlLGEO2JXb23og9+JAUyetzJ2BTC7PcIRZjNXuFrB4o4hFsGALdjT
CZt59HksiMMOeSk8vO+oScKUMEPMoP4d8N4Vy4N1lLgVaVPdUYehaJnRBfHBS5qAnOkN/NR8SS6H
W4rdZMmbkxMypra8DNNcoX0JlZfeBFzHjuEWRHApqakklu5ttl4GIPCqkkPHQCiXIzAx8MTexh0q
uS5KRHxH5OwqRIc04ve2dnqLHLYykONY67wMIm+sHhfAE14s6NuH/NIeEhkdGArfABFSCuQeOIct
7lRRkDzhBdPb5vVZdqZfE558TI+aUIo9ZKcfLnVzpGiOqbr3WlbRel4/C1MV8n0sHiw3eHUE8H2S
sVCyxKmXhYAhHhFeYOoZ+nkMgkbMmDxwMtbbBuy9tPoR7wWOu4XOwOtHrGUfqsCV+vGPw72HGL63
9lKJgiltNhjLNr5T/kstNs6XDWx2kQIRsfsxVZSYqaQYE3mv1Lq9m/yYa5pK1/067Segvia6QNhX
fX75GdGOlK7vrES5lkhTjy6j+DGyM7hfQ2CIHH+SAbGjcHmSwa/kVvVB3cSpAlXUL1zFjSEY5joG
G3jhXCjC+fDPj436PBd2AYqCU+uIWNvOFUkMQzFHdF+VxDCA/4p1/e1EQ8+ddxqc25mPlBEwIRZC
hBhkf/NqrVyzsFF8Qp+KpsEtkKdOBGx58x5utTiyawKsCU/nNgn5lJ/mbq8QtY1Hg18uKeLsBRgc
1y4AAsCR8xVLapKGrtc+yajUdPDdkkscLRUfnagN4uAF5r0zYhrotcf2oGdfK50owQXHAifT5GzL
6GyzpxwoxUgzZxPrDT1JZQ6TwW+YtttDqVCXcRrl3IOXRkaI5IWA1oOjTfF34F4S34zm42aNwHfU
iSGhepZYpZp7C+LtDIKL2AcbK/oAp7ame5Ca+ZY/kawqyd/n48jQB73eEA4CdYS9oiaFQNkuk30w
WCifCGl45LpW6teNHm3S2vWwTVMbX/o0SAFX/5F8NUBuE74QixCBuG5kcdyX9foU8Gm7YHyFZwZZ
yXbJUq5SI/Y2lAKuOQhS8Si22i4XKpsEKId11b0vFm7uq7HyxQQMvv28/s7uiPIbtOzdVzI6jW5m
vYupnB2CHneSyi5uU8uE4azDY5WTlxlqc0+oS5yb/h0LB4n2MZTPzKLhAFpgt4Ve2DtDgkx5+rn2
L5qz3zS+Ez0H6O5jUD7nYMAO3Lsf8sTREu8tNDVte4h6yFK+xGoyctyIz9baaCUwrvlFWv+Uf6dm
Xzuos6AhKc4zYaygmYxFnEV4hX/RdTjwnuSuC6CQN88/UUouzwkf45IBKqCLaN9ynbBzYXwYd6JK
XuvQ6xd+uYX3wWzqMC1e96Pah3jCVFbgtO0HdSd1OPWKe7CO3Ks77OQe018KfWq9Xle/PRB3twlf
k8c33aaSxJkgNSz7AQ4V3g/kUtYg0DIwUo71qW7VnJJXgdliahDbWm4NPB+F8pDVTuNRnLWCgWCf
nkDiuR5O6pfCAIZri9yRfkCu3ZOX21o1uqGr08DVt+kVZXAjkjdj46Yo6GlsT35su37dqBIQDUNB
Jv0XDQ1q1m4Nqvg8UoKOcSAP38VlEj+2J+QSVkhvOB05zKDsv1tpnLn82JV5qOd+j/sv9N0TGH5t
KHPAia6Mlm5A3Op5Bf+OxbH/08j59bjbmNewP+gCLfaOhADbkXsVPdwJG8vGorBSFyxDhRyWXghD
b2zR3pfh8zpWVk2TwCf+9Lf6MZ6Vp0gtcEm8qZ7gflYMfRjDo5a4s0oAHjg+XVSUBaahgRXh1gay
4UwHQ0+ZE6uMHlozxEz2kEq1w2ytokIvhMrjKpaSRLivUOTu/W8gQdcoNlP/7ZUOZGV5oER0vDcI
9huchJVjBBxp+P92PsCDByXLdSLYPXjE2hAvEL9cIWRdeBSnhPMNpMEPz5OiKhle6/ObOrGjXRrx
Kqeh3ReyZYFxYuk6X548zyFVJPvkZDLtYZkbp3wmHXdRof6gV45WeVt9nnyvbS5FLSXk4beAvrJI
IPZVzW2v2SlX0uFjwQahJz+0nSmDlcOWAMoXdE9lVTZFfF6Co5LaIHYcIiOnPmAb0rQdoHpt9QUY
US547khjhsIWg5rPEIoQciLOSNFaAwndJXydsvsOEfmr/HrEflXEACtk2bd/R55awQQ3SqQR264H
wMf75YUxpdt+pKK73uyo5tb2aICcTp4RdvOx+g1lje93fMpFROjYmG6DH3frd5Z6OgFIXVta31Dq
Ifmaz4xsAanZiu4SxwFRqf4py3DOZ/5aw/9mlYFqZktQmR/J27UDZQViZf9xFG3KbURXPSKaA6AO
H3dHJc9CEqxfV9a6XQlv3Fs8Kq5afZEkdfQ2FzTsY/Vm/0CiBHqycB5LcjcuWAT5kxqRCKbOWm5M
EMRMGpXetvj8j+eQw9Fbr6IofCtcUVxK48BisXqacYPJOhd7krUklhQ8ma9+KI6E4LF+Ta2Or2Hl
74LEuUy3/eqJN/qKzG5HnC5fnNd/Us9XCj0xXloXmKDDkIlmZoe53vTGbshtC6POkNwQPey+3yMu
+px+h+jdl8gPnB5CPoy3uTUTS8c0Mjb76PQXfE1misHfaPKvw8qnMseXJNjWdIwFuZAfw303ddVX
hnxhFysGBpZkSo687HOwpqqes0ll6QMGL5zjPUMT2CPElSfPXDYdJvdbvYUPmOCzYYzXPozWlVvk
mXyfDroeyyomhsivnk54BASevfgUjbbDbPL+LbVZZaMAu/Ef4q4i9viX8B69u8J9gVOAEZWO2lzr
dqzby9ApAyr+SIJqtFWj8vwnNAccj/Y65FfopMpcnB3z/B4YFXb1K0BbF2hsyMRDvZ73iJc+8Ym+
rvWTF2JTXLu+NqDEA1u8YLgV6FolLSp3ijrGcsm+8uCcCfpuvPYOEwYkDYpgYBMPR9OElkF/gVpe
/9lx47dAJhB0qRTo8QrPeV7h/SCeVTzH9/XpThkTH3XdROARaHaqwtuxZTeVu3RZAOBsovoxDtvQ
u28kmojWXEH/Kw3gzWgJkG1qFTl+ylo8VaN2XMBKbRpzebei9l9VzZnIv4eaz5M8QvPHAmF3K7KX
xQAR3unV/vcXPH7Pw+p0zwmvBFNNL6VflSLgr8fnN09p9irepX4gDIR3gQ7LI038DJ7lL0oU3Xa4
kgv9SfjcP0ZKaeklBO/txHRRDLS5nGnmr+wiPZWgTo9M2CpP1v/kg0Kenr28/yEqJffi5Z5j/sNt
eEE0Y2UTMRP6dQOCkUSdJw4l2VQ5AiaE+/BoZwplsgAVGj41wltVFDCCq9B/8y+DtMB7eLj6E8G6
3pagNckl+NUG9nqPIbdw7zXriMfub2OkhA2fcim5+mg7SWqnUY4xwjlyB92iTmGSVtGToV+8BLJZ
uTVdxTNkhTxEGXBhxwnbMn2qpkW0f61IMBkZpR4OnH//90QOtS2yDOrZkG9KZwUJrb1PR5c1MeSR
0csRhZ159xbOvUXv6tpLZXNJ99ghHZtphDUSX5DoBiL6TkG8U8VptL8OEkh6s9Qk0cVhOx8Al39O
Y/FLwvy5nyAmMeoD/VKMiInWgb4bdf9E9Wwd/XnoyniBsM7IUoxM3MQ8uLrxxMYjp7CH+IXk06ID
WdnZU6Mi8QAQ76ErBEVD9dr186XlqBSZuSbUcHx7EOTUrMVEAoyJ4CBt2B01CMDwBwOQLnzB0RP3
YbPrM/wCf0jbk+Y6mQzFYeFeYqWHWqoHOOUF35IepYh3ITAdOUJj8VgPyMRISYxMx/vvpM0/dBrI
m3l6VJMmA2PEHHmfGUTv6WVV8AQNvdVQ7+YvYHFQEjTZTvCfwGVv8N0HzW/Fg4+ts3PYfi4s9tsy
/4gk8tZFhH6NJ5JHGplqh5FlguasPugdliS7yDtelOTZGJQojpm+VcfkkjjCZf1eo4O6dM6Y+iY5
ZD/NN6vXYYgetwYVfgcOuVs6MsoZC7+h6BqhuJ5n0z7Xn48jC0hWsbGOfGtg4+Kuw9OtUOHBc9+i
0O79kL5rwUPSdMXFZaXQP+UGXrfcU0lPP+qVYTXbTPHtFqJH0CkBPVTXibMPyqzn6Gy4TTYtmoBD
ASwOy1wHVY8/q7XCM4M3Gk7Wp7/WlUx7nev4ST5csyR9LKP7roIJL/wmnG8Y7Qd7lJz5kDOJpcgu
ixiPIkPDT3mINF6vaXxuJM1zxQPpW3Z66XyvVrYkREkciwh8SHBbOC1QKxbuSSEQ0rT+jSMGaQga
d/DQdFJ+7jbXv3LgShDdiPZlsUXNXwlTwJ0xm5/p/v3xGnk0amliWBReBV+qfEegtwpcYzPmUIQf
/BgpOZmRlFIw0zq8u1ZHI+WMefEl0FhWfXjJnCjuZ8sR6ik1L3qzCiNp7CyzLKEhu9BkzxomA9M2
XmKfjHJl4MdkALvwRp/XfuDGo5xWhWGTmmZxay8b0qO5fDDAS4KVX/DRvRXPsTLuVHEnKHA4l7Oq
9+HWLJeojY8Lgzm1E7K+JkWvynZdAiPP1hh0gFLvagUdqSj4KTFJbCEZwjuDo1ivdBSK7cICnd/j
op4tozF4GRZSpfbfrxASm4Eqw9tqViEcSZmKVCaHObPgYqFRsJUB8PR6ceHbEtAUFJQdh3Xyb+j+
bW1tulgZhxC0bIb2+iW5g3du0EsGHKZcFGtSHnLkkHQplAdz0VJ5A935vO9FOa5ecqwdZjLC1Zq0
/5l/jC2NFjiYqRYGYpRH1PbR38hw4fMH8+M050FdmjwHryBQ28IO0x7kmxb06NFqA+Re0saf4JIx
0GPOwwjR7F6+A5kV4HWb5HjSbXl/uBdlh39zCgkoLEbB2IlkdxaGpMwYOkQh78lc4W9APf8z7PyS
OXPmiz3RVsEjBiHUU7+7mUmQpiND5dB+2mf18rOuDu2+10w8M0HFUm0QeElbkvennhPTzcMgyp+f
1g0bsrvci5I1l+X8BRu/XjnQUIgw3M1L7AeGYHDgqgIO5zXHMVPcoGx1JBCwhh7UD0vDHM1oDFmg
WSIQI+Mnync1q3/8OzfAnUk4iWk1XD5PrM8Vrjo1abNtUkkLTAGiFr7AaCSi+ZiOpyS2EooZgCpL
w8TPfvGz7hsyiLvBBTtq6cqzEJgpmFS3tlhIqfX/03azFRK368YW01Uo7IXetubnUScMcfM3T/Xl
qCNni2DSvk8Uf2+noSptKgp1Gf35ica2LaNGdAW0DnaG4zc3hybBFi+G7XHqYUkoNq9En4ET/3Kj
HyuYs1V7BpHJvmJxNsyeHnFOfYuApaY8VlzZvomV/f5f8TcTuraQPQOjy3yDreX/bYVeG+BgMRpA
eZ3pXfRd6eiOYNdoVUNs8OXJnDqKhg3MGxH3IhWJQOKNYcFO4lM8+27HX+019nxxyKtf+Sjuxh37
6o79jP9lIEFRwRRUuzYAUUndySVBM09C47t8YUElB+Hhh0qUZd3mlhU4OL49/GMZH7za34VmVhHP
qO7Y6Vkxv8pOACjHJ4pS6QqzrtFI4ONs0ICNnu54G9qU31sPfdS58KmnDHgKxpWhWmimcRUKFi9g
pzhiOEmTjgQrDtcE3oC2h3eXw7lP947vDmbquGXSeRic8eUjdltL9DEx7TEhdA6YKGGlaoxpH8do
kpvkZdnTGGs46xVhmGZgn/bqEOUuMmyz3pybru7g29zZ9UbAZsgXU5of2K4tM6dRmjtW+X7gsAdJ
vdhfsOeTsd3SLDKpsceHDCoKZjkBm/DpGiEFpHWH+G9NezqpuIuAFoLj+ErlgliVcSNZOlHyh4KA
B3g8I5/w2WCfHEQv90paMGkrx+a79B1EIlQPcPuXFTY0KjJeNAEvC6tIVQX7Q055cKumdd4Y+0CT
+qtJPapn49Ei+F5KCX0D9RcNFL7yGnLT7u/s5N65fEAyKk/PJMoePjonStOlCFCmkJtemF5qoaJC
QHWXC5MQ8YPxIyn7pYkVzGbFFT9Hovsndsmi83R+yEUP5O/jfaO6HNjTZa+MpCFzEB4gMQwO20K7
WQYwHRYh6z8/0Wayjbuw5wCdFKlGb6Yl9ORnjzY2cuGRNlsTjWa9tRZll8V5mgngJGTVsHD+FCLS
lQIK+nU01s6fVNRqfkJaf7PRz3r2VI9vFNGzIata86wEaTp07L3qb9rIvdKcSdsmwnw54Nv0cS2G
Tu+JU7NNSW0WrUuNZtIZUAC2yR+iGWhj6dD2tS/W0Rdv9A6t95zz01juOcnorRSit1tyMcyxNTYQ
LZmiaIuO3/6k8Qrp6f9xlEp9pb0Ec+wnHiHjCvSFRDWw7Xjehk83NEI72Ga1sgSYqfhxpF+0Omsr
cmnKfLVbtIY2VMAY6Ha4S09k6HaeMwPBj1KOPL2s2A9FxuWNaRYGkbHewUjNuX+G6U5gUwfF0kxO
YFHlKa0yvpubJRSoYj/n5MT9/k5pRiCHeH59xhHrP2kaTZ649o9GcaEwEuhRkkfAHZQGEipBn0vU
QtLmICnS6XwlukqvFvnmMmdMqdhAw19sHF3qXz1bslN8Qo/bEfl2nbYZ4AReJB9uiFKjJGyOoIqS
BV4zeI8c5GH8q+mA0+RFbGAvdq1NCw6Vg2Mc8Nt6woAL1ZIU+ImYQ4XQt4gLBfk0BtZumshs461T
ayHCdYG8+zMNc+i1B1Cr+O37g9w/WAy9iQK0oEp/8a9grFRq9VvjoqurUYGulc0vf05ZhLEM5w/2
yG/a+srPknPcuNTD5oiRFhNduhrpL38JIQ1DU2xBIT6V/fSst2kc7PMzl8pK7hm76Rwj0K6viKD1
obkkBAdpdk32aVpSFft9zWlORSIblKzhUmVWXps0REk9lYaiab8nQFRPMc2g/QU7uYuTYZJY++sn
WxDMJKmKXgjpq34U19UwlZ4Ev+Plct1DaCgydObZ4wLSykCWJ2ear5w8ANEcNSTqysu0O1Mh9uiP
YLAAtwWhysVE+G/gz5WB8cjOX00D+luOYDz/FYsigF4Cx8ufTXsD+qEFap4DSHBk03/KufByDAd8
Al2Ojic9IlGy6S9oE5smB4t5f2nFyeITYsSuKOZFTCW5l9Vm8Fc+CT0D/D+fEgKWKII4PD0KHPD2
ydFevehf2Ncd4LGYaNtr7gRbUftuQwuL23M6dKowWdGo5Ii6uVAeKy2hEF1jI0ZlxYuX8VD8e9lC
DzRTi9BfP7FJJskOXq/FZ3+JCzCuhrdJtO1KDT92q1N0b4QHfD42LOtwFJHxJ+9s92csaNw9elqq
AXoCmzqVFhxTqw8Do8odbdXwf74nSJVOtiyuPOrO6z9TQAnGseeagipdxrWHDweFNl0apsgMx20O
OOpCn8o1Hbtauy3JXy+MXBL+PZYQXIWB/yRt8a7GvO7r8hiwfUsukRF0b4CkPD0j/h70k61sslYh
SwGRmXWiVJw2hfT1oGVh7MobZjZNTlDujRfvm63R1hZ/Oj+833K3BUIeVS95fjSP4Meb1YyxK0YZ
w3puG/swVb7t8RX4yY+g8Ck+COsgbkMXkZnvdj18HT2Lvog0XUNUMjDtbOFnwhc0h/nUKQAxkZg0
nGNYOkm4ufMdpNNTL8BPHNQjPsQHPeqCWmCEIXby2hPcXCKVN9ouJ6ZCcDA63Sns7EFGQo3po/H2
N991UzemWwIElZegiG4O+5hrYheOtJCeqO0GnCovzzGc63EcRo5qyt+E3IMakXWQrAMTX3H2LxhO
tqbI27cslRCvvqaTZCwk/S7Hba+0wjtCNXG3FgQmifsDUs9f0ZTxB6ioagmzIjDc9wdio77NyphZ
p1W9k6wsyMWGKEejRYWtmMsARp8ZDy5N9U+dk85UmTeYJylEIU5MjOqEAmR4xhwEY2ohiqwZHOu9
QQQvW3FplyRBdL6q/lbNt7bzErYb1kR0Q1348Wa+35Q5fIV5UsWAheCXgP6rhvB+sPtMrGRPU6Ez
ZqHKkER7jIcF2D5IBi9nf7r1nTxaHhrMjuQtL0hJ69zfhY0ISlPaWeJITVHhFGbFWIx3nu8qRiSO
SaFZml+M2sn9nsm6lO/yrKVvJCoCRzOCn9nUxZHlrKQqLPwR6b+htHzH9E3+SBUc58ZcPWlkxYap
Bb9MQk1tAwifV8SXykyBKG+moCw6ARraW/jbVVlAes8CAvOwBkiBCadMH4joaOBIi40r4bFkS9il
g72EDV19SEz2IKszTI5koLUCepJLuorrn7ADe64/rDADRt+eh4PkH/YV+Ypn7HRbfbFbox+N2BTs
c+e21CE3zBSdLQIXdInZDTouh8iTgV6fWGlDkyvKr0HyTxurNtKg+iuuGCJs+eHfb7cPYJaNNynX
q4PU935JHP2n7Td8Ej0hEn/AWYi9y47WiucZ68a5GiOqOTNOnk5+mgr4Dbf1T64nVgTgazF51M0t
+KfBL5sQZUZxyLmum8i3HEO8wfvQ4qMiyC854XZpxfoXz80w49C86UVIlK/CHzuCNhpb3byYf0bc
mEPZPmlL5P/c5SouVSNHlgM2Kf9Bv0I/ebmL5NHEoEVHn6DO4iS3EM1VA1gEW1HCS95afNDKP5Sz
dMU/AzbNi4tJPapOuHUhQ4aGotvPYLQBMqfNk/SrYglQWj8Ic30ihDqg2LTuTnyGciPEjjloi9g0
E0B4nXd3jw1t8EZRWkcilW3k57eqFkH+qOBiKTmsmFbDZVFFbDNvUM0WM58VQGQGGOJbfijqHp3j
rxcv0DrZ1aufKWxvaSALOK87uCLRUcQoW+pmHHcNsKmyz29iv34tV/79Z7resTp7v1Pntlf8MuR/
9F2tyB4QlWK+U0cuBvYjLoz4CBG8mSIQZDqozf7jR4v9yuuYwVsA2ynlpQ1j8b5zyZhrYJHmiGRk
LOlKLHuhpPb9eS8ocnTdEaU+RvB/k8j2vyr1SuzkgnPw1yIpNqhFtzMkChJ2JpfgxdNe0KJvM4e+
6B6oCX5339l5XiDIY18d/JU1IDOAH99f6MTIvr9qPJj6oTcss00VwCT6GhkCJYD5cArZHUe4ueUz
Dww0voLZG42kY4wliWuhMe3gqHxTLU7FWNLdlUAjyuPfdb6T+S8cS77+8w3eyOCaN9NeKkDntx5M
9NGYZgK25EU6pxkv5bnzLx46YTw8UTQQjsbMao3fFm10RGpiKbPrYGERsqkUb/mTpB0chto8sJ8a
wQjNn/YiFPqEJwxjeydwtZxP9nGaG2+gDEaNPHK71Jeivvb3t/CRDf+geTm6xuqjaL4seSOJpKX1
eybpN3QfChvO8f04ylYmwFKItIvptNhyPiuMWhIJ5H0z5GIJHgz4kZK1+4xKvFyVlrtJNbxH9QqF
B779oVyy4+D1JfZPsVUKj9r9rERnGwSrvE7ASU3rm6d3DaPlXwbpCr2dQ81LtC7tVhE/A11z1V24
MKB6Gm4mH4C6aSpX2F/+3iVvTDZtyCdCIUPCBmrj21db5oezhQIJ6mnvytRenH9HF18+CN23c3DO
v+5gbXCQrtiDvf9Smn9e11A91qMMqYeGYSKJPPe9RriRKZzuABslCYxHg1PjdJo9+R/yXOybm0sW
GaZJ4N+e14GcwTfZuFtHxTrIKMcs+trseHVBySjEzTYkHj4/Y9ZxOHuxr7HPWTBetnd5MmHCDfhD
BiFVfG6kdJXVUKMqe44qjE3qWHf3CuU8F+C/xHRBmGUARPxlgxUCvBhfOgIg/zLgctnN22Lxaglj
6qslJ0D6kbtZ8LGCzx6M5lBlztFDcJnMIXhuXz66ZG2v4wZpDsq3pD+4QsGxhAejstviFi5NNKUA
2nS2Er1+ROoGoVnjP5gkYm+pE6PMRgok6F0GdihPyj2kEvc1Zx+ETsqzkVHBiCqxw+/8Z/O9T0df
1vC/sNYHClKFTkzXOn0rPnTrzwptrTtVIlKQqWZtolKmYj/IfzSqaSYF1L6BjBSH9WXFMMyOFZ+b
EqijQobXLNxMj0mX+SgAO8GFzWzMjaUBQiD+d2sRszmbciTiTT+OxkUsfH0myp3iwpUfCv60DsLh
qigyuKtk1gs5QzFv222f3waBNnpai7LJ0BGKLe6hlzmehPh2mKq5E0mipsTCihdiuZyqzmz6dSAx
jlOHTmhkzADpfj0GJbGJ5mSoP1IP3i/EPLlCDcMEvp/5nEbpSP2W01bkdVXhYRwNIWw3ZB/wAXJw
fmfKVgR1zwNnpS9GvZk22McMpKrpdtvAJs4x15dEfa1lbpcfDdCmBv1MSrerz9p4EdXWoj8NL59B
lFbK9M4lwEsmBEetjCgB7jDKPtApYOPAVurGOUyo4ElA1VAzYgQ5H+BMVpKnzqac5eR9wtWo/TQ9
NZYi4b3e7Seu7Krq4fJkeZGOl7mQrCb0oqjPgkK7mr/1/NAYPk97eSuA5HK1809EUmTt8ug/HFG/
buOmMl0jJmfvEbmoqPfrR2ehRWo74YL8/sZAmMbvdpXrtaDMN/mCaAaPDLx118590UZOMcz02yec
5hkgJSWs/FofAaF++6EfOF8sGifdTYJEGdPAgsu2zAT7rsWXHj3dCiQ9DJFVBeutKuzeq9urNYrs
tl6by/bwxa10jU5/Uy9A3pxbhftz3DaBD+DgpaHaVd6TMitef6rwljDklsZJrb+d9TKYwievz1Fn
n67LS4GduMTxv7uML8Vg73kfPYlcixZn67wEN80u35GNUUvElZivMeCNBUfvne7eFKLOMQtIct/s
NMx5wCwJUSW9N2SQWaDOIwOIl2Fzo7kHGaroTUfFSmAKA9SY9UeDhFMbxNY4cQpVyPBXbmc+YxeN
tDlVWIMqmxVXJeasVZgWyu1vumNOHXlhJq3w4cmpCR4ze6XwNU5MkQ/fUmDXDSLnnBQXLLSy1/GD
5g2+2SvTKJa/9CCoHjIdYSO4gTBQsglZTVs8fwTqVzuL5ILr3kEHzF74B34P98bTjgva1s4A9InA
yp2Efljm0p23vdinTGX0whzIX0j4OWq9ps5eEC+yMtQhN5gFORCMjUc3wzXi6kbWnnRXLK9ps22+
da8gNEdNHexXc7CNa/n5rtR7j43awxp6sT3wGLY48vatB28DkGuLsGDkcRXwrQYGTYDI5uqc/MzE
DB4yhpe+9COtVeHvtS+E5/uFGUyjpHqslOCRuKErks9Xu6BEzHVLbkjWaMIKKRPe2TNs64fxyxzi
T2sv53yh8gWsrOTrJDfqFvS/HtHFD3JkRT9oHSxpN0iBkvHCT96yG7/LcE8W6SJj+V6RxwBx9Jzk
r1ax5Fdw/+mUheX/NARO8dMXrFzRersqXGCkPE9n0Do+2akJymh1c5+tVG7y9fL7otkcT05ZN9uw
KTo/1HOnvOLKsgbUTE2RkS8U5cwrrHjtcIlV6FmgFXJcHHEqs7zfzrfWI56NlLCub+7NATV6kV63
C5zHGFG1pFxzKCijtm2OZasE0vKPX16br7oiO05PPV+VSaTPjtwf0OUFvOMLjqRs3GgIZ4xFTjdS
NF3T+pSV0gLhx4eHlHAu/pDQgBPZOMUpTJM+dHA+OQmmWdP8rVGPnS2eh0Pclpk/AwDyiUkCkj1N
0HPSrLlSlMSKLwiysHXjHI5mHMHRhS0XHKcg0+ZvZ9En2frrFq5Tdc4ismnJy5uOaTITW9xTfC5s
/EpZHACzmXNjsMB4GhMG2BLKae84VYO9hIZoFzaa5+q1tZkI/w+Qhij7smHlyiGLNMDO/EAjf0by
tFIMRRKoHgkhZFSJepbWtPVq8GVNPydyBjU5pfqpttvX/Ie+Q6lKJjMavdn4QTNHAxMj5AeuQuS7
J/6Cg6cfJO0cr8NczXwObKiceDkjOqDnCdHcqsuomhWu7IEoplB3PyaXlW1on3WEuO5RfFIpRfnU
2D+SZoU1k+BSONJyQKa9yTBJhmwP6pdudcLUzxMUVpWKOTHnnFQQk0XvE9lBBx0vPnYk+m5I9qvQ
NP5/4A2O3Ex6bvoKcNmGJwfcBJCYXtsJCAa6gs2O5GRUFM6WHfj/Bklzsi56U39SkDVveDW0nlAE
faY2Kh/jro46m2t7Yh9MsMkjdswmMFk1HRaxJbtxWnZKsylzWFG1opI0C2ochJ/4B2s0DaJgmC4j
2lmTv1wCuXsmeLkJEF696xFpDyvfkLdJq5GZYpHxXjBKMFIn7enk6hQsQdN2eC7W5fKetgTjObec
nUHBXdSypmPG9v3YzDlwVGISYR4QCvPQQXaVp1byScP8Zr+pw3f492CHAKzWNvRJNgURetpQvqyR
BONigyK+x9woBLcdpku/0XafZEws3mRtLttPk32CSBa6kL/YaZDAFcSOAbIge2B6zGOlFft33yLD
6hREW3PvNZGNFBo3xOKz3+VJjF+IUwqjav4QhnSmZvdSeVRE4kNGNl0RYG+ufqv9KeA5FpjqDUAY
/a9OOFrHe3a88lgsZnTP2K9DIGz99rfhw8qaqbO9gpwvTtBvlh4hpEJzbCzFFU4w2U8WUc60L56W
uz5QdxQNy5Y8/t45iNpSQFEJRzaCEPAlNYUJMCskAVvzmeblJvipT77F9R+qSV+hD/fOvxyr9i44
fGGvx1hXg7VEqvh7pXm/DClbCIEFrN45JPHkvX0iy6TJmt9qWc1OgmgDIVXTsu2r8yOCG6CgSZ/f
MbZAjeMImXwsOdzaXVjum8M23AVIrYBhBvv7WrH8cKz7RZuv3VkHcslZC7PJTZKDBzHmxXDMtbHu
W7MyWGUfBDMe3EicGIezQXi/Yo3j2lRSIMWKTo6Of6Io+BfDxSV3cucucn4QNOr/vMn1e3Jsyw0H
HowX/rsUJVtvwENQpLMDrsQyV4iG3f1wR9+nfVb99TbSAhxxa7RhJsA3ebXYRHNEA9LnTT8ucDRQ
28Q2cgjUW7V2EwMJ2knkF73xZLWv8bg0DNsPO/j5sd9UszSV9F4xKHArc276R4Sc0pNmE8ESL0uk
9Sl8y91/E9c7w0H8hWW3aa8K3dPNDe7UMQKJz6RTE3PXHwSYDkEukwxUqR9sHKJVY6XEqaZClHY9
0+fW3t+FWdwQjCG0vO8COu9O9j7lha0GvWgvnz8JRlUFmTURuh5Txia2ceT/P2TO2rE43nUl6VMI
cXmg9+UW+WhSBEhkrJsHu1FT2JeuMjlU5TpLsK/BBipsHJUnumE205ljrjH56xkpJk74r5pwp18C
3AZqr1uOOgzwEltsBIgaUcQhGX6bqosNXMOLnA5XHWAF6DFGB66CDt0Xc7NhALbJaIDO9V3sde+J
2O94ViE/+hRCF1jryzOKDuIX85PyFlwG2xQmNJvAcAeuFOyGZyzBctOMjqfKvDj0wMQq7+aCzP/J
oL77XmVcPft1pPtt16N2lwg0adGyc05yaru++uizRhRyuRlNhhaIkwekz0sCy17a0Hyx/iU9mdQp
4C0jOZCXDACSS1SocayANoqBJQG+/FBL4BIePvHkINiibaZOdRvfJLkqARDFda8ZhEAIX6OOlfLu
lb0tSy+gckUvIR5ZcXGYgO1jpzA0KysCMJElnA6h7F+l5dUIiI1WpyxaMPP0V8+a6CLr1ctAnwZa
YNGz68/ZOYd2p4ZXzhlzFTt+/Sdiga2A3sDPvdrxResxuAgBFhcfgXPdPU7MH9YrmNvrefLK+N1A
xsOAKNj7ifdvxtfaOqoTVO5YXCUEsNrWfKeYGOYj6fpr92sXA93Oq0fKf9u/izKfT2gZT3XBZRih
unrwRamcdWa2dbom00jZluOnXgLIeTSO8WU8Qp6Jgyo9A+PWmu7GE2YHRopLXx4nGpWhtlfhaxDm
VCO3IfK4iFWSLR6tl2jCpLM2BlEFOXhITu0KMT2kJSa7Dt5ETEShkwIh3E3VbzBsucV2tqK/42H2
GYKNPVWLuKOI/aYA6Gh8hmfYMUBXyAgCEQGs+wLJj3+fU64MpwO//QWXD36ea8sMCG8s6wgqCNnr
yc8BXpq+SnXiLOmViY9dkrxYgdGjaac7RpbkndkEeOPUG44pow4w7jtcynEAi2ECj9Yhgu5nEpgr
SCu4LH/fpnt24bjdBVZSlLnOLNYakEzMshOphGwYHcpGFD0FzZDjmANIrjahw8mcTpdT5QZnXsZD
FS1/Wmsis6rLpgsMrjwhPfklVzrh3kg0fWyTIrhlNIUuBtJnAv0WfWf/Eyny+dnG1UmHnw60PgFd
5zY9/O+5v1mKIV+V8eMMA299vCjhp1pb/fY9tzbjfnhjmXeboXYOTVM4ZrKvo1516sRdBto04DuH
tO+OMhQlyCtOCGW07qwyGOvyBApjxBGLDOYGqeGAcCQgPGXJyDCyEWLcOXbWhFe9epSjCUnxbp8P
jelhqmZKNzvJMlXofuxCRgWGzqibQOtRPCWKAHgECJ8bARBUnXorGRCrHPxSePRcMzcvAJpf94OQ
bkbdqZFz/R5oZhldtXEADx5NCQeIjllfT+ovrrhGVyRpRGfflu5Q8TritmWwGLuxAclIdLKNB3l/
lce0MhI+JpOLjWM/Ym0Z2JaZBWJyR4X5LGxrn044AQSd2YsRYbGRQpIsXY5dPEBql2uVgfwoq063
et/EF1n9IVjNW0MRE6++YJjiVDlLgQtmq7MiebV8CfZQ3r1jK/Fn7A7N/9l+HeuvfZEm+Nx9ql5p
bO2lgITEkdQXkZH3VTXneSiNjKyDaMTniyg7WWWhVkDjlLz68y2SaMKdP6WqcgOQpFGhRfMj3cGn
Yoh0AqlINThuy/pdcutBTV19s48/TOq4HDv5YQ+oE2HoZxA3H+2lNoDWr9bTGHxFkSId2A8pdW1G
UorCf1xWtoBPsd+DlPAwjyv3xNSjmFIQVDlnRsQRTPgbHqVR0rhiJAgE1xT1ycHnHvepq1BxqOf6
89xL1ZYW6TKee1nK+T7MIUS1zriKBjx71qVCxoMw2sSi2oOMUvgrS3AUe4nZjNdvKoKno/cWv2yv
3voBUp0Qmud5iBQMUy6b+P7x4E8XeHGZRH9q8oePOUZ4YouKxXpAMpdJ7yI4CMl9vLJTL56tvPWU
hMQDcUE8STAym5OYSEEIfxqXUsRuu5pq6Kuk8+GZeUq72Rhx/EcuyXOyexsUjusyg5cF3Kw+hGhx
Ul5RYuXOoDXtKhQRX+bo/iEaBz2hm4LPPvOi0Yi7oWZ1d4JLBkjAxq9KqwF0OGNESKNBBC1BdydT
mrIUM5VjUeUmyEXcFpGRY+ApyWrtT+YNoI+pOEJpu2AcSWljcauogaIGRTltY+wvTCq75gxnTpd+
rylRSG9OHPGDPJ4aXm/2DVe/JQytfOViXbCr4oxF1n3N91HW3NBGVzMr6VykKmVf7xU3DIFAU4hf
bZNzoh0sdyXQ3XuEIYwGb94fNStiEoK3za631VQWGwVfzlk4tY/X9puN9Sgecl1ZSR6KSdTRG/PB
U+XOWdByyAOM4pBzfbnzsRR6KoJzPj2xUXWLc+fvF19JlDPQYzw08kX8DobM5KQjBTF1UVUdY0y9
KCZO4Du/FAlUGk3aHwhF3jN3ZdTp/HTpPM4e7XrVcPJuQh4TJO8zMaG7Sb5UIHPmqS3+plvhDoKf
B6ecsLhWp/P93BhcnP3wx0YAdT6EUxHIQOfNa1gFNwBbDP/4DX3NN5Y2M6VtJtnC0UYTI7zIhe2k
ibQAneNOgDP7Cv9SnXkWfkbtFj5g8cIeAFjVuq/WbExtrQn407/Hu19FipPfB/FrYI1TCHloSOyx
wjOKxaMkuieysOneg+rv0lYeEOAp7U58liS/vlwWI3R4r8qDVUZ4bPqnHYrZq3yfO+jDtPqmE9Fa
1OhkJZoOpPUafZqJnYw0qkKjQ/drzK9dg1hpb+ryrkXxyupMJq8BhewV2VjZoREhSW3Jomh4VH2g
Qgrmg97aJjIhG/JnQuXKVJ4zIlhDpIiGP42zJpdyyLdGdHskNpo+T3NCvbBmi2gyFUcP+utWm+mw
sEM8Psj5LYWCHmqTIc6x/MzfjoKtQTQ0mA/pl01mwSM+5BDOTtPjGl0mhCroA5HEVPx1l5AXchSJ
qT01Z/FbzOJv1vqyXXpQ+I1BoDsGnAZSwc72MmA7KfzTHzddwzjXADMuRaPez9Md4m4kJY1IILul
AKvqYOefCw42MT2N4BTZ5m4n59tMnIre8LBp9PoRt45Xs6lDCfCl1C9MbFGkwGjdsAlF+Te6eLvG
+UD8ti4QmWeLz0z260k4BRjJfBTZHPIj+vprOGW64BO1twTgg8jJgvvdQSW/DsbJnQn7YwPGCczE
CyLqu2IOStcZYUUXIn8dcS1DmsTE4hCmC6Dgl1gfGpdN00jzHqWq/7xqhNTJ7w4BVLA1WIfbzRW6
ncZOqP+9npmj2fsQ27vjARrsZ4R2W4XJktMrJsBZG+Cog/8qrhXkVkqIpMz7uIs8gUDiT5vXar9S
VGit8daYWJYWg5YIW2vso4YtHk2uLVSTDQhLUI0jK21XWyEqfoR1gkvkVt5ujm4CvZ6+eezGJfat
Tf1p+IVEBax2xzhqbvwy2Fg3OlF1lVq4v81ABQhLQUc3K/ErPffcjbvQIfTYeZw9FC6rNtZTgT+z
w7Ys2qXJ9D99Ugtp+E17LQbs2VGRrLlB2oPxedDt7glsFq/H5w24I8oFMDI3/KQV9THCMytprs0Y
2CJlYFhbqTVua0Du1nCG3pnqYnBqsfe9QqHdr/QRARBs4iuhHXfNp7VcV+FAmeKC9ro3BZol6kai
jt1seVdOMGyAY25R/yVfX4uIRJANdsvjI6vPNW+MsPWeIRDmGuCOd2xoQOEggdveKvfiVKoOxbFQ
R4UT438tGM+twXNMWNGTO+MdYHAvlbzct6EzCVFbQCEUQ1RtiPoJg85CX5ZLlqlr7skegJEKyK8a
Xj6qQlyrWE/qiMGX9tkwYe4k1NC52jFumKtkC49rYg21T/KYsOGVYix6iOi6QrNCoG+3pMh26AkU
82FsmW0KT5JDeY+bhV2K10L2cBM3QGJcXj7SOkpV0kJb4sXy4nD8avf2R1y4zsyCGe46g1YEDwCg
e+b9xs0/ngAAZXwF8WFgKzDKN5MlV51cvfpIk2sdXZe66l76vNDIYbDpwtiYLTtCfhWYTBhHIB7O
tzck9o9YsP43HydruqV+wfWqmtZrDH1aWdXvttYywJXAvJIcj6+wqxG7U05aXP9O7Kc8laQsHlkO
ZukYEySD2G1YCcrkbD1KiJm9KMofpaGfFNRxH19u8E/doRAWVbOfqDCmQKwl5mQEUqu21ta4ILFi
WmToY8f25Ao2RaXgAd1zEpT0i1uOPjZUStoL27IAtpD4wTk6Plq9ucgNQ1JGnTtaUL+V+FBn6JEH
C97LPAKpA7kVgD3XI6ScyqYuAtgTF1DBuTeELbsVMZq13cs1QUnfiEny2ip00QnDnl8ykPTfG2Vy
k+WJha/DO4StOEvkTxRoUSAkRtMERJbZl3m8vxcmLGg3uHk/TTgcrOKdbxl5O9VGveVsC2fJS29e
CElETJuY6E7VLklD8QGFN5mHutmWvi3s8FIGCBsF9GiAL5yEXFV+hVMlpAcJYajw0DxxqMp13Oas
fP1J/OU7675IzXlU4463sJfYnPhmoPKRTb+Eyi2A0rCZRgAVbipzmAuh/8KZ8Nr5zo8KH7EpHt78
eoPtkAX8MElch4EGGtzbGN74dc4Mxe45d0N5qVE9wsqiG+vES42/7N7XGoENGchmjVigGeEHYood
RnRN5QlHC3PcQ11pCIpc9HpK/Y7J0IQMuoMu05b25cCdLcpQEFE+s3p6Ec4P2iPur9ddPVBQKN5F
jHNUqcv7UR4rg+jQ+/qSdBXJxidOmeu1zvVLAD+iEmeSkAVcxTekTplOoaVqKXbB27rMXG29ts4I
DgtmVJyXaa3AllnN/TX/7pcuC0SWXkn95rEPzgYUabVbjYHUNIMrLXgCyc06S05ioNQ0rnVRYHGc
a8mjg5aCVECC+PjJ0+BGGlbYu+UpxgszK9vKFWDmf7oSJzBzKe8TQyFKgAsiJfkoVvDwixAKM5YP
Lyx9LGXQCfBV1KaLcuAdFMpe1l2vG7BwDoDtzBVp9wOJ6jALzzE4sX0F9wkrpdPHgN/iPTbvmYE/
6WU5Ms7Jhy0ebKceGmqRezpcC8xp4++M1DHlfoycZ13w8kltSm8EdjsUTVfdPSMnR1RNyd4FCFan
BVGbtrwq91q3CpLufCl/7AZ4yZ5tpQwcTQgvzbdO/pux53GHHxBDHlAoUIJFakiBjzfXaqr2bly2
O3HEtLyoZDuogonB4710RdBypTSdg6mpZxIKBzhXfHBHC5SEh/5SITuLbrCzzZZ+6n2D1S/KWspS
vALDdvALXmsM43IrZJ/ssDHdXBIYrB6do012I4e/NbuKadwALpqtjtkFnHbBMoqjbb9VSUE43lmi
swp81LRx0m7Mh2YyiGo1s59uMO9ySDEiswHC4r2WUhaECucr89OZ5wnxwwyy1K67WjeMmggrUBeg
u9TPDcOliua7fvA1soq8WAcHXEoSjv5aFf+UaQ/irVazbs5jJ9mr+kQKwhSR7Jz1dX4Ew1Wf6foE
19Oc5bjL85Wah6d/XmICr35O+8yd4bGsQRnv2ZAj4At1/kHzGYlQX0Px8EkGC8kYCDHYD6IW1VRY
goi96Qxv+1jhtd0aKUHC+gewQVtQfMQKKayAAyThu9tCDccXG1HTFPDOaGV2Cu3hW9qsrArsPD7s
4pfFBJTpHnaYubIWS9cjkUgpoEo3gmd0NAs2uS5w6nxDrwrJBV/357kbHeOGEztk9vCjagT5oHxn
kJq+tmzXI0Vqc9kQNZELrcnTpf9wuC5E2CfBvmZhRzNtNYkUjHSjgi0i4IyHGL731wTD9MEfjnnI
yyQBRJMmAWEDwnIG8xAYsp5I1l/AY9ZPwP0+p8faDBEWqyCbmtD7A9vw7bbBXt/mrUAHeZ6xGrAu
S58DVhdzoyq53HNdRY9KAGO5q5+mYhB6BpRRcNwhcd5dHRV3FfxPbGLRGy73gnJGEhqDjs8IBNEL
r7qcMAiCcADbx1myiQO22XjexEWM1hcyMQhU+/+R5o7dzsdtcIzwgmAqSQe0zOMD0y8skS4qD3S2
AqRuas5Q/TKIa6HeDxXE7/bq+Ad3GX9JicEP8Z+QBQut53HlBlPgMdkdKJD1PswevcgjHw2P5Ym8
D/r5fq3sznMSv1uXKwsPQNRaO6LxnLfjqYtS7dGBWfPd/lQl6j3aY+D2Pd1Qifn1fRKcqrdc/Tdb
SsFPHwYGKS3IwW0Wi4m1DnoLFFz+U5qfTHw1TLEO3iPvhc5F1bFeKOjgmmMg0XIHIF6Dkj/xuEB4
ejs/+gzyQptggARXr4D0PFWcYao/EKbNF04+OJRZGso4XJ5OsiJNG5o+047PjzBSOwxYHYKu55fl
ONd3QreoJW5+wXp5+hpLpvdNLff3BPRmZENIia77Vvlc0hu8AanjDARwdtoh5jP5lYsfB1Qj8VYM
Ken2gJUt1O+qNaogB9PYbHGwPXV+WG9ERFFoG2c2OchSW/wrVK2GGpZfX3yX/uQ/naE4VFnYjwpR
5BZqB7L2LRDMeM/nrXd8obxaYIjpneUNbMEp9y0XyAnBR02vV+/Ma9eiBgUEKYfLGKsXxxLo0DDg
k1IsdHbe2bwROft4uKhbp9S883sIDwKtDgN0flPNJFZgoFzJCw8F0znZ8S9OPZRDd1uyD59y6QX5
gthCRnkaA4ifriUq5yrWrudfmiCrU/o72jdWbo5L1Hv+L/YUlHo5Xz5ESZeCvDI7n37oktp+QiWh
IjdI3sPN8zpMNQCEtoEyfQEaXPv6baQa60Uc/+7xQFnUjZMnP5HsQjFpqJr8jfKlLjhQYK5mJSrh
WoiiAbP5WYxJC+0E1FK6H6RcT2izvAXkG3aC6kZtNCFUWC2tTWAwN9mrIcXrNg6oHdC0Hp1STZ8d
aFRKOhD4i0xB8sbONO0KfiAnjqH1m9/65UqkCGuf99A6XG/uWstArztrpab+62xnjI/8iGiBdrRX
Fwqn+29yRTQyS/Ub9lrJKk5ExeuPLicOJQ9G4JA5wZGOpeVF1M9FNilSpggCIs6nTlH2ErGt/stX
wDmUqk41+0LL3O6DeZ2ZrVl0TkdjEYhXGSiKq/SVXEwiP9dQx5i+AWNIeGU1wUAOGZ/D2nWBRuhG
7bTidSKyQMkDkOq9iuS+QIIKmQe981PbHQSJoX7s9NnFlTWFWJEBZnpQmnPbvKs1XGfL4VRyAC1Z
LJfaPH3MO2ss5qmjxR3x4Lvuqao80zBzNLkXhqcz0gKz2jJOHKrDBldLszt/1M7VI5q11zQNvjGC
D/yMSSbtqPvG/NdQKUXbRG8vvdu4Gh65iynu4S2XJ+yUcmsC49SKYOl6BBpXcGQbdzs19eQvkk8q
Ekb3T1+ivR2yLFfxs8PsxT8ms4oFfIBWM5SwI3xcefsmSmMElYp6UYCyJ09Y0+krrCVUUleNvbra
dR8p5TxaWx5pwT7Wz74CpQ583nVUNuPNrH0iSrO7zbgBkI1/L4+AA10iIUzuwYg9PJ5jHuIMqPZT
q4aE2nbIQ1wFL2x37UZ/s7mI8UzA3itv+cHJfHb+Dy8FojgXipEv3/1vXvH2uSh8TZcmdsp33dcS
VW3FipJc54z8n8vkSrJD87lwk34/OMms23MmjHdckMUfu99HgDRoF6DCYMhsBGfVRHaJogxyIve+
q/4vZ6EWuwDp84DqrV7lJyXQr6jzlUB9W/WIP7mHpDx+0iI4aFw58c397Td0UnKGZDbE9L0+qxwu
Stxh+tvmb6JqrcEB/DKxZNjbAwugXHd1JJm6CokOb5gTAkUoQ/NnMLB3gHMtY4zQXgexUOY9ZP0B
PBe7kSwZYlPxqaGQptIzLCDH4TIq6Ijn7PMG6OgK/aSpXxbA5795ULvDmmm1At/wBYulHaqy9uMv
OHPlGzhMW+DAc130TxNZ7ixh41ePg3SrPRSZEywbYI1eyLKaBaslvUo3FESo1ccgucAiAUcBnHSx
+br41ublpdLIU1DX7n8Y/WYz1JlTXg/MAECKur4nArKLj7cv7x3ytS9maKGkkJPfxxQDmyRKQ+FR
6muilmm8Q6cEixunyOWDabfs/ALPKQUIplja3VkcCLxvgeikTjBXpJ8gFikLEFY0ta84Ztz3uUgc
HCxMG0B8P3VyJOA4Tu9GAGLGcpGH8KzYiAg9wgCewZe9kDo0Ywgo7JlFn2JOr0p55I+et0VUP66g
gFiB14lmtZvvU45ZtEFGh9VAUyh7zNu428JdHfVGgG/3UhWT3zUNFTwM2oYfM3tQzwx8FlkkUolo
dnkZ5D1DkHxaSaXKHnQQm1+GkLoGYtShXX5ON/qcyfWPXY1iWhOH7TVSqDKGgiq0eZv++YW6eRUM
wU1yTVOanLdOpofWMCMLhUub81e7LPwR0bz87ONVHCXiXSawI7hxVvE4hXCYJYxvMsFkOmrcu2yz
M+jkvaE1mULH7XH3JA9SBN2asu9dpP6HclVrECFvVYmSIwL9nMBx+VLtr8L2vQzPItBfZ7FL7rx5
sSh4J2ewtW9+pC4VFYCugSXUpergnjlJgY5LnYILUz4IgtMiVF97AlLmHYL0s6BOUVu6UK4aTiSZ
A7pHks+r1DXVRSJt//lDOT8RhGiDoonO4XUei5mEwk6bPA0wOfy+KtOKt0xq5mAxWXrh5FErg1r4
026yxgMOurayAJ3UtWyefp5u6Kgjb6/naGqzNe8hwMiV39vgSEC7GuaUW2GZMG231MSVI/ocrVXT
wkEYiXWmIMZkR8OrKSlIXYYBIsAkWuF4gWuF89AYBt8ueRFmmuR/3LaycjnRMytNJUUXZj5wboju
1mo2A1boIe5IuCVYgtwabOdtAKZoCAvEPtYVxi6MG1vLttBzIi7HGNpsTbEGLCbHdHL8NacFOBVW
Mfmw8LAmFxr+vQWDQZ+azhdk+oxsOvzAde9lYMpIIsoD1bdGu6bFrDlKuPYTKEfSIeN1KDoDMLjr
cK0CKrruE/A0SrNTlH8Q2gEtNX9vqnXm4yzqbAMRE70F0jLEgStqLZd7EIrOAufiiDG+qG5bsoeK
7pcwN+PiV6RiOp6sQ9eGkTkxXMgzeETLAQpj51w69t2q1lUqEGpRjPnFJPLcPseAcjSU5udrWimF
Rd6kVCeWExIeOqWDyHFElOd15ly5OUZbFD37kO0p3aXGLjqQMoj8QWH0t6JgNHLMiYPtAj5iL/K0
Jhbt8aeMZsqCtZjMkXnlITxHX5iHDWHuPywOHY6icP7FZqCgsl9nogbiSjtr4qxyOWZyx1YnVrI8
RHKlWT0fxm0boWux0C2Wz6lcCIBt18w43bDW1juy+BsbQJkojAwwP0r4WZTbsThMgFLjQH2Mor3V
jUR+VLcHh22AaEVCXiqbXKE33zN4eFjp10islZ8n1mCGN+MPi2vGUoBLOjgjRZVfQBVbOKogqC+B
d2qJ8upkDYTQC/eAYv2vPmsm+oX73ZlelLXEyzPMKWuyxyTkJ9ZpIOpJ0dOjW495o150zndyy34Q
I6Okg54hiJzWcXUHjv6JhfqF3chaxz/vO4A//d4yD/LXzdNGBlAi/prfzxdwBB2jyxCiWpUsPzR8
VJNknmLr+4Pkov2rMLCzRePj+MIiH2AnOy7lJv33TDrBSY8pX8053qBl/Mmf8D6LVJFZz104VPhd
ot6f/dJcYY2q+QnH9zVcgW/F0EM88kFnDNVKgTzsskA3hz17s7lGX5HiI5prLtKTyvbduDOUimdN
XuDio1HvlHGQ5nM4yGy8FALJ2SV6H/U8d/ryYRMFwDRnwzxfagSWMVZUXcMFElpbu35m+lrGt085
vNXFA/Fer5t+oKKhDK+fUo9v/VGYa74WU7PtJI/CiJ0iz+veWM5i4vuenW+woO1jQvmT704dI4pQ
EvSVcs66gS2hlUDBRaxEceWknUTYIbUAXirjL7496ZyjBdAs6pPVw/dXLh4vzs53y5R+esCTZ0MX
wA1w2OKIl4uQF953nzAPXlzNT3dvlzQZIaSr9JKQ8IcO/Sg/68zkyK1VA3t88lTDXOS09F4hXvIa
YIa/bJvPnsSkpgW5n2GFJ+d4IsKr3F46WGod8F2+SYlV8ZjtY8aD38vP6BtkwNJW9XWX6LTHgxqB
Rl/28g0TGRHjRDFjuX8nqePl97aeW4vKL1iRVAfbmaMzI0d3QqjtBAZqQ+K2kV6ILMr4MLQI7O6P
qLu4bgPxR70vrKeU07tVQmZbLClQZRI4ltlPvg75hASBKVWDQXlDKA7fHTOKb4den7yzGc3zh74a
L5VI20rYyyvCM4ihoPPDQeOmrGvh50MGr6t5MhlUFxuxCzGcSa7HGxdypSIPdVInhmSvtsZ7LUsK
m8DNcZwa4RdYAQBnFj0/AykeGKEr8YVcGFrODRCCC0JLpnaUC2w9AdOP9YaHir0AHricWrqbaPq5
brby1LD+UujaQ+3WLJZ/WlZJIwD0g5R1TWwjd/zU6xtNAj5YNqMi5zL+7Xs8P71MSlbVkyUxHYor
JRbUu34ULyTEf0F/CsYO2KdTD0unuX8IjYTRdpoituSCRtzMA2RvkEq0tb0O8FfLrIwTh2oG6RdI
rOvr6j27iAHI7wEaXVaC0SjE3GxtAFygT/GXVmlxB5xxUqxXETw8AVQS1+YQHxRiSGewHaj2L9F1
oCSz6JPFvW9f4tDnlHpXI8lhAWKG71t4/YkUYktrBeZJRjBrOKxuX3o5gy3Hvo3p2l8Cy7+sgXKB
H9NoebFSsdL+NaXYySgmZcibFu/qjk553Zp8MyquZ7jWodFm0sUqnSaTFvzgD6O6cY1H1oOIZs5B
VMNLhFtwBxU+TwAfnLde+1K9yAw5O3ztmX0kmScAjXQGPHaRefYNQOln81E9EuXZ0w2mWuFCAcCP
KRx7ss+XABRD9TXAKUXsaJN5bDFYDVmwCFFBpykXqIbzf4xaDNGxqEGHT1bxnMB2/NGvCp3dUg3J
7D41dvuB5WQSS2M3w+VIAtWRP9IqSC79BcdQxrYxwGO9KMtzInXVFv7AXtyPOpa223s9N53rEHZp
6OFigfQgUF/5ZayrmBozUx5KnxQVK2M4qzoW59OXk596Zu5IXLQPA+CL7qC5+Pvaj5RqxHslE9S2
qLZnIXto2L2PyM/ARNqiQGVxxau1zXb/ICEaZcUS1mG+6QeMgWWVsdpBhPIfaalTpl9I0CO+169f
qSj8P/pceOMiGqqbXydDSLmpSuJES57MhjtET3P+KTN9mOt+3tUjt9hH8a/2l8o/Kqv1IpJB5Odb
cpM8aUTcYiNVhdCxUF6sAHwUm00Cl0HFFU1D+0XGDROWjvm0cjuWXvebWjxqzHJrzuBXu+aR2AOE
GtLCfEDJ0C41DRgVskDrrvCeDYMjzxZdusqU3a28innkGJlheU3O2pyvopw7jz40Jk4WqxzUFVTc
kYXAMZuQs4xjneGFSk6p7NGckYN5s4it9Ibmcy1djHDYeBUmyQ+p39XA8K7d9qUh61NGCxz3qsoO
prlMyscwy7SHt6rggyMB2Wn1NAuSHnd5T3Xb5yTYg8NSGscyIcvNQI0HU15drwg5AdKNiy+fPqEh
yk2rU5LW/T9LcgLFjrIEsliruhzzoe4NqDjJaVXuJ56QXICFJKBKCcGaiFK0pNZvswOb+Jpz2WY0
XSoa2EW5h++L1Vbpz01FjwG30O2TNEcuSH6FA+XXYufZhkyG+SpDQwtsG2OZNYQtJ8NagN9yg0pt
S5z1t9tJAwSOfozeWPZeQJ507Nk91ti5zs4+Naqc6P8LFFBooHBPHrNGXmikvBWHVGWPfJFXSVr/
ST7BOUZixpw0H9QRnD4jkTzvxrIU4gLZacnkPi8zAwA/dxaJS+xP5NzBPSi6fZSopiBDU4VcLd9K
a2AtjAdgyhyA7KqsnZIbZhAoQyqqHSEb9rHX37pKBUvkwLca5vtcvb4R6ksAwzR2EOnQONo0OdUw
GOzhccqHZtCO/AFdPoXWolRT3FWyPJ3N7zUPhQwNMJZVsnYey8Cta+iOpFVEII40JjDJKkCVBr5i
lwWGnve6GrcS1a00er20S0AlYK+qr/PQtmDVqWDHGH9Ig0CMtE4E0X8rjWB3+Jnzgr6kCXAftcTS
TBPJkqlCQCLpqdJzzTNGiLawMhRqSP+Afa8DNXgor5Zn3+LdhWkyveGke6dessukwuLpLSk/sECb
HgcDedKxc+HG6KwXVCzP9MRTebeOhN6WR4tWOGoA6ixdokPNVpkqFwFVqD/PJDurDAg8csNiB2/5
Nu0jRhxMipHMDulGyQHHz186HO7VRRNN/kksUy3M0a6nOHnguJN1FNOpzgFKUzeYhzC7f2ChY4li
wdLRBVdvHUlv+Q9FCOiUeIhMVcM40Ec8VS9rMuaArSwNEnOwhfn8zvgVX0WqHxF0lnoIjjmvKffz
x2CoNWUK/EOtyUmWf0RD5hKytQsuGUc97+j4gqd9O6yktAc6JOR6pt1AWcEoq76HUaa1A8kULiTt
g7lSpYYlxElynmxAXByQhPTVLFcHXe9/Gf8/US2iO+qAq2jYyafmVyubmvnUwxzwTypQhHJ8g5Jl
pSV/cHmRqdU2a8VJn9FskE+Tz66sqFkQLQd9uW9m2t5QCs8yFlnSEKsAwb4QoAupEJEGbUniCM21
2/F5PWfcj7ZoeV+L2zblldVuZejEmV8cgQERzLRvG4jGmvp3r4etZsWDFy7kxuoaFk8r1hkJFE2f
RLv3TiZBLMO0M1zhO/O2GE7Z4zPvFQXObgi81Uv7O6BnnHSE5sqqd0KYZGcFxqTVS5t93JqPlAXK
d2YccuLKRGfiFq0QByV6UPJ1qA+w6QuRb2ZIdExamQCbIjZL+sVuw+Dh85fDumAG92BnV9xreAXH
Pi5CuV2Sds9q0boe9lYGeSiIwxEDkZSkL3YcNpiDYPvUPB1kfP1Q6+50cXVKX9ij0DNcdoKoHzGz
tMFbYJcZne8eufuV5AHXixy5c2Rta9RgIhMFq0d83XmBmi9nPwIVhhl6biPshH338alAD43uIyoU
UX2h2NOsotiCVNSYm3arGwWZNgrw2tlaNAikNFoIeEMaP7ZO94q5Uuhhi9hjLUsFqWCmAvn/yOr+
XGmUS2e3zXuTyXVA/oPbwN8Izn7iFWeVbj8w9zTc5ZIRsl2C22uReYLiy9KObAdcLmOUZtU1UqKE
b1YaJWzZIDjSE+BySDvclDsBpI/tdp73QlH/UCCsQw30msNdc2v+3/VQjJuDEkbkVnRENEHvSPH6
1iHv8YFTiRZuulZR6msvnHzHx4FmS3Y99Ns8A9HubGXKGx3LK3dY6EMxGh/UrYFYdLUVcBkpFBZh
G837N0MM0uBKwsgU5BhZ4VNp0AI9aJ8SyJm+y6p7QSl0bgYJzuUjhWC5SE9cw/HIyGuzLsOei9hy
cwpFFyZ/kQJFYvAGR15TPYTRGHbMqYpKf2wFR7M0I33udhSXE47iWdFGLPbAC7CeZ8OBg+pT9CEP
NEcz31yi3mMWotlT/pUIvGFQUuIwoPhDO5QVtS4a4Sp2M5WP5F02GvaViZuYyjX6j3h0FJ37r83b
DcO+w8orY6IunTEDX6Rf7tRCETdCoev0wNTkYi6EoyWjkXjRAeNZHd7PG73QIOl1BUDnoRLYb1Gj
S5dd3VTzYZ1XUr3534aWqSDagCiars18TSXfjMPnOzTOMOxHOml8YDizwbUC7IK1uK0doFuQ1TXa
u08eFR1Xdvivak3vFTRsl1PqfQcPmr4uylZnuJvHitoSizqHnWnZicspbTCm3Z3EQ5P7/xr610Ei
aW6SikIdA8AF3BQiJX5fNWy8TvRNobMpr0HpG8ruzg4kBPwO8h7umO8HPP9tVmj9eKLPjGfFKDLE
Yliy9TQJWOb8FtIOApopZNKhUQ3O8/5rO2t/tbnxvbIhSsX8mvL6+H/4QDk1yqWZqEUNtdgTeaZu
Uvz6xXFxRnwfag6jQ8hta2U5gkgvGwnuDIjAYa+rAv1Gbdk750tSpPWDH/sTiK0Yt/qoPEOcP8sn
hJOw9w3GzZErZfCPbrFf1qT+CT8CPjOPN5vHXm/kMx/b1LExJzBBxmuoo9KWB6oecRrgxu3QMz3j
pxV/C1h0WgNsRrStU01h4I+Zf7aNrmOun6/Jr5yKTSc/VwG29KNgi/Dz25bXx7+WK8EoAVACZAwL
wB1EzcMZ/w/PsBZ+MV7aQLzwfFESPTbnyut4KO8agORzkCn8RoZRVE0fjdFdqHxO5D5g9Nd4XkI6
RiBEx53s9kC0vvtTKwnugyofJD1cdbR5mTv40ZwLTtAcnKpm0tXa87jEs4p6XlyDglYsYBdiBHzu
dPxR8kuiQ7vDtMJLzpQRmmFjHV284SVjtr1O9ZevU73jx5Jn0Hv8sX7M4i3UG6ARr3HFauv9tg0e
Joc60ExUco30DlJDIpy2LB0m+ujwpK2/ZrzB6J4z0HxfLpf5+3uwS709Z995tGBZARX6rbDAVh8i
e6sne01o1trw9TG1cz9ckVqZZIbV03ZZfHVR55dDAD6rt01cuGGhuGpbMf7921TGu6R1IpzZYZVl
OK5Sc23NWACTRUnyYi7H+oh9skIM2Jy3iOlCa6sdWtiIR4m0RQu8g2sCTHL7tPQPrchZ7wGwtW8s
ffSW6ogDQuTCEbKr+7JARCpMVFa3prMf1LpeqdfmZlEQk4N1FErVkwugm3YOibS7Cx4mXEwYVFU8
Jeu5+E2IDFAoQ0zSdmMgjNH1/p0SrJs+3ExsfXkrAXFv6TFuPAAsyz8eeKAD3O1jbdBRVaZN5aNe
QDa47h8wj/ZEg3LpS7l540Lez349ewayHdbxLNHcrYNvGklEzCRIhiFux2rCir41Xd5azmVQuvUQ
nvegF2k5lYH7bpExTKA639LEPIOghlRVare4ADkq4TfUlfSIQOMgqLVKPLELkVUFLihFUIs6Bi/y
TkB96yl1zTB+jzotwAdKO4ZkE7HJEu+Q7m3Zv2RGs2PGGYL3IuMLPhj7utA4ZiGT3EenUR7n23+H
RokaFn1xBMXqTGuPhIxprLLKBxbfDVsvk2z4kecUY2ubYE+oncXpUGZGC+EGhRpUPhhxdBeMN35F
0EcUib2FrG9j+JybyOq3/isEWTlknJxOjESi+WTQwRpPqkx/GOxEYVJ+vzqpgZuT7yJvOPwZTbOe
p636plqJd8VsY3pfv7BI0d00pGJj8Fq46Gn0RILMo+bGWLWE+gEefvOabJIrDWWw1TuN3YEzV69t
xSqWL3ApwQLNexDOsKJFybMi8vhs2LDVhSati5fU5OLESidQuOoH+NDVyW3rVIEb3GL7pRXRaPEt
mUxVvcm1B/dGf51XLO25mszRZGuH4oHjzxjGbpCBHTF9kOXGyHUPlivyiJNQNtgidecunLwl58lZ
DMpG7cFxzpuPOBMwtaXfefXiS/1v10YfzFvBDEFzqIwrMUHzaQkF01Hhqe/50pqTm6i4DQ5qzHCx
WQaeUVxr1RsUABCTrJtCQXJRGYGSk2pIVAq+o8mg2Euq0tQjfxJAQZhr2WkGZEyd00bi4wdW7Eot
vO0b2rpatMynDO1UTB8OHR0iJMVf6t0nbfAlA7cFXhyyg9izq7/3dnW0DJS5VgDnbPD+OIJcCWME
C0bHulfuVyTHhfcFIqbhU0SifEyygnrMpScFFz+0qBjYbfzrnUgeclBvfnDREEqFSVV+/kpf1seh
4wW+/od2JDgVyPX432LoyEgglUJeZm/rwNZsOlA47LjsDAPBk8J6IQO9+net2Z8MJW+2cGqQeB1n
yB/2YvVFkprQjZ87ZHlW93C3NVmEDaIDaFit4kxsCmLs8U2NQi4fe+BR1Ef/5igO6lk2UA44drni
PgMNvvw9OomNWaK/divjl6dChCfiWZfEte5adXRgz5S0XX/g6h/0lBAHiM4LZNMifKmOJrVdHeMM
aeLiGsVZJKCdQmRsqQKUJ7wy5vuawx8sGlSHmedPtFpPV+Z21EaZkjLgAxxQJZtbxavLsBHqP/bX
BLY9pjBcXWfOv9ZqS6hAGtSjYQNjsHNii5d1cMqmU2rwySVIMkoS8JX0IwFu9+l154pLsQneH6pR
OCCWETf3d+T5AEJDO1eWl93O+PmkC0yul6vYMrDXqtO5K3+edaWYsyz7zh1pTFpQc+91IHz16sPG
7NdzV+lffXhFlBd2rFvhtPZCSKqKB6lgTESDPOJkrK6BNwaZSXQM24OCl+oH26mPiuAezJXqnOlb
qJVMfFDH4PPoeJU08/emrrcvtjqmAAmhk2u++1NsiBmFnvBuUZwU5f83C32mHHNFXi+6ro+KaUtV
J13zOfMWgw4BuDn0NIDiRrsSdnAE0/Ea/NTFSHV2XEp3429kky6UnIcDOGwZ+TMNSAWuMmpo/Gx9
CAfweh7pJz9AL90Wsxla0DVdDnUGmY/jM5qbsd/OLND7TL66nLfK0Ihz/BSAYdw1UrlEnH9izjk4
dBCmu34nXiZxqQJX6u5/8bJa8d8i/T2sRDq0UAnrofGKJj/btGDKUfWwS00454yFbrLt1zzh1w4f
OpQqCuyxyzZfKlUzY/qQtVLcjHCH68gU4FHRRVA+ei3IqH2Yhdvi8RW132eV+0phKvPlWqxFB2Dz
eIcRSUroJxrF8yFwwGD7zYkniYqen6nW/jovY5oOaDYUXv3kDRq4YRWSVYCkvVAyFaEJrM+ej1Iz
QfGwIESXyEtbzaUT3h85LHpHhd9jPNsoNFkxWKFnqG0QdGFSTx5oqbQG6p+9Tl0dOG4nJdWyAFx9
XpAnDinOTZQ6wK1zarbz/x5uhurGNPcjevZxlAiTbStezu4itAuF14nP/TL+xP2AlZlzydjIgN9n
UYjzirtpmAA5LzAdYgZOBypi8THx6MosVxz/Tv/54YtMciQRmp9eJgEsVj1dwn1K6bQiYIPylhyJ
w17xY6w8ZLr/BqddhCQYmhJmIA/GxEdaBJTl9xsLq/CQqM+BAdDGRJyc0V9ohtw3WDGBYfEn4e0v
wqJQjTz2OXerpBmev7dfL0zxkC7s/+KqaQlOCW5b0w4gdhn2BVfh6fOF/5ikeAmMUV4vPy2bB+s+
urkcc1QSOMQLM+m+k2U+liS0emF+qOMKg+6Mbj6AuUNk7azFadKCUNuOadNrXBA0FLPhScIZBUSw
qt5zqTtDB/r9+35TQFCIZrcccBHJudDJBB7MvsuUwDG8hkzIccv2SG4Pdt5aLCrB1dkM14v/8iS9
jewbQt09X+pw9+X9ep+HIBmhdYSG/ccopu/qAFVtui8FYdgFqTpad5dcsoTuy/uyscAnrXxTmbpn
CpmYr0F38mPyIeEGm7aoGCC9BiXyFRvCscUNkxJCaJwi3XtVgT4Pf7spjVMyjxFsW2wNVJ26Kq7n
hzQV8c9xWaNKJUbNmqOCLlyCi03RfQljilhm5rMZN7TBC5OfIKKR59pXxDWAu5vLGW9yx8FGfIo2
+JXtGq5Q11m7W7Wzc8xwXf1ftDJZSjHKnMLiDrhCfkiXBWKapo92KmIMDIKXNTvCmZTeg8+rBNTH
HLdN8Ipp23abUluA9UrLS6R2FOqDlNGV6N2SXno+fyFXG6zBcpPpOdyk1TtvRzPoNNxGacS+AutM
VNnvamz96Y7WXc5CSAixAYomiavyzlWYqAYDge4y/CPM0GdXN2JpHNyt79IsjNHG4vUdF6xAcOQs
NJ1uUxQ60CEdmDBsdiXsmvuawtBZoTbCF5AVCa4AJwfw+/iQ3mAu9AzahQa8l/eXwLRORHkgfhDZ
FO60I/CPJMLotQg4FXUn/Vmkfl+EB2sYIHTwd3j68mXcSw+qhwc9Ky7ORcE89Lwxdzj1U9W0npF9
m92EIkjCZKfi4NXtpPrvKjVu1DoZc63Ljjs0aXJISLxyVH6iAvw7KXJeFxcQRYj9xb14Fu4X66Pv
jDUrI634+u9uPfgT3+PAg70W8ui3LhIo+U5tquhwrsDsrX3cn1eLV5B7g9yvWRGRemqrkH7N96TK
lu9suwU6ss9ZjVAtC1NVGbkdjjLvScJP70dgQzdVhhRAplcWJhrmk1xvZP7tpbS6NhDFU3VzZfRh
4YPgSe7g530ewWUvMwQa7ebrnJu3UXgfVAc3zj2O+rVOZvzGpoPJrFmZzKd9kZ+S9WEYhZjKF3Ym
/d+IUWh/N51VBf4dGaDcXSgUJOobseTdCawEUSYXAhw83bPLlAb0Wyib116+lPmnpQoGv3OhTYMH
9/3CsdmQpNZRp+jwZR29Ech25dexWlYQULZDS13o5Sm+G+jEPPbecgECzoFxBsES/yrWUY/UtcIn
qDeehGsaEOiEPkCpjaoyHbmK5v1HDKOtlrucs5l93XdGEeCc0tuba3fHfbK01HgnglReVUNOq9jv
hB2EcR8yO1XNpZfkQvKGcupiXRCn1WEk8PoG5M11Jq8jLOy94MfRLPtZpX3yKqo8O8oqlzu2Lztb
LBGsvYq2AxHEQZTdj+fEmu8Gkvd0GNCmEZ5eKpoDyNDMCdWWmoiBrjY4XJY+eruL9v+pUgw78t+9
lc4PLcyb4AMtWzqvavai19ex6Sylsj3d5WwDxkaXGooBeKBLcoPjQq7RlR5O6fx3tLD1OWUeH4HY
8k57pxrVmCnWlcwPp9feHnoMKyxMUzZ3BfNTh3k6v7yFhjaKuTnPQ10LmFl2p/6hC0svt6wx1/Zv
olSZm1E5k6caVYRh/UY+GxtzFAmIqtMA1R3Oe4VV1RPPPeTKfEe3ECApL1YvVVhuFQmZEbgoaMtv
v01n4j7Sax1a3H4T8rtG0DQypaoYgFqPdnuoLBY4MslEOTLI0718MDica5wd9uollkAIZFSqqcDt
Q5ZyQuDdvfm1mQLlH02q89+fmM0dcoKbSIQWM9D5ncIHPeUMsI5/jfTEYnqscR5HzllxdHQOJgEf
DZbx3dgkREN4Nc2o//esBClZ8FiJ9GNk8ResoUx7cChxwXOEOzJImijv83ywc5LUMNICrD/y51BO
rEdtKkHvJqVFsVzTmeCOpKTrEgnUbrJlvijCYGVgMAEEwHt8OXydWeQ66l7ipLNzVCgROYPblZ/1
Tuahu8i0G8IEFFghK77Wv+2op8n8y+xmMMgNlVfbcwt9q3Y1f9mUsU/AxNVDfmaV0LeOmf1Wg0rY
6YvllPjcS28ko9fSnMvT+d8NwdOADtUN5lacWAjK9GgHydRnIvLas9AcW47/+eoPLSkw0G+mdNa3
LKGHMvsUMgfP+X8CPv1/XO1a8ibaE966RbZxreIE+JKOCGBDuDyrQjtHPx6XYrqDrhgGmR3UO5h0
lny8PiC26GzTnnfnC3Eajl13HLuqaqSosUI8pc0I0Yz8uVlgj/y1zHln5fr5GvimiNThSoeI4bY4
XhmgxmTK7tHsHGr8gVc5eV2ske2O2Y4VvHpcPSKbOtOXhVp2u8/OetqgbubWwX037fNP8SdUBTZo
LLggt+LSjxWKKPHVSu/uihLLJ2adAZkx6oqeIwzZmMEnfCQ/1/++YUZeICiZiSHg399iib46kAIS
4dyc8RNlbYi7//UK8IWyh+2ePudzbkvI4qXxgbZZyOntRxxVfhvgLiaTC4TNTxiSWi1iSKPliByv
bQDCyly09h/FvzDxFZ2LHzhgCErMSJngGeK2LbWgjc5IjFtEbRRlNSe9eDbOjg/f2+YVG7x4aqat
SYzgDkGO3dyP7Obgk5FO2jqydlC5xmWFWxiAc4y+9FZix6wEe4aL3CejE2wcOU5qcryzUaG/YWWV
Zl0KVixMcRh3JTPj0oH+4SpK4yQSssXnBFfTm3vtCA84d0msO0be2m1AOmeyHwtmZWm/4grxkLLe
j3bDkny9xvvCLxmHjsON8ZGWuN3kvs4yI/ETpI0VsJTDUV6SjXj761HGpmyUyhE8IfbdDEO8Q617
Wpr7k4L2yMUdwTHOMtPuzPwZy3zUufzwLWVIx/f2d+7wTwI3SqMCxfTxVrqp832eoQtwuKx1mRkR
NgEEZjqQTw2wn8g/stQM7eaxrMKcKN+hVk3E7PnWOmrXS/5UffEprlKbtoJmJwi3Iluy5OFiznJj
lcQVoXPHc0No31dDi+m23WQN5xwawbmkGrCr9uTLxNVVZxHWME0LD1B8aW+arecSAcscXsDaZhG7
+aFaT/N10nZPKLudKiOvPISdQZF3vRd+/QUqCvO36E2Vhg4xV+btLsYXmXT2aw9o7f90ux8BIC1g
IDaN/i4b39nCfQWr5uWGZWdw+3ZR5TA5FbPofQJPWA0zmt/CnPUWE8nKgypnNZ51PdqsRrkRU42P
BPAAGE6xpqBVDQXb1Lr0qPQASoFIh5IcgBHwsl3HGnrSDC9NW6Co4PrcHypAqu8rigwJ+8sXZcTY
6A61Cjt4OQNrWlf1dLCvpMaaH091rtQypuJOFcFk0OE/ygM7KUiIdkk4Gkxzq35j1HCbd7ZWgiGt
787OVFvws9h4JpEjGhtqBuftSp0+jCdpYf7cpsvXvG6dn5e5ihjEmz7gMDPD9ZfGog8BCzPehGE4
4rNnGyfC+3yY6RR5B7zAaOe5w9XfVs7sgSntxgFVMLMPUWdIWoX9Yvs7CW0XuWnAreSk29Rut8Di
q6h3ROaZ9B6g2Xj1zRBsKw+hPetBTbon6ZuSQH7sqfd2CLEMkHD3oBOq7G/0S+fwKtR+HjEYT+dA
f5Di2I+NEJvzZlY1KUik6WBDHsidfBXytQWNx0wnhh58ASfY5P9GtvXgG9/YpoIGp28SMpylj9vU
HBC+yjNYntW4ZvqkwoPByKULzUC62QUS5b9V23zqqRnYiD3L++ZE0mi2dtx0q8gdNoKb8yuiGcW+
ua80MVZEiU2rbjpnsx8K3YfGvvv8hWzff8j6QszdapOP7PYiLf9EwY9+Gb8o3YEXuN3FAAkrneeK
BLlUOxW8BolR0fAL7KHqVVWiPGv1qNr9GEMtnXGZdvViwrF6w73o4UN59OHVyzREMDKTDgvzIEFk
N5riL+S3OkY9lJAjFaj5sk7MBGWM6TLMSSkfbHw3Vf3raupnjOp9KHYohpk68zA1FHtVmueo7hhI
rFPoIyaW46lkSrgl997j8ETPLdxdUqnXOvq9/qtitB+gX3nqZrlFjOnpi/UhzM0Vv52gP+EpEWY2
cROVOGszAu+H3+JtBSlUkbhG1E3UkYtw36FdaeZuaSZNkVQuGPKZY6HQDRO56+QLfnpXQg9ysDCd
3FVzlPIRV6YhfHO8dlVCFY3lO+yf48veIyyOVZACKYM+cHmfmzbvpXF9E7HxgAE/43dorRoyI7qH
RvY/uYfXJVY7JLfL+Ao0EdY2+wWZ9/HOkrlaQObeA+VHjRdC2xKx6v9mgzJxp5uT4bfn7lPPHD9d
rtCsltRuKySXwPV/KnXTuQj10yZrorqGjxgVGZ4VXDBcvXzm6HSUAfgsAB4xhKa/RLOgjfAfY82I
oALkZxB2P8+k1pfUFBl/KtX2aDRLJvhFy53tXoH7IhuWW4jc9B8+bo7bonR8gctGRDQRCBlmFPl9
VADmzfHbTwd7ZncVGy7a17YQojQz+7ax+OaoYlVArnmWlXMMxahlrF4+qOA7QhFCq2Qcd7E4Fozh
FoN5aBCEJHkQwkGos5jvY7HtThcB5LCn4JWRdrZFlHHDEGE9TBACGm3Yw9BIivgZN59b5eQ91v39
nU+EuXRCQXMUp++YiUdXVyJj0ThXCqCnyAtRyvXqFrlAjdOYAp4USitK4qgaJtcXlTQiNoc0w0Ne
//9nAZiwtgt4/omYE8usnAY/U76jetqxM+aMlUt3gn8PMesI3caa/dxELmqu8jYzD24sIsiiX4D6
Or2jNEOTBZAJ/wrPP179pd+cB07S/WJElSt9LgeHyinUKt0rDHZ0behdzBAy7PfzHIgs13jIl2+k
mTh4WW2bOPm9NMb03uJm6qUi4ciSfKYaC62WRU8up7nd+YwykvC9pjOVH1qfpePji+PQAotM/OFG
2+MADb3/WFYAOUXkdmRRy02LfklCxd//sZ0EsQMp9zaYlTSJZ3YcC1ccz3pOKD/cA9ZXRZT5bNTH
HOa0/gyd94/Xbh3fd0MN/I97YkfGaA3+vEPFGPS7bCcgKcvzqNDoj/ulV9jy1Su1LXIxGRdzZBIJ
tgEKtYdO9JA71uMnWVtn3dC+XKIqkvENBlO0E0Wo5KeV1m/wRQ24a6Ca1VZCALU0U6+zmeS3ngZ8
Ja3C+xUQ7ts6nn6H0AlapF/DJg3uNd6ghnX6rzKvegM6Q5y3qhdmD3IQB0uVY/z3f9XW1DOyzIwq
Dosr0o2F81HIqJ8X3KEAF60+tKSb78nG8cWneDvwOFPwo83jLPZGVo3/yraVV9QDEylixF+66vV0
Vdg2frVnc/wlP2GRxc7C5zB8vvzAoz/fsNs8c9EOjyxEeZFFUirR3s50z63XOf324xJKjBuGiw+K
TaVJrLdhh8Qr8ZKRVxJt4fgOvzTssJlhuTGxb9ejoXN98FuehH4mZnJh5/vPV7CCimH3bLIJJbpO
Y/a6ry/43Ktho3kBs+eQIsTZU3u++bkNu5jlVHBRzh+UYfifwSBx/KuPmbNXGYNZEdvjwxhruWxG
0dOlU64fNtnQ1pg8RcEdeSgBZ/3YZSvp0tN6l4CYXCKniWWXQNTOJlLP//Xn6XUPHQ+VQsx+GFHz
rzcNKx7jQGIVA5BXRIPyL2YpPkBfTxMZRnKMuPnhNNiA0YEAy4uvZtyllSTUfwCncknX8ugyVfJZ
Y/mq4qQ90IhP0xz2IRb6qr798GyimgLzDa83KHZOTVz7w/siJ7/eSf2UXAfUx0jwZPGN4RO0vUA2
7KjY5ub1739kGw9wxz+vurtcUq1X7e8ICWz/7k3KcIhV8lpuGYeh1GLMzNtH/pLIExpK8lyZkqRZ
QSHL7ks8cUG3Icb2Upl1LAoFHISKOvWl2uC35rumgzAeV1KpHsQRC6qYSlM/nB4gpkNIDGeJvDl+
01zfM15//BK6sITNYdM6AOs4wyfevfmvGjtk6XemQ4qflYsx/NRFzDbh/yFMP8y2/AErSdjn8unj
axaz8I8LnBtizXu8jWTCVTfdkkvYJzpyZUhDJ5VhsaOns1J5aIFxKnwIaXEijcpuTkf4JO91ZvWd
ELNW+8ArKFcMFrGlD7ZpXt6jrSK62fON48umtmbZ0nr2YFJz4QS3tHn2Uu4QM3MxADS53qDI9Hb4
PDspI3CGnFsALlr5JcQ14gRnaYbT51wBi1BQAF+sraLYtL8n3lJ1gyAPoe9pioigQBL8tTvbbhgy
2Y9u+tGJwQLlYAp7Y3vevZCvS3qfSinZBDaGzKeELhDk6LT3Z1I0vnwkIKIINdpOI1CKFQmv58ui
20i7PSOdceiSMX5E+ImkjGby6iLw3J8QtTjiNuqpO/wdh6kCCHcqIuc/RkGSNwRB9lFsKlH5BJs7
E/+whHgmKH82A7DA2mY38s9Eurj6kIx5m0UrHS+uyisYh5pHio1aUUwFgAlyElCbp7aFWgeDFRll
kHnJnI2tFRdJsmadl3AkeAuS0juv8TTC6yVf68qfLAGlWvA8Gq3xi2hO/5+j7+CLxQ4DX5hHBtur
Hp0wIz/1wK+akeYw1OvYh9N7jU1NvEzKaQWc+0ZAnXgLetCVhy6ZEIygvPnjeAqARiRiD1YGkWLG
SOAWMTPNCDry4AKlCm9hjEhMh2JcVWwS5za/xLFK8rTnTp6rS4uMvXVw47w+CY9j0ttw1ya/QK96
4Ag4ehCtnh157up+r9YSSxVvPXBEtD/py0yK01yxYGcdb6w5pPxqiiu7k594U8vcJluhAxlP5AkV
49Luc3E6fjRHpVyagMoulbOqFLn7uVfYwl4jXtV3P11De6HgYftGWMGFG+G81KIucaaYpSB4TUBa
pL271EBQrej88WX3oHYSgH97CibfSt2W2Gwzw+TifrlYSTdPJf72UDtb7ew1R48FGeM58X/+Bmgr
Fmw/QkLVLEPMQk+jPPJL/4Wk3b2R6sglVHOT0CIlKHpj+7ARLs+4pO0lzwcPt84kfqvxxpSV7fOA
LxfS7jpY/UjrpIO13DcvjXlhMV3qeTASzyNFKnV78QF7sXlRtIygSlQUeo/mp0ygVbz05qnuLsl8
G8fmsxplbOMZIokWAeiE/YS9Rf4rM+Z5VUnyGkz51N4i2q0TTiUhLE+9T6W+sj8MzgkFd9vEl2DF
geXi3Jp1HjFFf+4k/a8fXERjfa3bw2ycASQaKY5Ta02ozD7b3dbTqUWCqF9kdyrFGxpoHwav6Ihv
yGD5zsvYenyTouADsA43dXYwx1350JPypnDIAAQcfZSlkkLl+7UajRVaVFyCAhpbjoYAdDC0E6AI
QQ3KLPQgmc3XOvMVMNsV/JDT7EhiRgtAfvWIhJqTMS9kJ2viXIg//00uoY8UWsxVs3xiZvopbD0o
E4KQT6KOA5YbQ7jniQNnqRnhgL985Itjs5N7zJkFtLk0zP8p+vedFW0P+e+Gx3Xgv4RkLd/yqb9f
UbxZ7Q24SulZJa3Sb7gib/c6k9/zbFRw5L59DvSqwXeQONkgSfocI+nrWZUmQtLlmm4PFp1IIc6s
yHm6048OjgkPiOWTtJOCWQqlFPTaLb296B/DMjBEhRVq3lCe2CxrCwQNwW+iOhhN9SbRobFhm7Ox
OnPfvxwJKHYWJW9RQLiUZEOs/0DsS7UgpgvExL+9FXfwW72iF1n7evyaktG2/BLpC2GKFkmKfvKh
jrwC0c6AhROZgOAP/X/qeyevlDqu13xwFckTu8UokRtTcNMeN6x/uCq5bpzc1uYr/kM/ng8g2j/F
IulEIXE5Y44iLFb0o6ubH3gtEhfeAbUnAqeDhKh8Az4A2Nz/BDu0JriChPXrPKPCsaZDVlUYE1r6
tb52qnpSIRANtqzTx4hb7DwiPE8BWb4uIcAllru7pQF2rnL9GG+UjUjXHzOB5jzWXmpW5AkqOaq9
tMSrFgGrwKkOxcq7Mw9HLft9JFwCijm0sEtsLZJ6NNl3Z35EkdvDahWoGMuECYWxBeEeXOO/lCZX
UCgCII0jW5CmD2RB51/3QBtlrCPa7gDeqWRbqDmTJUdZi2bVvw8w7LKdwppequVl5bm2lRTvNb1g
vhgO9IhhD+NMN+uv6ePDaREmO1jG5r7EGaEJBNAG0gqLf2+N1GG6qBq5GrclFtKpnLrL6CpcxwLG
YbDgrVw3Gi6PMplkAOJ4oz0gGGFOVmJIe6KOCtA0tnKjaf7kKFJGOoR1fDKfUuIjMy1GLRR7ZZ7z
lS1DvVpR3aGXT8y0KPDKupdFqh/XdRhIesiHtWEQko22Zu/nTbg8CDZ3s4dO3YtVmnn5tZR/AxO1
rHjV9lLzFj/49embjsORk0pyl6L3xUZ7dypXJUiB8sjRgAevhNbLXvu89qsbyjZFYzcNccV7tsQD
MjFJdave4A2n9MfHp9VoiDfjYcEH9yJoBYk04Z0qm0Xq2lt5lKAJ5Kh5gMTPC6IfhcCAsDvSgG4h
Ev9P91rXUQsXn2yRG5G7RbOftPYlra5H0RHNMipXmWnlArxqvMIHWJB8buZSK2vP3xlQFG6SWV6B
OCCVFoexy2lpOEL3uwV06YptuSgjbE+smbTidWLmiTspyrkUBZRDoNjlE/1/TtWmyur86V6c+JUp
pPoY00anzzek1qdqBcM1QkEfdbaAnURFt5rBq0RiE4/v62YfTKJNMoHQkWmh2TQObkpiaX85uvva
8wqRuGb+yKhxCzHKy6Bj1S0vZY2c+Mh91gW+koLYAWWDwHKCuzCKIY9/18svWZSFIuLcqUjexfqW
qb4nSX6KIO5YkGTwKYJur3gN27q0RXoT0TlaRdzXVLwqQqr8Dx7aLLChjXYvqL7g/d9ci0t1CuZX
7BwkNyMuRVr7z+p7YG95TSrnN4are6ynSBpR9tVCCyGotEBqnAy4pEEt85V3LH5yeOceBvnJSlq6
r5YthgTh8Xw81euSbXipRPHPnjloGUieTZ0AHnMKeTQdA4dC6ABqlhDbexmlkAJ/rXTk+AiNlakM
x8fgrQSVG+eVVB8F9LI78cMukdf2bShmjzMbUcufNCxPaOU9WDpeWCqkd6Vh5ZSMu+Vh3xp/es3W
m+uR0NJ9DURbEQ6kwNh1MII7nJrD5bj8ZgAqKiUOv58IfZTZKqhXrC5dL1EkIKh4Tf7X2IDZHJJH
mDgyEZABYNFv4XHrsKqyNJ4BpdZLRHtODyLomD93R+W0kYSO5R5mtOW23c75dP3Hw4woIa805rB3
VkyqijYcBSyL+NMOs3v0wrJzY9qGmZFwK244EPq/KvbHWI1GLp8I/GbicbTnm/R/vGtcyI+9hg4R
dAM0ZCmc6p4AKn3PRsso34B85XbAY4HuSBVdqk39jkvrkHJn7LIHGR8+dh6TqCNxcvSJOryZYDz3
AHpNr/ky4M1WXHpBOTEbQGQLOHRTrbEAWFyHJnqpnt0ApwY1je4pYS2LTRdzxiy5+X5QKpa7rri2
Tb1XN2ZjVjshbjI44HLRxjAiw3uESPn3OiUqcmQhWvWiGxhg74MYzkBN6bbrUX+DEI16iyzHoqmN
k4N3p0FC4fHLJNjs6EppnJHsbOD13hevhunba5gTZ6+j47DOsV4QEKnDnyyVmZ3bS5iURQtSmfjn
/Cbn4rOcJ3JIYNog8X+CFZIQz+nYOaKZutfN4q7kYaKSQVotT6vS/FEYtS/Asacp6LVH6W4kGWXS
U/fQRHL43tGTsykH/XZWLVX3lWB+2u7+sUlY7rJ5fQBDy3xeStQ8qjR+5U6YAFmvAD6F0COIKEoM
YpdGzyUwC2X56zmKNKRHCLqjnvgBu1kypEYuAptWckmA8FjRL43avqyhBpYuirDOuJOwqKMNOBWn
fEJxEkErShrQr4iUxV+ZfGbttjUiaLgUcBvCC/rCr+gNqFK9O/y93mXG/OiGXwhxn030x1wjHnE7
A62CmRVDnu3KH9vvVOLAuYc+HeCCsPVM5O+447A3mj82hkknGVcPFHHnAv8NnskMwfuHtzHJ1D+o
mwWzXPkooT7A6JeIAKsIZsJXD26sXgs59szJWUknTQHN48Ewxopkw9S5J6N/YxfTmBhRnEFEjzd4
nSWG6VN65W5vq7U5Ji/3ywtiZx/tYTVrLQNWkqxZsXhg40egwgG6kNK37yQvva7cR2GdMGhETi1i
5nxYtxNyE1IDfVvok7SvjXa2cf/C4x7lzg3hxgJZGlUr/YQ+94ud2BbL/OPEh1W7W1ReMJZmytUc
kcOCQ5Zup9sSG0PJsv1KtP7i32XsuWrHBKD1upn8Kh1X8vcCRKMMCghksXNF0Z0WQEJteO2qGu5H
rgtL71SStlMnGt3krdsU37Bzn11RX1Nms2qqHtRPS+MJ3EfCcshC23Df6XjH1CcTH9BUxsl4WEy9
1FewoAgRdzOaUMhz9MQGORgexOqrUIouk8hBUzfCkLrngprdaFyeH9H86CXPbrPsOzg+Oyau9dfI
DFR/PXPSEimE19Gv5VT/Ds4UkztDGU5r28Ckv5vsVzAt6V9qEnN6Ztf31m2QbRLfwtWO2xHu2PC+
YhMBnUvXmk8SPn3dSQ2/2Cu5YqFX1HZj3pokuilo/npZSuTlZ4wutdMAlCofGmwWmBZSsIarD/hf
4/ki0KTaejD1Qjhft3LaBnVRbZ1zZoERFk/zM4EtkEKBJUSnBSZOHk4Mg6SLY8CNHIQ8hrZF3w2A
yi4IDj2ZAftIoe0ePCE4NWlatBMUpJJ2aOCNmqNsFaObFQXSqE9eF3R8Lx+uLxzfnr/l9QwHcV+A
g0uHeDWbKLTHqh2CQJFE89NE7VN3PyvjdFSqnJxMoXIgvK+1PBTkq24Vjcs6IaiCxLwJLzVsbVlV
w9nB8v0Ex35IB7WbKQB6gTHL4tebRCLB1ZnC+RE9z/XnggtGCU8Ah2ykGlmFBv7hWEwPFLPgbahk
OmrSkARMwp2qKxVJXAezYWKeLZxEqp+SFYCZROF0KcdFSTulzUhB3QHtq2Dr2XKDs2MRPUHV2AcW
TJ0eO9cnyDoZoyibjVfCrqVKDB9EU2CRDuh/7VsN7xPtotjvurKcR8id93Wfq0TdZl5LBIma6Y/U
RV2omeSdcokuQJCfUCzJ3dwj/984AlVhMR+QKCRp4ZPF/gZkuU7gDPJ/RURGXc6YwoJ34f1HVhdA
C8vK/5OktYy0qlHE47iwIoNtUbIv90hoU4n7q3ZRBHYgVKEoqFuqheHQPOsLgzVrr++0n3BlDRxG
xpNg+LRF/VO8DzafdgMK9RihgVGzxMPV3RKqLiJfuEIdpXmyVmZq8ovUjZOIdSkyvY4Pi9OVMm7L
/fNIqRvC9JFNUTXB7j7sxCC0xdNBxU6LQ5/yUc+cITP1FMZwNeNy+hRKMQSpNvkcexkt9rEm6vSo
fPudiRWkhxtZQ0x9iz5qDQxBM5pdMx7+PnBIgKYbTakar0cGBhH4SnHtZAkOXQjywDLFUI54Rs3I
LheBItfNKh/KZuDuy2JfuAjUyh1aAUMBmDrrDgTfyPf9nH0m2MmtWW1euuR6MnbjQlPN+U5qM1m6
TvnuMHoAwxrfrYDeGx+ymSaj60djHszwWW1sEFXhVYaEq1by2AlyP4lt8wZTXCOO1+NOaz+SO+61
1K0wPgmoyu2WB8FdhChwLtjj8+tl/KIEpmH+va4KWIuikF3nIuKi6aCKvAFD5v/WGDF9+ZNKt25X
sab0d1fpxkNdKYi6ltSrfcZyWxt0G8iqys+3aTJn1Fh7AGVCVxmXf5xjHis5mxYmnLUQCM2msN+i
w9bAJHBVbnvGIsnOp8aL84DquzUtqOqRT5p3RevbccJteaxtCrqLttQE+8iE1bcf8VxRXzG4ojkx
EILypPN0pLVFH9y5sO63UK0077pdndFqwoLBcM4eB5X2XuUWsGawGbTt9PwKlc1/oHXxO0EXiMqq
b7rIsycDZxilrNqJZejq1qt3M3F+PTWFg1/rN8nKsgtpebIN4pRLtMI/x/5qdhAA8D0g3KlG8JLb
5Aj55epEXvZrIUopndb6T6v4d4S6yCVPZnO1dURQSnnqPzD5zW8deHb2JlvkW8YVrrzO4rXRYsIh
PrxKRxFaPRbm47g5cJeIEAXkRLNBl3yrNQ3DI/OsjaIGTeqqsxIPxx3EejMCNN/XK/s3tsS1el07
2KHp08T3+eS85AaohTF5MTs8Qq2JEtsbIVTgcGRd2oJ7pP5+NnGkI0d6kNiMLZpLYv0BzhgWJHEM
rf8R1uovEhWZ/4DNs6O4V+rN87X3Dfwu8RyiRXAmNoOnLllZBk13sPArGEfrheWVm/dCdgXiu3kb
b0OYpJrV/LhcxZgHtDei3yQv7R1Adp0Py4iECXRtFcl/8m32kR91rWeQEX+cna8LZYcm7liyb8Nb
R+ycHq2t0tp8O3/KbbpJvAPdLH4FpUrRkrHvoAt3MI3ax2OckKbV0rPRTg+cID2CCzTs509U4ldV
Y4+2cX8vlNqDh6dBjNGchrQsS4E2/GdB2u+gUeVWI5SxE3P+DzNdjd57T3odcZ9td74AYKHlLo8F
qhPf1VJ7dYYZziDKDt939EBTM7nN+VFkWEGgB3ReXmDFXQA3Qe605rOeRD4IjZSZeTJ+9LYLO8fM
0/z1NS1KkZV/5vBSXsHBK7I1FrWZG4CoT48mkyCm0V/JMxc6+dD77EzEI6+OQmR58tlsvcYhkOuX
IvswnphP+0oWz6N8UrWcKqyf6us4aouMIt4KZKXoCv2GCpjkuOc9+KW9PSOjU7aZVQvDyR2H+Ica
PWr2Ega4JwXTmvccEB+E0DpM8C3FO/8V1qcTIc3Fbkv5dqGLMMvJOJ+BG6wxsKNQxI8Nns/4UHMe
A8tp/Tsymwd4kJUy702UGvYexjPu5JsxDvqA2LQ/9tUNZhZv7ZQDvcrRBXuQJaYvPdr6q45cFRV/
tlNnmEC5tliTtF+OphAMKBRKiDJWiqKwkjXyh80fPs3EAHrtJbFec1h/snYv+nukbuIx/SEdFG6A
VbTfOTPAk4yTdhcbmcAoldhTHEZ27OvSKLzXouOtcoclbxeoROicLlWsaabA2946WvfaRSlmA+1M
doaDMIICQgUKdo4EXbEKut7vV4oU5VsjihoepGDMybsTLJw82xVog7NN1fTBkpda3WEuEfCrya7g
LHeUojGX99XKIGQHJdVtzisHTjaQg69ybYi9Uy44tsPpiZl8aQc8F4srL4MwZHaqXX6M53MG/gp7
vYzL9H1KKtRRrlJ6+PD4NibPPDsvDO10ZJzPDuR3gXbAZ68WOB2ZhOnvEkQL62hGab2MuJl3L0Zg
KtOwpal8E+op3MN8KBDhravUi/Nt5Gw35FlifmaPBjg2byrrXYOqUwz8ZF7faDkYDbRUyrSxMwjY
swBVJowjIy/vHOztxk6h/yFvBSNTy7a8t1GfiSjieqr43UKiJU46qfWpzl2MFh26AIXHRqt3pj2x
ztgT+CVI5oIxaI61G0/4lHvaGNhmBSki8YJngx6QrDrPsoACV/f/Ncnnu6pHYRoTeMwfAm77tdV9
Qrm/m8qdhC3JrBtOnUZXfLLcbS70BiHLmZ7AEMuluwNkKE39mXeA6ompBIMmPzCxAil6KEdr9INz
rTjdk1AFvV+0oSdA2GEKvDjhDYlqkWcA1BolSeRmnwitpD3YsGSigPTjz28OWk/fpoAdEvF3hEO7
H/aIK9KI5pLUqhu6bH9FQVuV3ZZwqtmwPEfnrbAA/6R0xf4M6EbNRfJ5OBJVNJkwjBz49XDooU9u
N2aAVA+7JTx7Xa4UYjkGVzTzPZDDr4ZyOi48X907TNDU9cvEZTLSzdeBjWyu8JTJT15Bla+yVT+0
7rIPLLtpB1lSzwkLpVJgdfvojWSCdf5dkuHNO+qRZBM249uxOrkmdPDuf3nOhaSa73Oq+6vZ9IkI
6u2gyqlj1Xo8YVugTfk22+X82mojcSCQQluODP7/5yB7GHXCBLjEo5CHKhgtZS5McXWZO8ciox9M
2XixJIN47WBI1lbFg2DDzROE6inTFi1wcB2dT86n+iSSD90ngXKeqcwGeSr/HliD2AsHXQ6jz3mT
uoSN0wtI9CHVZ+NfWKyggJh0AMBHwpwQs8RG4tBn5ISl5TnoRxTuPd32Bu0wq6ib5LMgi8l3xNUK
Js+4fFU9lBsS+yv143A0HwBEpd0BOBz83Ng6UhFNs8kzRL9ImYU/hUZkJ9WTm+tveHPAwlq/bLrp
ePbU+tQZad8lueLrIzUKh8x4VczNQv6Xyw49vLokz7dw/wWEoHdsi8TJ2E9Mk+WZpf58qGkllXJR
6wpkv3m3I6Nr7vIYdJvqApl1HOCM171S5B51xMRzmPI1Wj5DLse2pLsH9WLsp/33A63LtPevAhuA
MAtVaNGm1AGuE6wVhs2yJz3kK+w2Ce2VyBz4og+tY+5/fPKvdVurFZkzBJeQNgWD1wyCMxGCN+yP
S0yDoXMlbhi/c8av+tTQyvNZj3KfYxsBd6B6KVrgEBB605bn6NhjC/yJhiiYfDxcyqsuv4UmXkZD
0vTfUDulxSeBU0iFo+LF2jiDsqZQwYRJ/MUn9h2MP+8Vu/M3LF/nHpmrNL6cDvp7zCfmSGJbmRw9
pGgl+3UHkOD96HMRQTo3kNsOMM+h90482UHwFxrNVNaoJvb9fPUIcoeVeeUfpmNvz0ik+++Lkhnb
l7AH4zZNKEj1VUbMQYnQNKDfwZe5RNE4I3ekHau7K09fMK3AesEbKmNy896ZuwjdzHjTz7kIJXE+
XkikuiGY6MxMYT79+YyEoLmi7pYJnNvfMG5aiJQcqxC3KXEsXhgWdYy5gYudhtFWkUhMxGwfAhs6
tm30DXnwe/8xOoEH1HpjSbstI5+QpVH5v4DujsxPINwsKhbOUFvoKscinHBr328qcow56GpiQqBz
2C+9YiDnTbADRDOo2waurT+Rvoy8nZ1H/AqTuA9yhUP/vr/qNZwzXxTb+zBp6Z3Ih+XUxudItLFY
nHDgZHdzKNFtF0wXQ7fyxun2ZcSN0rOkxd+jirODv+VsoLJOHBc/iv96pOUTEkDGOFQGMg8O2H+y
ORYJwxaEj1lWpmF4PwBG99hc1QTymxj2kVzZ1Rq1oKS6IVJjQq8nOPB1J4TU0v2eBPvevmdu0mKc
P+sRscP6TrHx0HLeFKVY85Z3/VMa/aZc6r9rkO+fr9uYRDvAqevwRglar+1zZzOhrJyh9lLna0ge
SET/jXU/Z1tomItWzsIuW+0xoaX9Sh+4StobsylQDsQ/k8GPW4V1Pt2QO2yd9sgaK3AtwMkqT7Fk
7RyMp5Ck1aVRwyCHY/Ho46CiBHdZtE3gPiDL+xIuftskxlDka4C9BoPZM/fvHlmlRgmJcsHhMCM0
r0BFDIAyno9MmRLzIL1FdPLmTqqns5Mdv7MiwT9U3j/Boh5Gf4BWgOH2sldMwMwaNnMkzq1JvmtO
d2sw4WR0WBuzQByvEUV1Gv31gs7Blx8mR2V4SGaXqLCr8o6/GV9s8kCrOyR3bB7/hGHoJ/Fknfw0
zzyEOa64A/j3EB1FwN7XKHeddrxnRilRe+dLQCXQYIO0dmVt64PZQGbmTBD86Pr8odsG4yoemAfU
wZPVA9W+tDs1/nqnErof5swevKbxDmYoLerG3/fiXEArATXkIxZ6ZB7JcEhtQupsE7C/7c3nzw0y
ONjK7BhG5AQd+21HGXFwE+MO90feY5Ae1yv3MkoFCJtsG/a6r9lmmOkc29Sj8Hn8u7XyfiwUczfl
jdThyo7BU0/YKWZ8GTXfoK0D6y7EKM59yRFv+jcfm/FOXL7abQ25ujFmYmA0X3G/Ku0DN1oWy07+
DsdxCD8QGG0s0KyRc0ndZRb6i737LjL9n5zF/8k30RMJP5O66z4pzYrQdNgEtCncORMrhNagZSgM
cArR8PhW1uojt/XM115IajOY/aQSpRc/JknfHsGol8oV9KU5IteRTJcQ7sGxSnr6Mm1mJRyIpyKo
dZy8OoR/3sEe1OTI139PkI2s2clGzfcSHUcIY4eiryuoQK5vfEMsQhljL7/p54yXfIbq0Gxl+vlf
JG8dQkAw2UM+AIahi+9hQaCsV/3q255stOTgQ/CxS+guiTLJnWUChbiAsSQJuPQDKeSC90mxbNXZ
41N4W73yPP8l4RxVPNEJzOFA07i5oiYYfCoOujeJALg1/ijkr4YM0LRepnk3aaokX7u3vrxohWx2
cVdIdRUMomG4PfI9wWXufXCsk3NclOoYikXvMziC+CeosBdlY2XyxU8ievxPD82VQFdU7LzmtErw
jv2pU2XNY59nw3Ite/lReRWspz3ssDF+3HWfvWZO6tQvs5uD3enLn0cAf8s1K/iPc6bWReKSK6FP
rhQQLNE0emEf5J4lCyEiVzb265D4ebTLVNgdjG1OYOZTrtvVmYZvYLE1H1LtA/TTpMAAlT0Sjpte
9PvVEvDfDMZjrmwgzY6kbba10ZuxhayNuHDTtgK2dNK4YJU9X00ceGuLn5/fJhs9IWx84VhGOuTB
C51HsFEQS/ZENKxceC7gOHbV+uUhQrMNPtjUh2Qh7nvDTXGzIEEcB4eGTkgZTZzPBXCrxrGUnvb1
iqAZYAEYWAjOioJFrs2n3sUqCFydX/AGCClNI7oOarCZ3VtyhWEnKcXS46/fvDw3/TWhM7aZXewQ
s5ycDgeikIRsWHJJ/Zkqkxn+8Z7S+3YYWzjEhkVC86binpxqKsotM9hjCF2lHE22leiKQ14g9yn3
L2VQxukZwGRfN3l7idz4/FcizhXWJbemMQZ5n/adt9m2+Gql5Mn8NCFC/aWkMLEUiXHVDdG+C4BN
vDu8TkHd7RQoXT7MAm6LX5+ptlpMjwzxdcOW4K4XqY0PT9MaDDeWitn4Os5wr66/GRwS+EF3t7eE
RWZAg7khMvoM9wxLTJp0SgxIr6Ui1WVSCWw24LnBdK8HyaeTs0BLW8ebFjyIQbUWVrLPGQQ6lCRh
QNGncsLbilmnpV+wgF7xUhbnrDqxmx7r/2MbPZKEpOQUuRYHYexuj+HUKi+FJQ4wpirnZGpSkhI/
DnA3jiyNYR9Dg5B5AjZcklPsxCtFHAX0PDdogOt9Qj8y+an8NJGuugNf3yYiuvFDaphfoSmNsi2+
oaDD+hzi9pszCzql8rdM2bxFagDmmbP8kRC4bBSUKKrK9NyxQ8rTOxkLzi3siUbFjglQ5tLS93rL
MGMTXyJ1v2flodhQbhk6XaAIRFtI7IBoa2P76Ky/jQ52/x1VZ32OA67f7d6Jhq2HpXclfnHSaQvj
p1OV5402Uehel7owGGcKZczhGc1qwitTfAmfyxL2aLz6Zkv/FlyMJ/FfnWvR2Q6S22IgTmezZkI7
H8L50LtbyYHD51hP8Vn9i51nYR2PgTirx/NTF/ODzTAySswVsKBmvSUEzOvT0ZNPhOo4rA16vUcY
LXJpq+/gdvB7cCgIAJ+iitDloP92+ekNcs9Iv9VHDS+Ll3eeh8koNGsxnYDuHs9JWc9uEk8p/YQY
50L0jJ9AAioIT2/Ey+jLAilGpHRBy2gllMmBdhaTrRyv9AfQ8Zg/VDjcCrewDu0MoCCaW27HdL7A
YTLb8T6QzLtTTz4VuoA88Ci9+bBYInHgg5fTYoNFQOPWtE7NyQbIL+6SFSAsRK/vZZGmj01yj60S
A/KuUVRQYVAMV45Xu0A3s79/cK8JwKVRsloc415ULCoZZhJHnEyVoWrWK8qxihh7LJG6Wk/vZHK5
2u2YT7VBmGLSQHffPSKXj6kW+QD1SIMS8uEqpgg5ixt7d4c25aP1y7S/qUPw9bFf6zU3V2LBlUKc
t7W14q+KXB0kYDPkXgbAiNkqAhCcFPlBBRuYhDMF5ezW7+2BejYJnZE49aSGr1XEBZUH8b0NeZgf
egzM6osILq6V3MtS59hyTYT3dEFOxz5uFlhoLZiDXdQAJmKp4myyxK0NcAc+y/IXZkv3eGjHSGu8
NZE7xyuh5ERXdA95x/pQVrnj6qITXlaqtUlc8JgAe8j4xp/fxZ4E4hJfkcKYHKznYRKtfZLQCVUj
8DWMQIsqsUhiQsPMV4K6R+XTsIaXmzzt8CWZaO4enjcN0pR4quTCpAd0lAagv42yrorIKkMhc8Cl
oJgi0WhnkL7/L0DoX7fQd538gaqPIylsEnaLEd3AXH9CGn6BKooQFtjF1bKXaRCcbrx9N+bhduBV
5ig+yzIqTlnc1LcDCYCgQFiwzmemZfRZm7pTo3eOc+nbLq35baeUc5TfRcXhYux/icCcfwYjBR3A
xFaAlfPz48QjwT8eOBKrz4pwVOvwJO2R84bilFpN96aGDZPUtL0aGkTQPhBuDDnBeSHLtaza/Lxh
wHs21FqKWmQPT533MYFHozNj7ZQ4V94ZXbzGSXUKmowGn3XvsNkXVjUhZRlqFjp0gRpI2FlaxQEB
xZs8nCNsFuudMH9a/uZV+qv2S66TCctyhvzx3ArdE53v0jdtMkyHEb8kvta2k3uUIZyr7SOCa86y
TIPhrblfMMWPGkvl9gAAqWZYCw2ZvxYt1WYNPDTsXTQsd3f1cLNxsmIcWqlz49yBCG6Kx330e8Z+
aUtjnE3fz7SMl5lXqe1wTXUnonPMyXe2yaQR+5vRrAODv4XTb7hfYMHfyUIKRZErzp4M9VwXnqDK
yJZowUVuh7BAYRVUO0VE0Ug57bFbK54UsnIISTbMimq091oa29qyrC6Tmrh47X6GGaJ/HqZNsyPe
lT/A4gurH1QJD5Ukg0QLZEilJVA3xbA7APbO5/tgaSzo6JOwUVpDW2CN4CKIAOw1LJj1mXeDANnU
UNOV1ydEp3jbdl+V8NzHjHQ77p0FA5a4XHdaN6gDYyAsijKNWYfOkaKMYyHcZ1RgI58yN4VuLRZC
w8rsLuFrwVAVueZEHdDA9ncQhrzn/HfYFW4bzXx9oKYXD730mZCEmNeS80lpr8QBGthwdc7Vysg+
tx8xNVg5+2C7NCifFwbHFTh0Rk0OPeqEcaIavOVPpiYclqRlhwmCYKPycyckvzQNa9vwham8gb7g
MOFqV2pa7sED/KMRRuZUcu3NExq+jCwlUp5bi3gmtb7J5CCVggK95FM+ZXDZl7Ql1zAy4SATlzYH
orfPVQnI1f6UWdcF7Bpmd784F5S80wTZRVbFEbQmQ4FN+LmETaMxlv4NZsNgWujUeokrYnS7FafE
2BVxjzxFHsCqcn9RcBrI8d7wVJ3JrbOurEzhAujoMXJTSsOm4tzr6ClhpyYE28ySzfGalxIbWJ8Y
fHDaa6CkfgWkvEZJp3upfAhHFeFNwMuP8SP38SmmqXUxFijVo4afXaOdkuMgK4xgeUxD51Gw99B6
7RMWmTVJeJp4LmsAzO0K0Q7bjucgVht6f52esp7zqO89ZudeWCnlPYJZNt5ZRsOxyJMvKsLK1Lk5
infvGnYnknCbJMHYskRunYi4oa9fyNbKMtkw1Yl0YrTIjc3YOjZjX+7RAyL/v/4pbu1XzSd23/vO
RZYQHADQa49xw0DPv2zFGTkObaXQrVwWrc3fHtPedXHwDnuY5MqknZSvm6oynlxsBUiC0n/5S3hA
NO8IKTBTyd76ozkAOfiS2fs4J/Rh8k//yEdtnFGWamtRUtk5lDd/jBqlsyyjHUGUtvXGetj61czv
xYFlT89Q3y3XCL9iRP6+ZbhT1qfF+DiMBx6Ds4LBpwttzO94vBvkyvVLYWsAdvJp1x1gRezoJITS
a7r2EddrEbxdRgKsxzHM5L9/zjLXZRc9YaNEk8tgS2zdCqL+Pd6C+ej1k+e5Z+HwSeT3DuHw2VRB
EmYMe/REYvH/bOrL9oD1TI/iWr7j0GA1s4lhlOhf7S9w5jKMEm+lsB1xRYoeC4bosL44/otIe5tk
uUYwiMzVwYAS4PcvXi7CneQWjo2DIRe975vxNqa0FTz7fpedDWRV7W2slreXvzmoo+qKWv94gPnC
hirOIPfdFs7Ht0Ix5RVXNZc7FmHl0Q/vgsp8lEKgmPSBbBtrqUOi8OWCNQBgglAK2Y/VxVxOf1tQ
sFKql6+tRVBZIMt2vBM733GCDR4fss3727dNc/uW0/6u9UJh6DKaG4AGdbFNK1JdzmKmpuaCC8l2
BE2Y0Vw4bR8TYejw4HucJWLFkjLYrRdoa+Itxi2rmZ+IhPl2NEWdV23Pbm61pti6pPby9zsjaHCp
I6CJvprxNIWDPj/v+mHZvgraGtCzygVxAlv3Bfae1sL3M/mRRYn+vCm02DsywDP3xhfdnvMP4S6Q
35LtRm/FrSpmTnI2EEVqpx3ppavI/HVcerFuFQhzhagQ0S1Hmw+25c6eF3FT6eNtGP1cAU2IMTlp
zOPk3dhxoiyml/LNtsB+30/rL4TRXTo96bYPdkvQUraZTlkbNnjhDILniDX6rAUTCJJ40wARHPAz
WuDDJ0gj9ye/GBy0lqirdyiwZ2/suUvQNQ3Ch0mJtlYiUT+ICc0P6BkQCUQe36/+dAdmkmVVInlm
81NgsstQ7qRy0NdJxCMVz7Ns4uaR+4+RKO0XXYDhrrBFW+aUhG4BXHYG5w/H5QL4QD/7a3XKrsj/
iyEtTZijH7Wwf3kJ6UkVKuWRUdrOXZBMBYJX7inLPSLER75PhutqmuOsNcSTEYrE1s+eSF40ipjc
CWg9YJ6+fJp5FS65AZunkAe1wVl6hP14J5X4hYu3gx3avHgeViTvP4PSdU6hlKesgsrI3UeNpnZq
GystjUWtKquqv5cmXw2oczp1s1+9vvMNXn4dIgVsLhXHJM9Cvbkhzl22iepssAc9qmPXP4ZKI7J5
GQD54fj1zYGRuZWgkXSmYIb0UKAeWSb8cAL7THa3C+qFVsh5pbaoaLHRXiYJQ9y6Waw2fs2ammyK
FG88lM89jc4l/eJUfTG4/0Bwj73zOhdwD/+YlV/aIqe9OwWI1WCDnVjt5/tjRSLw2vBBBLsj+mMl
0j3qo7DBsYaRAUlHD6IditVo9zbupMGCx5jVZGgLMYSTzZKR7zyhBhm/aIdB7yYS9VqcpS/lj9+h
9SOi2slz99VTLWhp5WLZazfwwrXM7z7aot7YoN/KOeQsDceinFGMxiJR/kcB/8h3+GqPhKCyAfh9
/Pf76JP8TeBRGYpAvCqiZnAamzbV7ZLMkKyrGQELGwSty2KKMAvjkWEMlKMPw3wYiJf7AKBmErma
2fypydzEXSXKYOa+kuEUZiUDsAPHyYZ4rPeKG/o43NosQbGr3AWTZIjz/Lbiql38V5UFrabBsM7q
XmfMPhuegB+2vuFDpId9KceLHenrYBsIQUH7AQf7p+sf9bg4U5g8zkTMg/mW4H0YV5JPIa5/1W7S
vq/xjzkeMnO5bY/KAmiPoLYHbcK6HwgoT343jVqdu0L3nEigH6jvQemSjI7q9MdGQH5N6er9R4ba
KKlbbzO20xgH6iTKV7sF0C+eQTjpuDxfe+SNCH9DsFPc6lbni5Lds5H6orxXm7aZ/VksUx/2XiAc
9xXwzdyw/HK5ydBbxbxMzxp836scWoFPsbMmcZhyFd9zuOT8qZqmpyfksnGYh/LcMwmK4pj7Gzlv
1tu8LQCeEmPolfHcdXzniWOuS+8dyaJKczq+SSVQIJEgDmKGHv8KAV1tcwvOQCCbjNgjIkjr0uUU
jrxHEoNiOBMwFztgIR0KzPpkmjfsP1TvedHqtD/h82xw72RPDzQA0mlr+YLmaWs9sqxvIYB0DUDz
wl1Xy3wC3isEexCGhfjD3v7FFIbQQYqEF60oAQkEf41Nong+gS4Lf/lNotFfk1M9pekP/iWKSzkY
9InagV416joiivAxE8xsfRJsJzr8BSmPUOU4QabO9Az32bRNXkevP3kmFbqiI8Uv1tW6KVwXqkNf
qK2rUG9zM7m44e4xiEGlQIt/WqiEdYnzsPdxg4L9onUhDHuOFkned2Sk11QaddQPRrr/M8D300DH
Zu7kSvBplVdkl8cvzzYGsYOWA+xlA0bdwFJzu7OSIa6dZRQuqQlEb1ccq+7RT5qmTWmCsiTwiumY
m0krA2VYnVZe/553fm8Te1XOCCaIkvxZrI99z2jS1Ojx0B6xTCXAGc90k3vihSaa3BKG6B9dSokR
XDDQVqGpYcLvw2MLleiIMLVBGyfIpeK/r/rvYnudYGcgJHdszLEEjH7khiBiy9Dtt6bqK6vzyrc0
DOqqgM+G9l2FtTxGCfRUUUjCq0Q9jMtipvaPJilo+7vzmPmkl6NKMP/2rA6CMwalSh9hCpogDaF6
L9IMENOwSzgClkWX1BC/lTHaP5q4MuUEuuQHm2MkLT958dAQSpzIr41IfxwXV1z7b5kh0Owchsmg
uDW7DyNNTaK20oTL6QeHkOU1M0zD8c4HQQrngF/DiRsWSSXmBMfPliHuIK53s55T1L1SyZmkGvC7
nkgRCp0VYfLdwO9VbYd6Qf3J+X/1mOHqMhSsbKoJWleJX9YZL94dswj7nfot3YSCuwNtbTvF8FoC
qgz3YBsoraFd/RgfvWWkF4cWIZfeOYQJhnYDdaAUOfh+usLFqceEIw1IHzenq6zp5+6GhpvsTQov
Tt4Z1g8wX1q1y+ASAObRemqOcUSoWFY6cndw8msKltLU882O8tS3pQttmYo4kIYHFxOb0SqrqTlV
yt77o/9F69OdOmGAUjE6o+IqcrZFiUSwDf0O8MWaThIWH3UjDdAyNkn0PfgIqeu0z+qC9Dsv0dDQ
kk4EQx6hEuzYL7slT679QrB40vCanFpBs+mvhA6YzSZsq3154plmYdPFD9jhYfK3JTt+49fgIjP3
iRyCBb4tGoYMGEozmBWUy/5kiwnQdC57BUHJKxAMwy6Ynh1OfkBNSRu7wSnI6KbFdjul1Fw21Zby
+01U8PoZTxIAtL3vofEWM4uWF+mzPrS2eRBd2FQCmdursyNhzD5k09JtxqK/JR9eMLDUUv2deQEo
rQiQzvv6O2PSS5KLlvAC58inBLJCEJmg1r04L+R9a06n5mbat4yC24UquoZUcfIuYB/aYyv9v/dG
+r2lGXJrT29qVftITDl1VLcv9UVTmx60Hw8wZkwXuN+FQS3VLR3WNP/QnJlDo6lJJmUAgPEj0G+K
NWJnRV8mK7NBaxwwDsr1obDRww3DQ0KvXghDEutAOYPt49ritw3ycwFySzOCQHm2hxT6ajSTJiGU
BfvjOg2NQ38I9ECpFvvqwmhrf6MHy0aScrtYhIaOVJRgo/rcmP2FVqURqqGYsWQa8JOBJIw4jjVR
PgAPd/A/hBLwfYBhEm/mWvKo7XXT2YpaHkP9YMAJ0jH8DLyBxVzsf5ZlDF1s3pLUHLiPTu8rYGVu
EJ/gkm6qs2UbQunwj06CD96K6xMuulNTlbzQExwgeHnjUppgXPYZhor/pjPFfRZoepGXsIcND0PY
vA0bgd7zzs+7TBFfr6C5rD+waaWU8LzEi73yCOVBgwZIcjNoZcQg0a9t66zj6qr8tGI5soPrBTDs
/ivHfmPt9rCNcYIzvdjKy3FNPvNZjKsBggrZc43j4Dh2qrDiBD7vUhvf/vHZk4Um8iM3Fcm14s3u
wal2tkZE2ZAyUWzlsHoUh9alK+FU7pe3VWoIDPo2m+Tn0XWwKsChX0P0Zky6scHPbmuIkFeVQVVV
h7My3y5h0u8MZ8kgM0pUa9bH/XsrgP+A1kEsH9k7p1vCCw5iMjLXx4kIycO0bdhdmN+4IopAAjT8
/ugiZ6kLHw4vePtQAt07GxqT/m+jTghU1dTssyO2k8F3D87X+MMPowlamC1vqoS+qEtM59WqFwGZ
nDGzDk0/0+DTkBcxS0wpqDqZNOndJBenBTw40/MK9xTQ6Ly6HskFtz5NdUXeL6JLoN1EH7UtDPbD
VsGqpD+fmCckKi8zNwCSw+BgRxuWoksaj14DTU2Ic/QGA323Rd7AKXxMmYz3EmjqlvSJMIbVAmt3
i8ISKh0o0QHVFA+0NJsO+zNBTxWMp7SCJgN9K9oP9MWssGXR3n4F7tP93YN1LEkZCt9zKfURk2rW
G8dWpmIKDv4ZHbyHrWCgjw05xSsgiJd0EOKqPX9o62/5R2R5GhIDqCHmGl5wx0pqU3eIjV5r7yJQ
M7dydiNTblx4JJ65SRw5WCkWxRb3aElOTkAjyUM6fk6j6Iz/7f109WU+HCLAoW0LY4oJDaeNdtEA
SAvRhyxz1nCO9CzpldRDU8+F6iasI+OJpzuYHJ+/0Zyk2m0uuOQYq9zHhlt/4PsBwJ0/pilTOKCS
lSyNCvHIoyBEHL4+l0KMyrH7p83ST78HrSWBMBGhqSDY+Zuaq+8pWWsI0zTCYcIu9ISovaAWjGvG
HvLq4LT0saGfZsKKu5s3RxQvn268TYUDzqDLqV+OEtFqOqyy1w06qlKCHrQApM78Uqu0VPoyiCL7
pLT9wh/5NcsfIEy86bW7GUlDtWocotOSqoU4kzzqLHYhQCJjfuhNkGapg+xpBBzcMIPgw2cb25qL
cWxPbXLSpGoih2mg51Yg/gV5WJ+RMcdxFuKtJvmaLGDSt/9CY1hdNJYJEcw6TsxajTDdtD1W3Xoi
ufsmLBhm7ltInjpUzoRkNYaTUzMc5ItBQxjNuVTZkPlNh6rBEoheiDzJzEAuTeWtDvSLwAyh8hhd
KUGlyvp/u4d/DMyd4JmEFm4ZAYorw+WH+MDJ5ulrThBUTmFtYAgJreIFpHje/w/92TZC5tA3BLqw
pgD0PX29We5ngC0OtXML92xifw8sqxMRRgqdm0WiJMt5YryP18+hakVAn3f9kP3avP2nKVpzEJYf
n1HYzP2xO26RkKQFcKLGR4MIPKp5HFwYtlHO+V16wWB3fRMIRYEDocY9DdZhq41CQR4Kdi+2cXT+
g6e1zUUrdrWeSuya4KtXTb74p4iMdiKnxVSbzmEgXEaJyQ9pA3/7h4W/EgpQqw3x7I0XEzCUUPoy
Zdn3rEzVA5tnNDzDsiZhfb5KY2WJBePrFE45oAltUC5ZvgiEf66hkrxiK0KpCvtjNFQXOuuggPUj
SDFk+lWdduKfri+7gEhfAVFcJzLeXiwcn06ep3lToPCyqtYM/NfxbKOEvDt1Ivg7sGl9yM8wYRM1
9bpx82hRCSKUiZCyouKzYbw8i/S2VD3AMcxvpEOG+k+UDcJ16+Vx9P52i0h/Bhsso2p4WxpgNryY
vyFdoRNk0b0jbefV+Cy4CcKog9SGu0hzG4HD1UIJJiO9J1Fy7KoMijVvQaLXqgsR9RleibKlbpH8
MYNwve0xydnol0w+7XygQ7YHET2gCYHHL69kLsXsaIKZVP/t1AaC//vOQ56rhKJiDtHr/ko9Bu6g
J6NWgHfHLG3vTRMijMmatCAhQdSAAtQ9ce627ZIBsY0zRnHjVD9wtbK8imkzsnHc/DEDDT7Q30gR
jmEq4BGQ4FLgnX8ohEB/9KF2GwTOQFl95R9VoBycMP0YjRGOrO8c55qJXCTt5RqdLT3RuOX9uhcq
6EXhtJ51pyjLxFrEOnghT9Sm+wUBs36aWDXEIGhUnftTp8F6X1lRzSvnDgUV8TvrGnZhRNMQKXsU
7IIoQBOOeQygVYePpIkTPYjlIlaZrEsdi4WnAy/eXzrGqCCfr8taCBJqDwehI23zQ6GKe/ckCfkg
HtaEcNUweql1cDkwOyhnCgsVCYCs8sVRfmqhqduBqHMEtDHX5tRyW+t6hKqMYT+XUSvSOPqlG192
lJviCG7nLvD4Ync96wYtvUiR8MkguDVQT9GNUudHbMiVuwdx/UHJEUzjCJOLVFXlCuNiplKttTD7
hHMDIFLOWhkN4dUmjadug4tkZwsofVKL9+k9RlchJcFtRV3Huqom9wtJMTI0er6644GJJvIqxEep
YccFYt0V1CUHH+4v0DsCll5VkjaM1u2U7Q1rfipys8wQcnBEKalQ66EHQaBxVUC6wP91/8EyZSRU
/deYqAGoV2BC0Xj9yoSexZB3U9DAp67Ug93e2tK2Gh37RsT0dz6TDNyJI/4sDd9sW4n/+CzCDYgw
IiUjDFUjl7JbdykFv/5i0Ueg+nMUsvvBBODZ542relN4g7XF5uFLbcUhwBpHnbfNbHCb+eidHFVS
CO7T8h5eptqhPppPgkXMPw0w4kmQMjveHbF6BjJ9r4eRkR+EDNg90fu0OWYu1cI8UDpZuBzexYri
7kK7XydR+B+qglWCR3+lMNwgcA8hl/py6+YEIBNgoxCb2Vq5neYDfAGsbuLDNQeWrqeBrX0INhdM
G8WeRRFAmm6UmCTLe3TWOSW3hBv01lFnxo0IINeCW9kVFmFs+uRndniSWIM98O8UBARI5Ho6Ezlh
l0NpStUZkgIARlOHAHfMyvWoXcKz4075PboDemNjivBmYJjzL1DVSl6sXwETTtPYMxbzgurIvl7A
+KzJgSjWa/qS798JJ1IZiwNpZnXDi2oCx0im3w5MWJhsNGM27d9HVn2GO0KgNeRede8c2bq963Xk
2g3xJaYmiCq4zngA0Q30QzsUt9tmc8/PRzX73bGXlYQuNT8S6drqvmU2MAa/mUK7v+cmmTkrtq6Z
RKzGkdM+gUBcIiqR7eivjyTPMPk8TnozM3ClR5jVuIQoenb4qLioDFb3cmBETDKBzO/HwzOSQ9gj
zCfVKsdigu6359m99QfXU/qiUemn+fouFBLH8S2cyGFBh1ZTWqbHtz0iSomd9TyHIvr4QXOtJNej
CJfeH9tPnaH/iI5jVKjkp7VwBlFM47fEzKCoU2aMMUJon7R1eps3cflX/C1WroKO10WyZ/PXGzbz
8YtiahN7iyP2GtmHhYPWUB6R+I26cdUdtqw/3QHc89bP4VJ/XlLqclthb514X5ao7jFoZ5VR5Poa
haptKYT8VQjKns4tWGIHrcSOnpWafHNw5U5EkbyUrLG+NuhIHxsypXzaKh1WR9j/JyNyt9CIdVIo
7a7lBVfptJwtZFp4e9OtiNoQ7eAvdADPS86eeiTPMprv4bba8V/PsNLxFj1ZfS1bWJkHOTiPGB6Z
gD8qYNmCPn/ucldBMkfT2ywT3E8pfOX19f4zXBOA18sEdK77N72QSRqVq6ybxrrHmfxaAAG0bT9t
iy3a1mZOkiVboWQ8fQUxCNe+AguY7P18GZs39KUllvc/6YhzmkrlcCvACzNAOpqpjejiexW/fHGq
KsjuG92AiIJbcItRAcNhE3VpayxHeKfvy6gdmVbLe8WtiUsQDp5V9AOjLLO2LuZntzqFVg2jSjGv
MDuY9CODIJVf7YrVZnsK4zcpTOdXeB69stBZUXXF9TKwo56KyJXf8Cyk9zptRZj4HSTSLnXOiL35
Q3+HlEx6BwzRzk50TFEYEOCFmFLvLpBTJ5IxFFvkhcQTFPbula4jTobPkYhhv1UpSvZkK5F8bWVM
ynIJmUU4oTS0J//DDYpzmEPFzp5j4vNOvJnopW9PgpM4624H5KWZg4VWGBWAxNoRyFtQpN8SDlkx
FUr7hnQBlvoFr8vs2iPcInA9ZJ1LawiV02biO4khpKpf0d9HluoN8POse1JFjkkjGkS5ENNVev2a
7hotlQHJNN82NO+JTBpXAv/CAMQkemPnCpxINpp2dqPvxmEGjWfAZyl4B+ZvM3N9h0RrKpNf6tW9
ALSsnQHvLIQzxJAOosUu9Jrv5KOST1wNRb3au2PGhljxL0mwg0OcLiCj0bo8dPQOu/gkA49iV5sL
ymzApwV8UyzNmvlXvpAoYpV0Q6XLjrTrWwhQu+JHYnpfRQrKdzxoxxD88VvOgqfZa4zqFgKXncDX
8wSv0hkPcH1gJaKl0epsFwFn2ZhDH5sr8j1Zbq8nRAy4kI4iyhs7rZCLK3IzLkyEqfA0eyiuNQmv
eL/aSN3o1D/bUGAdoQ84gH998UdIspWMrNr7ae/pYdnnzIPs9cC5j/LKXSvNgtSrL6JYMYngFyAH
AquHs0EtWLaSrfonFO+mBJiOVWcFBqHy84KCtHZa+h4sWsNtz6RVXnT/nF511yx76umdfTq/55G+
qofA9qP2HVANC/STXdLMZO6iHQMN2/cZjsqZJ6lp34lcmZ1SvViXsWiTZTZ88FI3HNtVQm2OA0R2
lepGDSAg/OGjzMu+YM2AjIdYv4tz+VqhRzS7OCh1LUPYKMejuhR7hGDY4McqE+mtsxMkvOUmOqmS
Fw7u6tMb0UJP+PdipBpe9fG82Y9iskDSjnjcrLW8nZzyEX5dJStbPP/g9GGvFhBaTIk8YDgSJ12r
qBAkZMdkMFL0i/pB4kONIOqr4KTzw7UmNkiCgIgCiv25uxOA50RIQelu9Q65wyUT+t7jN7HZfRRk
Gg/ZjSbhRXDcRBwBF2nKain8mdikLkUIEIUDvxu/TaOuU4NBYmXazRQaU39el6hkhPG4f1x//WQt
UQ37Y6U2VdHdZqPXt8Q77wBeB9fTJLDo6ekQsDO8NmRFhzc1yp153LjA1q2O8cAbWKm2gUQuM6Jz
/81Klf6SO8CWvAoAklMkccnnwdPzf6euvKClFrs5PIth74g0L/MHdhsYDLMZrLh1fcN54zXxeM7J
66JUw5EmScmje3q9XvYO2ZQb/zSMc2soTVFIHo/VxFAizzgecUaAkmymon5Q40LydUFV/p/KUpFW
oR3vmyrYCekVNGTynnMgxATqgIo3UlsZiK4H+THBTsAwCHSrwdzBNL67aUZZHnr1MpLyWJ8ey9Dd
chkvD/4VFzltBNhxiUjndOG2DHhPTdlMjsYEL+owtjXIu6VuOTFtqMFGgeM2QYauy+4tlZkaYWPK
3FyEgzouTkHdlnnWuMitC8Zyhe1Ouek1BQHcMt8OX1hXcO7rHUmvgAfW/NqTd+0Aa6mlSuQl6zjI
4eyyUAzQ+P76NGYOAaNUsSMO3t3zE6bFofokCNiJKQ38P6bgmTnuKUopVjeksbJBWBd5NnSsEpPe
F/J0UIFmzpt5ZFrJrzDaqk/qofWWH/YMcHTJbZ6uVYv8KMPyVUcUELFQrDrtZH65fWk7cdOVps1a
XCbWQl/GtKMkrD/2LFJrU9gjq0SzJiyMSxGKl2XZOoOkmG7TSIgrRvuWXCHswjMRUNTlaTVTZPts
/r6W5jXaL2gNxy+Z3cqcH1JEQmT1fce4cZuqUxeCktgYGLQspzkFfmbsEULl2vTwtCISHSLxKT2n
/XfV43ZXgxqucyNkMMRk+m1LbcMuV2nosifQks9MlwA8IHEnWrP/gUtO7feHB344GVNu7IPqoApY
qZArHOHogAXXX4B8ydjYQnLXjRP841G2x1ogDHBDXB2sTSBuXrdFGYgLqVaJc3wCNC63ew+sjwlM
BZV+/PLRUra1W0k4glk5MFKy5KfwwSY96e+pcLETTxT4XQsTryLUWsC7rCzYGL8JEY1LuQ1N1OiM
3tdMKt1i72+T6jUQYyud5BmJRQM3AhbBpq82fB/ekwRDhyeFZIzY3h9Z7YAXBzuY2b+7n6CfdNCN
mGluxWqNe47SYOzbgL21zn0ecHVdxRHruqCdwdP8JObhlqZza1cA4R6KdpdcPVY1sK0twuo5kd5H
X4kUkHAleSTZjfuywvd3xrODZOcXvK9N/k2Hkci7x6Z52vTz7Qe3Tz3NegIiM5IdiySaSgYmUFPr
fOGsbJnBO3KUl0NOOG/oXmeWEYfIw0mDCsm79mhswPon2Oiiuz7HX8rtakom7lODcPSLCEuQX/iA
vYWC16m+dqspK/OLkoIwaqT9xInpLhpdkDNcfetKaQNm7OmtMK5fkiTZy/yMUbinSzBvtNGGGD34
FQ0eKIxH7OiVZwj2pO5ArTpTbsKppsBuEvG8+StHVsALk4AFUPvfrESioN20ieHbc/FuLxKAEWK/
JtTKeGEAn7r707nMdokGB5rb34zDpkUbT/Invb7zgVeT/evIs/O9FJstwSH8Wp4YIdQOH7au918Z
AyMW5TKTQf5ZcbyQijcdQrx2e+AWoaeWadgNSRMtYlyhXXYScceverbQjzVVrVWu+fsg47K6ntEh
t2EoQVn/wKnAYeLq2qT/7RYyn6Klkz557r/Y39r2IEHmrMT89e4m+vJWXmFgjotmcsqMh2Q4gH8b
ylDAKMR7dfB/mFuTL/Zy77GsugW0gxLh+blR5nC6JaxGoY7TIOFLoOHHKTMxUNxHz9L71VDngZ3P
87sgVjanbzzTLFOSptF4b/yy3YYXVwxnmiG/VeNqW1LckW3CLuSCHjmgjFAGccBq7TySCWjo12Yn
w7Fav04WGlqOkE3LoIHnCTIBm86FT51IPtabJKNQQ+vTh9Rd9uZPfLehWvoqJYeXpLn+Go0eZnCB
TVNek8NMLVpII78NjRp+OEnW/wbMkRv4zJ4z8QiUH3aVUwLxoVOE+1lAFdSjb+GHNG70/0ByQRxT
jfPEyw5PnyoReid7siK5Im7c4gSYUaWnl7PFak/Jkuc5Qv5USISuPI/6b/tUm9sLuTA9S6x7YG5E
KVSbJNxlnw3JfYiBc4Q655eBgEzd3wwgw1V6YZOz5mmJ1HKc8JDsVh5ac/9K0/CCf/9Mp99/uNIL
pjGC6+6ppGRrfraRmMzP0H1QTitongryf92YL1F8+0ToM0lg3htWzmeIhakpuv2vwq6yPrltWEJ9
8Zrd4+mvflZMwbyjicec2VFl4IW1a/FlVG5wGz6YuqtEBtbOHDxn9xUv9KWtc5JeG0pMAHpZmI84
RWaMTUoHt3oZYEWdDfTBNjLilvqPvXaG8lvbkPWm1rN16nZKW6/FVjuTCHbPsy30d8axpSBKlTl/
bsVVMtzNAxNf0/erayZtziQ0dwU6HAKw3N9pVc7EAPWiBjVbbRmJF9wjMo3mKLh88LobHZx5PPMR
WTIuq8VkNu/dj91DkI0+PPp9dIceiG0acbqGl802QZu1PZ8yqkXlEHNT/Edj7U+uEgCXn4GD07uk
XVb+6CB8C10bxEicgLq06AEHKmmOdZ0H9Rfy+/p9qCCaXGu66H5OAi4AY6BSqBA0VpQ68+hDIM5y
CyaWCN4BaPjhW/J0txgCTld9DQaG4LLSuWlfmXl/YlgRZbSeaZ+d9ytY7pdR+Y7ZQ2K8SewUgXR+
t5cQWm6ntj4NHblAdSlojQBwvtGY1b5hHajO1iuF0oL5G9jOGWVEGjPLaZRb7Jq/zWjZvmEVYI6V
2gG0U36RluTubysD1C9LA9QxSq9O4y38a8mDFYayxyZAQaAEqZN5YmGEylIvQEpdmX4t7keZQ/1a
TIKEbnBNRyEYywasz9WP1V7qaaDO/Zv3p0VsHtvJMloD4jtsmlGaMgPHiJSm9EdxETyYIq8YleOE
RGHaUjueE1QAqwBVglI0OFjcoPnMZOx2Is1HU+VmM+dxCU+A21nxDfsUtpJCNa6koP4S/QT3NGNv
JtLW6xE8+n61iI2f2vIngdd9QE2YN7itoUjv5S2FHgWTtfjAAzgdx4Ke5pH9ixmIsMttzt8W8cUA
IodW2noXC8EnnXO5JZfV63HT/1xuMnC7CxTH/anhDgiXLmgRdPN1m8SBunszbjG9OcqVrnZkO44S
S6Sfdft3XdFn0jwa4DvfR4rvZDojO8zrRsh2HGnfxLuRaIehtkrB/9bKdf7MK3jMbMN/fymb/5Rw
WGpL7N/ow6pvfMUk36WUuwS6tdjNmS0ENbDTZ+jrDBSyqOp+41eO3JEGNzeKEUfXFksF1PrEj0Wx
xt38hGlLe+UMTtfw+gqXggBD2l5kRX8EkfaBkxrqd/lKXfFziJBK8nHWHDLTlBH2lCeGB7Ic/HOP
WaGckoDbLrrg+1X7NgMd9HkB6BE7wL3L6y3aA27GeWYWcUR3fffB377eKrKlPsiJTBkcSWh2OnUv
7BZ5ZI7ESTBecrb5BEm0D2BC+7n5bmCbZGw+nvZ/eijvdQQqNYpmS48HOeBMmcW1z36ev0F5uY9k
R0NJM0renUcD8/9Y96CFfNxA/66GW+znLwzEREGGVsZgBi+yTixQMGQV4dGBvEV/3zYRLOJnCxP2
GG3JpeTCyxdahMgDMRN2/e2J0AK5FSyf5GoF8P9nrgDpWHObEb7LfucC5Drgkza4d0kfwnPj7dsC
61HReL5QRyMcJ8eg67Xxp+RVe9weMRKEwdGuGMsmwawh/rRlZyDTV/f0+5emkQLOvWIV9Ei4bkZk
oSmMzAmp/+t/2y7ZR9H8p0tZNwkEB8Dfhnj3dXHFTKFfUK6xHyBGSFGw6NmmsmMa94rWyfq0U9oK
6myQTSir8cYXWUdv0FtKPMuPcHu6xAQKcCfTNs/SOyDGtnJA3nzPIVLMCiLGbOcFpHunbI0ZpPuo
IRFSKiIzi90wRgrhRRVZTkPZAKzgOjCqnh7p/3ZmdwQymMIM4uTuB6leABUdR4ofe0P7Ukdnlti4
0S8ZCjfKDlvcHzsrVm7XYkU2vFcvZW2c+GQWiiJqWwP3p2MYHBGhldENjuPAsXXK6gG+iAZkb/hZ
CZwLF4hPoOWvYGpW9MnsF38NKPCxxR3DMwQvXwNmXKKJwrShQ9X+3nJzEab7OlHK+OVK0ZOhVGe7
faUHBIfA/tJ9Yr0/OhfUM4zg7K/aIzhAIspF5CFu/Z6dAESMGsGNElyhc6i961bPht4zANScfSXM
JY4iykyXFmlnj54n5d2nbdBptmNOERZ5B0PEcuZ65gbKAqmIkP5495KgE4vAwvWSKAz3wRj4YFEv
X7DJI9xPDZHpqnUwRp8dTwHmrnQicEhclNtcxjsK/0Jkv12M0JvRiUPnh7wXdnAAST3kAybgRdBC
5okZG6WWT9fCKWhR6FErTYv1+G6b2IBhEFg6ix+8cC7HKY4oYlJrUummwfrs2t/pQe+ncTrr4c0U
XrUN8kJnczU/Yp6RhjYgLWsmYtcom5bq7RHP/4jJC8fYEqMPQzsuvyA6YW6woEjSoRL8N7bo76U2
fi0G3GCMhqxDFeyIp+MWysEssacaj4i6DVtt0Mzasx1980uTHvs/76CN0hZv6iSLXXCYTFo5wrUw
h9zFqHBdhOgg105lmfgMNNp/4C7zDqKxwNy5YJ8zcasm1tB/CgUcStzvn2tgJZvz3tM0PC9MdeK2
b3cM7/Zc4PJGh/yOnoWfEsAJGbmWbODXXTuv/iMSRjO9tjbglyIqVDjtW+1GJF6nyaCYGdlQRfMp
Tbs9XgjGIQYYz2t8wx7evp1/XvQqomYo3ZQ/IF+yrmE1SPXkqqWCpqVkO70L23PzENO5VDnVaPHL
YNE8sfrSP1nL8RYlPIXMCLdvpd3XsUwI9k28O8bUh95HGvSru8Lo3CVe2UPiP6a5s5iL5hHSos4B
u2qLdJlj3fvyf0jF+DVQlVuiF24aq2VxXMCzcQNEmeEnFirduVQtw9T7UMZFhws0jI3Dm21Od2Ke
tUtOOdfyyjQoQmMyFctJjOBnZCzN59fFKZSOdd34vBYjxwUpjjiZDnDsO2mnnXoROAtLuchvVSqH
7HAJurqz3x1H6Q0V+JCj6PwIW1DTZXrR7bzdWnxGVd4gdLk2J990uNdWZeaFNX9YEA8eQj4yHCej
f6YEutftnH8jVv67g+7Nr5nFUxHJL9T0bnm/bngWkqB8n816glHCo+IbDlbdDioEidNghODayquu
+5lr1gPWjPeHwHndOBarWU41o/HFrrHcFCrBnEvjXiSavHYCoYdjg5HuKKbyeYiVD78qH+WL5+LZ
ytuWV3hxKsHKwLc2yrpDphRsd2b0SFddyCF5C6+9mEvJUFa+4EFgMHsCKe30OmfB5GA9QCjLxL21
Tffb+9AjgocafUD9RYtkRbMsim8wSAZh5dJl7vZwXVChKka1/056NZFXfE4UhU0Ha1DTQW73Wr8J
NzIoZGQOSplns6nMNM/6rP0ZR4gifrYra/H//JPNBvGWk9VI9LJXBFHrkeoRx2PoxCoIMDgSz0AF
kTqVlAGLpI3SfLPgkzLF9eZrksYL1krnZHQ53beEWlyEUJBDQHhu5Vk34HYos42x4cOO7W73/obZ
kGw5zRiqHiA0i/rWlzqaQMPAe5ZiCw4GYr0zBiQ+e+my/2GOaPuh9Zbzdk7RR/7916jgWSKK8nYd
LU1Gs/SUMLbAle7xYricqm0gCsoM/S4moJ+R6VaUIworbVgZkFtcu9139H4zt+LXSnjz+y+PTbXc
CvxYg3ABjp9SpsRI5e5KsXGjpZ/HH4iruZLHRUdEJVclCiIQzGfg3/5KZ4LhJ30a0naG7WkCR/QY
wMI1I3tKOJBuaYX0IksbN535FNPc383R4RVmRiBjZO4Dsi037wRne0L+UufYxjKCNfq9EBymQb/I
inJVnlMamEGzJBCgfCPvxhxv0SDWFf7W+P7L0cLQVEoSl8Ph8ktGTq/hglMWw320KptVUpAwHyK7
zkMWBckwFvYayo806H35uTya+D5Kr7vL7ppQtGns85wH7ad1Wqc51bhoaYttsnYzsPlWDwHs0DGn
MvW1hybjaWOqgVxRpNlLIU95eHlqQ8mrz+e2S3jaFksfd73TG1JKxXnpU0fppuZpryAN1Z6qvW3x
4kBPMlBrRfx70iTpqTDK64qm0ba824BXd379pCbE33Bscl1oGmjx6J4BeyeYdxdJfh8+VanzX65R
FbDl1xI4hDl6ULKiA6EHoHBohRBdkoXSfQqX8rO7K+NBlCiloeLTXoxY8NuiggzHWxf92748OWNB
aFy2FqHGTnZTsq7ciuTvY/+GKX9X4Tm35qrZtJjRZpRIrtPa1WuzLhNV9syFPEFhSzvUkzxJa9Tf
dOhlqP2MwTRka3SncUypzkvWl0deKLyKeNamV69TZIcC2PYFf9Xd6F8akTayfXZx9jZiGJm5R5Qp
OPpdrpYBwkw7KZZDpzwNO9t3boZqXHQg5uBtFNCo6SPgZGEeQ7HWRrNn0UXuSrsFSNsvaLMuxz0v
qM213P4llSV6a7wgiJnX1bEH5p0N0uXcRW+poCBZ0kPaDM6Ko2f2o3Qdju0kT1h/GNeXJ9kTSBx9
/7RGyUY+PcnqtEIyH/Rpj28g2x9oX50n+WGoNwDTl97B1HQi1hE3KYU93LtMNKLMfnKA8IX3M+8i
ZIKLsd8wytPnn0HO/d0rK1E0iE6cKqeeZlPDaVtnFKBnIyMK2qM3Z1pDAH+W57B7F0T7jzKgItsE
Rwz9phoqKYEsu9uJtK6XqBxOat03ecyhRwuRInSt9Nc8mDXAjqLNUHpLkLPLDnxDyeXno31bicyj
ESw9yrBh3j9Fkx7u935F8kS9KFiCwpNGHdtSULYdL5Sojyx49HiZGS9Lcytzc0KESXlKa7RnSyxW
lohZPoyhvsWLf1WDK4L83WSBCrVbHrp7X4th3gYYk0kJ3xf+K54YJvSSteForHV21rcaeAHQW3kY
GJmfxtuBltNhmjEoxnMpu8IkkGUo5i+VEntxIC/kJN60+pJB9RT3KLO/E6e3wRFswt1qQhb+yjTn
sXlnzKRZQk7/uaLMIQjixTVKzL1CciCWdfrtcjT2rjRkt4pQWhJo60vCDg/6SbZ+3FyWu2a1P/5e
ScsoohxL2e2sYtsKr+iDQm8ZYAejHZK/NJpBvvY1HfXZgStwFj2zat5lcP8wb+2z7st3yniyDS1/
ZBv/ELykWV9NiU2EPa+fTV29hv0KXIYLahH4lVJxsgzhdn/KP1ATSUKFb5I/10U7oEMs3zLbkah+
PC7yvtRdLwvnfopQ7oUKgIscD9BgwZuLZ6DlK5QVsg0Ulzhjnu4ODKnpM4BEfJx0HQRJQ5HOF6qA
yXBnrjagO1pWRp+dRSIi6jJTYYugfe3A7oPTIIdhWxfL+jYX0yqAvF/H3T3WJHQXpfK/bbP/3Qhs
tLB84N1lR2x74ACgzlVwB36Ocr2jqmmF1QOnUZKQ4BtWCsDXoLnzt4rrmDBvrL0tc3vV71zxvsA7
m4/0Yk43kegy4nLUZUVN+AMcJAzWSnSsanxWnYZbGL0Ztz3miExi5aN2Pfd5xg5q5FpE7KRGs/3r
+BAtcds7wahMmsVdotrWm70z99a376ClUwa1GDyViIAeeMEex18E8g3DX43YKj2IgA9f4X5l7Huq
xWIhFZjtcT19JyEs7x4R76D3T1z2aIwwWY47vT9NU145vY6WKMH5SueDJ3EIESuqEjA4XjwRLMHi
bzufhJbgHbnlkFMpxlq44uBmLryfMQLoYbxgSTbcTR1jUyP/Tj6ZGb7lWrETrgc+cUZ3aFAqCvqM
Y7jXjBpzGPkUPNVmAm4CC7NusvrjnwjgwyOOd1f0muj92UbIcyEZYf+AhRarOn3vrTQU1mTVCg9f
MgE72459uS1aZ0uV+eSwMQU3THZ4KRMsBGDDkhxfAblDG3w9iNPwRD8GV5ROenBLVDPJmjWmE/i8
1PxcnqR3pMI4RZs3ppwAQ7eejH27sxMnfetwzYjorLircv2/O80t6mQ/lh02RWQSK0r5NV9Xub5L
aPsVomCJMhtTzC5iDUxo07UcQCS9srkNHPg4zHPS8y3HzTrZiDlOt1JSAN4kOz+vVg4mUvLuJb5O
twUfPMK5diZKm6CivXNZQCZtMO6wSIx7aPfraemzqE0dABvmmfvZ/8ssZokygO5Kk6gHH5VMkU69
RCDSXkco3b3YMRQ4bK292acFHhtey3V/EEJE3gcHVVy7FnhzBeyyg0pnyvEo42pckAkWF1b6/5mE
E9riv68vlv2ctcEnRGBDsxB9z4ORHq9hAE2Mv6vUn7QSvqdCkZZslIUkfIR3wXCJH2QLxGjCkg4f
eEvdzmVXe+X6yXHtrhI+O+ettICMyaajJAswy8fCP+zOblflr5DS0SF4zVUfO/F6t/xXdR/oM6jU
W3BwIeqPpeK4ML0nSN8yWuqjmn7PNmchSz891EVtqkE+Qaat3f4z4vf6bn4ouFMBYuQkmZI6CuFz
tIGB7JBoDsuAJDpE1mkJ+FuDsT+xoIuwaXvExG654SPfLVii6U3+frT+rKzPv/y5B1RQ1tXF7rRq
LXnr3lNSdkHFPq1kGkMFXs0qTsyh2z8ElrgwbcXkwQ4BISDZ9qT+x68m5xQ9ObKO3TXTDwGZH2S+
ilPkQG5iivQpHp+sbne+BUv3uSqQr1/cdxe1g+YmGOcoCHrOItkBEZO6YLBxd0ZfX1lNzSk8++nJ
svuhQ6wvfKx/Z2p4EwxkH9Lvbamf4GVDxQxWUibe/rZtQ+7P5fxlFVYpMubDTnlD76SWPHLA+nce
2KtUdsRaoZKtnWDP0Ro6OEZDrgOtJeoPZQdNO0prGh2Q7fKzfqB3niIKH2IEX3m994SkRmVfSY/M
N4GBLPjftghqz4lslE/6ckQaECqVXaJFZG5Jb3gR45p2nEDP4Y0bdXNrG7ftWzcXpsBt+NTR5BzN
u+caxfp5phA6PkK4G7cOY4xv3xl/mAWZnTWFmAfMUegtbKp+qzeoUPk1YOFSLrOqpRGuqVfLwfka
mTR2uh/1eyH/EEVFZ2AHYIgMEOkFMmEeSe7fFoIYlrN9uFUNXnFNm1chsDmOnV0i/ZAyUz8VuPvl
AC3uIkY3YvI1ZetSmfy4HbIlKF0Vn3H4Ynp7740rmpVVlxzgs53iEkd5Ie8Q1RUbzgFGPJUUNlTV
28x5xCgKCb3nvwzx5QHLCJYjW0RQA9NXc70+67CWFo87vjZrJgG8COHAM28JdDXvMokq/ZzZHOB+
vh17v3Q1vu7QiaVn0uSLqtBvWTPdQT85HXnl+3rgDuA1VuqB5Xdio6BBj5RQqvqUPgSNoLuLPLHY
EG9uXHHOctyDRIsqUwp4czT/h7bPUq7bpvQA/U07DjLImJrVfaN6j5J3jDYNAPTe3+XENjCXD7U4
YzwJozrIfD2CkLV5lTEKPgp72wRwq5cRq8/PVHtvCO1XrWczPLFBJ2xwrZi8Ua5dIlz/fsrZLb04
FWSsVL5z1KS/GIbyfmp8HFydWiRCABc5In7MguBs7EfreS7Qw4Y6rduQ/Q7muug2OyoR3ijaffIN
IAuYxLmPK44xUl9ftqjQzmu3vMQysV0tLZ9aJ3dIh+DME2PKxKDjs7UIuyIs6bMuyQnzP3G4HXtT
U1kVVyK+tZOyWpmox2OVP8+aP2Y0tvfytCZHlyAS/qpi/7WRzqZKFihMPfkC0L/XljuLvvHbUT7Y
rxBhjL67Bl39ml1iURoJs1KW1NZlzwbckgkcsYTjJkxW3Y/lLkehaAv2tgAASyM8Z/kKnqBRD/Xm
TAV9ooGYAZO8ustQjshQkay+gxSWQEwib7jlUuH7UPCx4tLImfUgpudZvPl9CWC7TWUdzej+iftb
IjPLVsUGe7b6DKBUEmzxwOOm9SyhdaqVY7NjN+vxVIChf1JzW0nBsZHTyZ80yABmv1iB3dyuOByR
3n1FpJvGWimF3rBhrdNkavz2QSvm4OPx+DdpMa3W2fA+qFeSAyvdWdK/fZuuSYatip9YsSOwMYes
CvTydqr39x49pPxguGOfpjJWm1LQPTZ0QLr95XbylbnkQD6rTUcMxqSqCOF5718e8NoAYJjVPs0o
3pVDDm8WDVgbmmtAL7paB+jil1aeR0BhnMma4sQC0Rpx8pgcyc+hqS5BHPCRxXlAPuvqOY3MUyMV
m98MasKqiqWgkl7D/nsT2q+p6oo0vt7m/ywbL94Df+FQxazFJGt1gagnhnIevdA3xrwd5MvTIheT
QiX37m4TcX7H0yTsX8rhyRXWm/IAJcte20gHjujlq8iMMIGSwLtyhkJRKzePWOlmik6hlVUI23p7
m+xAI+O8oPbbFs90idaqHxUihEj5Xjz+LR/TRh5UxhLZ4SA9HJVERsLa+BT546npiUtlHcBFQm58
uaMWygAuqk6ssBKwMBtYirgOFO4uIGibLXw0WBkBkzNjS9ujyERD9oxnhsEy+vv4+g1L08Xs520q
9lh1NABFQQAzPkkv9pb1My3jA4TWH8A3SIq+3ZOWdNC48m1y1os2tUxeSHJhok9P+fTX15TWUitM
xNHqhDRUoRafmpQcKF9Y0QlHPpcxjcrLRmzEl40TBekrKOlftCha2vQXS+2M0SqPIEHPKCTDb52J
HQGSYlzk9TtXmAHkabtBGfhXpgB6D8Mb+g9CMtkO42IOwpC85IcvSFl29uyNQeWo8FmcTR9DxQs7
hQpKIpHJ/aSszI8hz/D7PLQ83LoXwuMs5ehMGpHQxJSA3/bX4n8UF8/MlIqg8pHUbm9pWLUPWeyj
G0dGU/nsYGPNS31w+LZg/FsCWZA36dUnUErniwz6AFnp3UGcXTddWCfveVgezG1eUOGvxbnbRSCM
2VEpMS+Sume9vl9PIv64z18zC9SBJEntLBgxD/Q86Cb6Fv0R7yyuq5fv0zFS78K9Kk/svig/65WJ
gMYnl91t44wX6RemXTF6f23dDZMXF/JWOWObGp2SI9rishh7UCOvRCQtdJVBaKx740j8Nr+JJVfM
2DDPpq9M70paZh658pn6MsdFRz238mRX9O7svFFSIUKmEA2qpyJZb60MxuI2H2sbfucQ62wKtX71
0jnzweGqYIBDVSwW3ArJWOSYPAZkhQMex61YNeAoJHVe45FwHfesU0tDsZcOvBWkUWS/NmobGfgf
LmmFW85YNNmxNwDO9eujI6xTmTxiPNzB8IDEeHi5b99fxt1TnkezpyaTUqgJQ3vJq4yy8fftIONe
GZcnG0Mugy7dlVZ9K8Xuq7FXMf5kOLN9HgNgruyIXKKO6qKWtLusSJ+AQQcn9u3B/9xFMwpUSUVf
hpH9brgTmh/dusFVcCdMNOhJV5mfEvoAo90WDdVdzYXegI7E5CNhTEse/G9YgMv+iOgMLGFoc+iN
0PlWPz03yHcAdroUWXry6NfX3PXx3op0yNK3QTkj+cdX0XBbPSbhE8MHBBVKhDCuV3xLwJYH2Ybq
S7BDh46I3FLKJvaA9KKoEEjaHEDVnO+tsFE8oOtasnsIykT2uw+ikmjqHFJFi//pfuhxLIil9MLQ
k5Ks+0EMhV+6LZy+6uS+UGfdXI5k4iP/YJ2Pp6OWPLjH2ws3VNTA4sO56US+nqIqMRWMC6I7yYzL
QqonCGZvUEtC/0hIELs5eV90GGdlCycR8L2DsuPj8myhQH7JlZtlAHexCtsQ5I3uaht7zzSbJuGy
GjHW3qdixmiAHW0HnCm+A58EF8lqzjevwonP+jJbtUxhyjZZUGwLpg05IqyrOuloWoas3QXCG28l
4p2xAwKoQ2sbSk5CF/w8LZH0Ul3gkjbbtf0CluH0KLNFVyr8eGMZVb/bq9/+mei4EkpOCK7xXzBD
QcTcCnEeSY8PhpbXRVpQIXnqaTH/akcLNAl4exvulpz+WUq9rH4Ss9kJ5cDpSKH5VFx4UjJ35lQp
ljc+NL1QvvIwz7DRVjRBrHRBOlNWq40zftHrkvBrZZMwaFdo85SIjgcqDZ7BfVQPTXUg/Ah+8om8
bqFkxA3BLRojb961//y6Kx2KqhXei1Ejd6vGAYUyxmPj5oaafXc12K76fPjSrU0vZA9x5kC33/XK
S6rzn8+B5+Nq5h5gH6Dz94FWGsiykiFaRYjFJWNjpT4OcEdcgbNGQtNX1v4opu8fNfrzuCEklqm7
EYFKLwtNIi4EwNxabaE7WQ2Djnqx5L2Y0kk4K0cmBMKUGXY7wIqcyvn5TJ/ACj5Rmd1IjWtPvqUs
CjO45WRz0E9LI9rim16AsYPui2nJbJnkvsIl4kEzu1SJAL/MJ8z+cB83HnKXNovInMc6+WJ1+sIa
xVw7IQkwJsl7d6qOZPQDR8Sxl9xVA6BIvsk8OlzB/N3L8soOMMFyfF6HiEyU4hqpX+ftj7GvTqhu
9L3P0X+WIyhW3hBFTteJGct1kQF3DSHwdcer3zlmMPvCm7PHXN7iKnHS+y+tGDgjHWvIi0n5ky3x
/7cRDQRJqQYJ1aXrxPwm+unNui3xCn/xudEpwTrPhWk3DOiJnmaZwHVIFe6SZ4tUfv+fuTotr3vm
GGiW7ZpVgzGB9e8Vx5jeik5/6r04MC/DvZ9LPSfl4XXZob6vbtuwuhe8q6hyNBjcvPXO7kpZ3LhO
RcT3UCOR1ZFcujP2nU2h6rct8qxX2WawBfYfUFgr3MmI6/69y0oI5RmDXuEJJjLECxV+FmrYd7Cf
VoW0IftHbJvxkuUsoX9a0CprYxianLxOt4kQAfpJKvbGLmH9OcCa/5BS4JwNkM8hb2VkduWLZkYS
IzXHEDBybGPqCS03f3pUwD8QQfkkfTXY2SUFDQIag8FaOX1ptvaV2wv5IRFBtS/u4Meu1NNkrsg1
828NWK3Ipv0LBapPHON/nAVUhIym3Q+k+uVd2kpwwYuMuRsSAsF144HxABBXR+/DmqRfRxUw04jn
MxR5uyNy0u/1oKY80akOWjoRxUp2n/lnmLpfAFM8uJoGElH91YXY3HkSSTJZGF8zmlln6prkmYSG
iD+TXddIyrzjDv1Tx+HF2wmFoVvA5I2kIFTb2MDV5nFDAL7hp7mosFEKW3R+9XPdotrszuTSNheJ
ezWcCzn7XjBaXbinrn/kA1q7IjPygr7s1WNV8DkeXKxJIkiccN0eYWudrDVpEMHCPFLVqmoyDb8d
IXTVq7ogW+o4RITpjqtLAIRDggCO6EI0+Ob1rm+zz4+F7NXwEC1nooCtTIhsoYl+KLxyVPhhYbi2
rIL/FlLsnEaiZJovPK8hTQQQhqsjSuJm1iKO+QjiPxF/dYmLVkQSBcj4PeA0dYWnpNyrqLURZMmf
UgxUqJrI2M1BkdDVVY/aMlE50y5qT7elrjB5dNn93x1yFB0PGno5W2S4KeVr64uVSDGrinhtS8t4
mXAgucVUKYsf+B05TMcWYCCVCtJClqWnXBPIFZmwdtFXFHqWuuFKKVNo6x/N3QeSL1CGGxc/WOng
PGHhAvrv75QIrU1d/4pWayeIM42Rnk2ZneHGaPM4djfGYN3OmPssdkFBY0rW+QXTz+ZvjQWcaGX2
+U1SU5cmSckoW+5KEzDWVCpWOqBLfL1AY7HZknwOTRbxhshi07nG8QmVboxkJuWnBbwGggxvcfk2
YEw6wbcd8MLQ30k9qkrTkdrZXoeKQxCChpwuP5/p8qUlaht+bIseCLSFfhombmNCS01VPvB15e10
5nTod/jAoJch5dRJ09HHP4U3AyKTlbZ06qh4MichKCwWIUWQFQ9l7gqnROR2KLTJtnE158xYghNv
dVVrMbkBZPql0ZLBZPJ7hLKOHOdE7xdIlezWE0+OmvFCl/9+uBiB8i30xx4/B6JE9SaGwpdc+ASc
1MuWpWvskVAKN5IL1sRTHP8v/rV0y2RytYbpCRLcufwd1USYhPuB/uSdt9QRzyl8V/pnBQOXUzSq
fyRy5NL/n39LcpdDWWELgaC9tCtgp5pDgA1aczlnpSrwmcHdxuZkv8F8HRcN4CbFggq6QXC42xhi
YcZWCO2Upaz0MkyT8jDci7oEioOOZkcub0HONT0BJiU5J7efL35eDB4CNZR3jAcQw2d27F/eEmfD
PW2y3KwXx2lUY00BtagMk6YZxKJnxSiVlbbzdgW8jRuJnbHotrDehBwrzM8okyBUe72cBnY8EF46
pjeHRNWzuAicH5H0ZvtuiAOl1TbtYWqXFwrTmPF0+OjSdHTKQwkczOnk8WSUF17zAS6PLSDp3pqP
FzuzF1HcP42VYBsKZBs7tM3u5k0hak0/23eKdqY62HggJmPDcv9JAq4IfSn0r6sXAdWkAD7vMQ6X
QisFsdsQeO+9QkFuq9g+0HU5Xx1EcRXSaAICVVQZ71Sj59wdW2vb6/F7ULeNaSAlN4bL/i+nOhMD
zHoAFD231tlt/ajY33gS0FQ2yOeKTx7b4vtjB3a+AQsPxMLBScVyEdeGSRNoRf8scg7W0pvFo8bO
CnJgvfzEwFYUhKUREoU9Egy/49F9Z5nsjn/FXUCPued4VH2Qtn1m70q8G+IZ/KAGmuWV3g7TvGzs
WIpW49oyLt1zX4vB9Q1yWLwvKOZtn2AJR2JotUJaEAkHwErGi/IYvvqF/678WIj1/hnqJ+rCdybA
bujqFLAm/VBhvXqUaoVuTokwHJa0LxdrjctgfSQ5GOGqVZ6LkCVdQ4gvai6cZDAQyixn9x3f3X0C
aNMWHv24DG8Oz1oLJB3G1dHMvNdX8kFQpO8mGoQpiUrXi40a12vdUIltRnueAMaYo3kvbLa+9QhX
0EHB/v7B+2yUdVOp8InLTMLr8SuKNtbFVYxN9tPCB3Yf+Ob1Ofb16VGtW7b9UeYDRJR9UdE01yHH
WReRS+C9E9lEAox9Mpg0ifsWBt9jssjfWBzgmzZHvYBmPKfI78NMg/wbdH0r7Ftvu6CPi8GrUso5
zD3suHz5JvCpSTx6nh8fcBWG9lPri0bfyhjKM9X/85FJWY8Ccwyg2Q0TRR/jCkn5cerGWi5kOSiX
0w/SJEvxvWDDrOWtYaz4PcIlBBz8pWXVTXGXvOA+C4KAZmdDTSwO3N0G/FSABMQhFyJDfsgY5OSP
b6KbWCu8hz7jel6SNyrM/ZCGX3VnNG/OnnlzBXhdPoo3QuXxpEe9lc9IfvM22IRIzXqW4Crtg5v7
+nV8XodRnGJ3aP7nXpOKcwu/pTOD2UiNjNwHkjJ7F0o4nXX5TBcYkmwtDhQ8FmHU7dTR7IfL70/v
5F7FlEifUKj1g5q7+Y7+vGy8Zisn4fP6Gws18uWwcILcDDev+6R53AsL6Wc+i3mvX/IaTRx6Ji2L
I+oWpi2EwAKpc8iQFXB6bODImLtQ5eX1QMRpTiGKyt6Y6QmPycwO3J8dQZd77gjvu1omfoesRxmm
s2+UUaBbsnNMzhm9EACnqIp7mng7PTh+yajEsu2VbwyiVIaI4wzV7lmwkLSR5Bu5pcT8J+VJbYdz
B4oW2SrPR6wSiraDUgPYVxANu/VLg1ICfR8YvviVQ6w33CNbcOKdovV+R2MADvTy8tUC9VcMGrLM
eZln5sBsLakq+SdbVsJ29gpP1blbFonCmUkPh9RfcudPQ/HC+nJCSkuBm3MV3rV3LtzD4RgDiUuA
1dP80svwOOmL07oz3sByMflJO8uYqGKVPqbj2mOv+qqcaQn1Chzkiou4uuTfsxeB0ME6SdgHh26i
nJVTsxHVHYRFRaXCn23l74+ciUdWNO0i/vNMfoJnS9e58QEjPYKpmIqmswwYlKRu4yqADampIRfT
xqlcYPYxopQZHrV8Ji8mi9A+jiHRFIF6g9iPiA2iQLo9gXlKus1WpDgDUtpiENHU1P8VifISzUw+
SyovW+i3ztHKz9YLcroKYJST+rE+b0Zp13EVCEhDe4+4U5u+jUKbCh9DXq0KlinMdWDkCDT+nxBP
Wbm59iS+fuu05MTUKf2cPVQcoHNwRj38umtlbRq9wAjQEjd1Bnc1gIBCvKZdDVLCStboI+wPCC7g
bfQw7BzuMLQACZvJgRIKkGtmMUZVOh54m14xRSXEbbbOLIg0S7KdFH2Wx+JrbVZ/klMCnsuKaqMq
txhitarKJ2FEy/USRAqNj50b8SuhOKTXcTQVXYiIkcnYxSvnimqio5ge3wT2P5iMQthai1yD74LH
X6Ht1XzPXG0L7wxmoy/NRIpwqG+W1D7VWPamdHXwd7Zt01oBafZlUNIaLemyY8NXUYS8IMgEbUUI
TllFcj0z43XhpQH/O2WMSBMTr/AzEJ6No+LnyToti68ufcwOp+s7on2sW7mbFq5wxhnuVb5vHRek
YM/7CTaBHE3PKuKDc2HsAjaqEEhRJ3tboot6aLHJI9PKK77PS0hizhYYgOwA/u1L5bbzIrtSXAuQ
S6l+iRGtmp5rCiwpWKwQY9k9nR0Mi9CWxdJnZqwInrGZX2LdIzAbupQlgJN26v4fIOD/DKBKzNsn
eL8qD4/la7yqyBK95A0FVe6WtA7y9y4mpfkh0FoGWR2aW7i2C/jKRGyASgRmkXmds2oMJICn09br
fyX8m8+EajF88yFmHHSk/KtzbV75Ea147+K6rniBTBsrz+1TJmzdLEnWvfkNHUl+U2Nf8HLvvpHv
HpnINOJb9vpPg1wRq6ErpHy+TTM2NlnM2mIPDRfcTxMsIbkKrfkhAZCBV/JnBPbsbT3YuEWtFlDI
f4VPTfD1FBC4xqIchiyu0oUqsvvLBPtLX4rMz8EPKW1j8OUnT71E+Ehbcg0kbwTbsF4Hwmo7j8r3
b/df0LuzovyBJbo3Sq7nY3jaUtYkbD/nEpXkB0aOOXYSv5qg0MCCNUyy967FSq+GphzFf/WbxQjg
bnEumPygmPjargE3wW7goYb42IkO3A4J0rK2biSUhurjAYh/ihjyT/aP5EXyFPL4DDXfoWnfexla
leskKWYBHPmm/41z4fZ1eCL/GqJAbRerGLwAnuVlnlGsKkQRoXP+a3aUEv3iYr9q7PtDtxpdHTFb
RG4tfH7mL1+K9XSeMnjnd05BdQKiYvWdLCUp5YA1R3/Snrd+e0P7dvo3sk6gNhctaxRgIbEZWUq+
ek3liuV+fYKXUpGqTnkYMLyFkWgbc07AkKjwoOC5E5a46O9Q9DGVykpase6JJi4guFK7+anGj9lH
/VODQdZBCyn5mid+MdDoEdpn7XCezHsItNcqyV1MCpwBn36xdzroUqe1RUJxiDDif7qijkKdGBUr
FIZEtRNL12ZpJHGkdwXwH3S9ZVgVM2wWcGlZWoshC7iQPddYQJppuEqjbzrBWbh2X7PSatVcrS6G
bsCDKm/ApP/n30XEMt8Tn9rph+u6ufLYmNMoOkRQ5jsTARph7z7+uqeGcpTbPqtPxMCX9XgMJ+hr
s+RRtt8MeK2zm9ob9546Z9PAgyz03PiM4OmirEkQTTXk0F4Itl5tedmGDThTUmGtueMFafjD2db9
jMGI2Njk5456zs84TUKlTr1+yERnNCOjfFMykaPEjpG3p5nZcyXzqMmvAgkDx7cxeRw3fS7YjfIM
9W21NziGOlaOWSN1NQl+VhsE5fiKalGDzeIoH4DIPkKoDwuRv81pl4Y59ja4UlU64+5qYoJuRfc8
APjZKw9SW0h9RvK4IFjMqpHG5Y/upsZOlRkApWeDv2lu0Vatr6lpHoZvvQiO3yDjVhUIzN40kHEA
mNJEqvcbl5blsRtEANEOwg1TMvSQqEO8m/jondwgQ/N8+B1HPLT9brmjL6ZhdL7NhM0FpVqrHTme
gyXGPfHzMj+j6m5GuEKj5jo/LgsShc3AOugrCZNv1oODh2rNnnF25DUHhJUK+Ijuwth21h890vcB
6L4oVbDCdAG3Z1/MePAcVGc/Pw5ZytNQkpIOdJewCio5pv3I+3tTeaWUHzKHC8yHf85l8t5iDnJD
yXtEx8M+AqgkhKCf1MjQg6wrbdSn9eNsf7B7UvPjPU6mvVoHYHL/2BNjK53Lvr1AucOFvFvcTK/P
u0sbvj6y6rq+u6VycGz99ZA0vFZEpYbFOaRKCXE264GLRDBqKEi/pIZ0CRfLAl9AYeo03Cx/L60q
qGMdh2TnuHr4DVcdwJSX6pvSmJs6Q60RTyeHeQoU0KkrTGynnVOyxDLV/1YadxExmGLdt0wt7QMH
PAQxO1LdM4utC1gTm5fM+hYq3CCiWw4Gs1ts66Qd13mKasYLMDJvxLUr9DKdE+lx4xA8hscCMC0b
FnuUMgHab2RSAPOPpJQ7+TDhjzcKNZwIPfibrKsEg1MEQ1AyxYGV0JlAf9J221npjg9OmwvM6xV9
dLHXToLbf0vPLjMRhzEKfk4RZcT3TR22VXVWPCsRv4rDRsKlEzY9GVI6f34Jl88VKsBqry6nCyew
vuOWKCqi4ieqs4Jh8PgQn6H65Z6MDsy4pAjIV7LgeDA/Fi5n54iCAN8EyYDkTlIr6srQnX43rzIr
pHRlb/TiIGWLTeWmIg+e5ESzYP37Q5vZ1s/Yqbz50h/m2olQw9WuDhQ80jYIZZWy2a6FKRdGC/5X
HydqmD0BdLAmzlyD4EY7GOB27nyU0xiM12tbvQCiT82u0gLgpZr5CfREnTw6zEK4LRGzRVJ9NwO7
TiFvB0dzIAF02RTWz7LrxhxemcxrDabcgA6SxiKtO+u3f6rjgWmuuFe3p3OoISCTYoOWATffpo7M
akfcOtgolAhFC5emz/FtUyzkCTaNt0iFjS/bmc9Kv9WMNVIyWy63OE08asWeBUJ/43iyWtqDpuFn
/4a5k7SEYd+Ua4ytQURXe2c2pxCADK58rzTgqRKHArSEKfPaXP9wjx7srh1rBIED13vziojRHtn3
Dfip/z3ZUE4PiFEDGO9Qed8+gLl5eVDSqTUG1KHiyip8za8CEayiCuY/CqYEo4D7VOUsNFeIFkMY
tHnIFKAXh4dqjIeAYERj7FqnoDOWGRtQa4aeN2Xw1m7OCmLJvnJxV4Ry0osbtL7931HDQE+DJG+I
fRimZEh3eMmD9w6llwfcQ0ii6MOvCGZGh9h7lwOcGNnxRsqrH9YZTeXMEEVyjUcIyyiDAnYKpcnE
L785ZW/+hLKIY3TJ9dT/sPiPOVu4KHX0GNbrk1vZ8w7Kn+8AB1a2fMld9O2d4U84IXXc+ds76Xmi
JDmqYCf2aTef+sj2JtLdxGBAbZDaddIurHHDUFYRk3Yf7N7WmS/A9frRV3vPSgnqAxqpfEJhoSAF
FyRut7yI3pgPahi+j+Ax7S//WupQyE3/VKpi17ABk6QabPHOvbZ7lW0IKhmnIhFpWXcjDcPKhWN9
JTROAUtlJdcn90SxdL4wLQ6yXomZXLIH1R8OMjnqSd+GkbAL9afDSPj7DnfCAnHOlIxPwKIKUwV+
B/LyyG3OgwfHHCy9w2+aZbMgz4YDAEdaFMkLX+WFqLxKSCuUN4vWarLX2oTxnsvEzubIO/gkDqTL
XdeZmUw+lQYSSoZYXejaS41f49rwR5IPnaYM7q0+tfVVUXVMn3C18YbUQID1kqw8+tUczxOr4HQR
POx/rAyI4MEOHOwEI8zD04XGdWikLiguqtc2eaRSmScxHEQr2Rzm8XPwUjfmsbqme51cute0N0a6
AnYKzkV9AG7el+/6czpmkR02yv04fxWTC2WOZFoWfG/jtovn3VxW12FxWGIvNNFhStACZZh7SnAn
vps5mj6hpRS4EdLa4dc7KFwKmwn3Ht8sRIGT+oVFl5Bpo2pmFQ1MP8wOWMLgMOsKaHPbMdikHZCM
4kQID95H6lIzSIzhwenftXNZC2Hg/oP8o9p2c+7B8QU4HjvJ1I+1BjOeOZQVC6edU3B6Ox8sdHvU
oj+8/qoKj9DkLLVF+pvSVyhPmDPIWFj+NBAQt5ENdtE9pjTek254FAag5y9p5quSrSN0j1uyglyE
heXlXQMAZ/X92M7ffta7+u5o+yUZoSEA1J3jdGKNSTzGNJAMOn2JtxiWTBetjbkizX/2rZzCxxM3
QclqGMcojtXO5q+TzGeWrx8G9LX628VgOyu0ogLgwyvyg4qwZg0Cw0W8UB6MB6hxWXmH+KDCpSoP
83lSl+26UOPJTwPvgystYKYgBhUp7Kx1niXjO6B0dCbvYKTiZwM62dRzJujaMzRCV5qwru+eXU2X
+9yQmHGmuYqNyi7XjiSKyj56NKaZmB/TF286aovOZQNE2HXNRt5CnvdypN3fa3ql/n+uX24oFwR8
V9rrncyOXnW3H8AKAzhYwbXSWlUWkQMTk/HC7YaacDr+uAWacez+fXSmusoUfU3Z3UwRkuDpi7zS
qkVXBtN0Hb+QIMAQ8xg9e6+qTC1dRmQ5WziaA9ueknbhQlwpQnuydqlfgZSkzmtQnM+fvWHiIq9C
/Q+xZpouPiQJ937zVDv0Fuk0ghq2nXpZOQaZSj2T0mhCkm3Yz8hLFPbY3QwqCcLwFjA2mS5dZ+pI
FN7+hkMfiaog+GAVpKbpetoevuFKSWRYbOFLUHi9wX9iwWvYXiHUb3Q4aOqjdFhF7wC//H4BdWh3
MSFE0GQDYFVa9/Y4YMmvZRkd/rheWF8RcvmxrWNVLvqm+NMv6Kx8fQun2VUlgIaMJwOK6aj8PHxQ
cSzaLnd8vFIsQyrCNNdyEYP65yXJScKe9Z/X0CxZ7Cxm8opUNhNuvLxlbGuh92QRkwxZQIA5eaeT
9Kx29XwDy2zBW4N7w6y3QAZcVoj9hUwSxQBde6FMQS3pOeJiaEqZF9404SoS+vDe/y87UDgJ9EIw
1vy1NacPzDCOjxhwc2FWPOpTPYMUvJQEboJeQXn+NpRBlRY7jZWKzLpyWwZA/Sl14HPm1FuqscTo
KJFqk9oZydDiVuLewWMKjAtC+e+3kigfphOWJyZAJoJCTfNP9S4E9OsNLSxLA6EjWQBrxDTg82hD
V/ZC61ZE+TgQkjvyQTkq/snUOUYF3omg+1n/kc3+ba/Kt7tpd9XJWsM8KQRKlP1AXTV2IWpfvsBu
uLydFLyX+kO50Ewq9SK8NUlhGiQZD9pHGr7uGQpbwjvwM7cT2mOO+3OMtuvPbeCm6GGI7B8ZNSao
Bz6oQUZz0mzC42aa6FQCIwuQo6tJ3z44bENLl3b8UwJ3w7fUUTmOLv79t7zMi6PHjf4TmkVfvmVK
oR9y/ByX9KAZ1LXSE4rRGC4QRhck/aKzb41Z+AdouUJkM+bD2dMQXXS7oDTcG+R4GDSGsBNzUA7V
FpSUh6bOlielbeAbQ+Cn53nC3/oOpO+v3Zvk7GHZVXc40b6gvz4xv+SCTnrGs/yFs7/h2HG7mz8q
bLgiTlyz1DzNs/PFj2mUxF8QzXol2qPqXMNVzdao8RQUnsrwHIeuXEjNzWi2aKzu59vNhQovt/fI
Mu2z967H7DaSXjda0ytc4lk47dg13IyBhnFtEESFzunAqcOpHG1f46SJVEMyQmPV9W8cXL3nLol/
12tsm2+5sp9zXcwMaOTo+KO5t8Wzpl7/BO4gRkxIGAllj3LMVQgjJur7Kv/cfWwswSuW7qQKy3QU
fj4r6uRJOHiG1RoHTqpaMt4zxgXcvxpuTY4hfGZnvEnub9PKvByPKcJUEh/H0kNa5dOqKbarQncE
5Pne8GfBQbw5xu2cGEUvGj2oCUFEFAY9y83aH4Lj2GyG1ttnOW4urLRWx5zYjoYkBjxZ+xA2JOEN
pV+SJDXZVg06MkJEDmE3F7GQx0sqa3DQIEz3hYSTgfr/nUiWpwfcTeLp9Y+I01s7k3xLgWsZRc1J
CzEcZ9M+19Cr6wN5exWilINt/yjq0UwlnMatVf8NvG3a7xxhHzczhAg2PY8ynK4VGRmK8u6GekLN
fLqFbARv7SboAaeDCVxBykiMKROb3fvatPVppQwHBYk9LBHIRGMwRtRtuiKyvDrOecGpgPyHjxYx
z5Fd5qe3jhx/CROOvCPzzrW/f70UX/x4mvJvdS9rJ5hfRDvKsIvl+l/cS+tqSfq4mGUF/wjv5f1B
tiq2sp/c5dacS/z57u70WRIe2liTaolEJXseuPczEOtOBE+NEwPM04ujLHBp9+V5yZlU2H/7voTA
lCIB/ckO0MRWRBmbCUlRLMj6BOSgb7v1YE7zqgktNysAttdiCbxGktTXtd7nLiANAvIO0X326Xc/
HNaushnzhv3tphkXJHI1gWLhZtcPzUEgDCB+0mfA0FmU53E9v/aypDNPTNzxB6T+JNvVSUKSl9hC
Xxh4fA260cGxyrLfsmoKEFLTO6cHp2dgFeTxnwjJQfU94VWy+m1t/0pAFnuGwQTCNvr6GfnkNMwL
i/S7/ec+1Q6LdWfYbUImHiQonXvxPEOiEJ7XypCpsNXp6OIFKwYr+oinmpz3EkoGkqvMVutNDtSU
b+YxkYtlwnULeRBYjh0fUCG7RXqgzE6vLjlDiKGrMuck/FRtmbZUJDyOJEcDuGHGH7nMN74jrOup
fhXzDKQLiqh7KshFRRlYWJlYJjkvh2yaoSE7Oq2cINQ4Cdf5qeLd0qcYvifbSu6U0wMCgEqKVcYL
5SlPgz4kbo774aiNfytOuKrxXFumr6+vgU2G+TptnYRmkS5dPSjkumMPQMT/YKnDZJejfKhpQQrj
jejmEF3InLr/guw2VFitWIaddpc1yvwrs5Q4QU1H5i8I0A7K+l+/F3tGoX2TnQidg9mfpOqhX0cb
cj3t3O/g4m7ZsYRBZs7Gi9DGUKiTgVuyhRoa8HaRV3OBFBGYEEWTPpzIpqcnGR+k50vpzNi49tAj
34rTw3/OjKQJC1xAPZeqoHyMEVH6k90QP6VzMpmmOr1bl0jRdYUDU00O45pu5cqnIe3lob1MMx1J
k4KAr4Ig9IFLuIs5wGn7FsmCk7vesgJP9/AZ7EQjYne8Db3GZCI/usDwZ0KsrB4aPzRB6ey0uUGz
Ee+fJpgwCUYyVg3CQJlU0MEvRNjBBOSS8x4gM3V+F2+OUCgSxon/7YfBPSSNndkKzvyBMRK6mYtF
9wkAh9ck+ugFSoFSwXO2y+xsGuXjP3G3KtSphP7u072d/TlLLS7xzHz33fqRvKYhsFCbG8uGkrgd
A+sRaHzAZ/m5DORktFt22hYyuytD5HyngkqpZ3F0/YESNnTwDnnHo05r17D75IgrTVB+2K+BBGHH
TfljQg/yHreV7lO58JVpsIUWEKSfQWn8Dsvh0xsYAjem8Jrns8+KNKYLcdjsHZ/gLfwTWuOzEFTu
oa5dQn45ud2uS+vTxfbeOF+/+q5ylyRumlnFox08iBryjkb1M7W5a1Ni44dfElbYn33pftqbn3De
EO4EXBWebOVQLLEMKFEaPlmOrQf71c9LUkrcGyEHmCpa2rQ4Vy8t63lSpDsTEEWboZFT9PZcaVPM
RC89uxSOjsNrrEZWSXQZNTTGANPaI8atCSsVqfYpTeCP9bk7rBrStAcqnGoEg6HwHaNjjks6Izl+
o7dKE727Zm42rOSRz95xSd6F6CkzoWe6LlxtI0hIkkUwUVq8IwJpLH+SyexS0tBmxiRv+r+CHpw0
C772ZIGfFE4yeAWXzHcU69J3IW7LfRte8u5LKJiUcdt64y34E7g71afyq3aS3NcJk86NOebPXnRU
JzwJDe4bxoGm7FoCdvZozYRX6e2z4P69PKuslip2E+UNTN998CWiktBOabM5oUjmdwXsxey3Y75R
z0PfOmJ6tt09JVGVFlf/NIJmt9f9FTIVrjHJs74m3nBxagOm7tp972ZTEkVs9cP9PFc1DlTrtteM
eVMVbwdgOqcpBY3LjimE0ukRHAIWre1XzTOlU3kBaqFscOEBqJzX3wMPP6OCuGt+WXibCIdC3tzs
3UWOZtiEuUzdcToeM2nAh8kwug9ZXiJYlGwUEbeTEgywJC/gwJM2BXMi5vTHthmpv8c6PoSMkGCI
N17R2Zh4XUZi2AbIGRhc/UL+mS5MHZJ/4UISIRvEF2ttt4kbbTrOQt3F1AgEPkedciGarOK5vjdj
eHdcHjZ16Y/64KYdIqBzNX7+Mzt+HuYcsa8yPxQ1RU7K7Gzg++iLKcCQdRxZCmscKoHiOEzp82uv
Yg2/tCamqy3n0kvrqi8Ax51PxQMTpM78da56CX7nApoxdpnXjRnXmZ8U3Ef8NioarCI4lXvce+zF
TNSpypq39TSgIwit094R1wSHMWB2odztH3EV7WN8HjUHzqIBAIRqKt70f7Nvj1OtZrLMhHRMkq7U
YEbu2UEJZxfxt11u39Lo5SipDYBmyqWqjtwzcOzAnpsq5OWIqHsKmJCm6GujW4f4KNt21VsdHW9C
wZf8kW1k3IKcsTNb6DmlMPcuOqn+NaMKd7tqzJtNkUBAnUiPnQ3+lWTbZtjS8hIAMZuvI4M1zxI8
s5saics/GqWOEwpb9bEdMCTzLeW3HbmMBnSrQhRmxvL+1ivw0oy1mMh7+516wwfK8Nl/aW0mEcEK
Dj17IcM3+CTl3526Vlak9sNuQX6Ws8Dluv9PB1tZQfJxEp4p5NOEUZeJ7RvpWRTxvfLAcNG7vTTS
VTZKgzUrGMZ/AsVBU30pdGugSXe0TbQzwYI8YbFiNkJiYf+omqARDUVM1HsfzRmzelY9bpvbt44z
ce5Wgqcu+KOfpnhOIQ4GPGKwMoXJaxkvUix1aMFEPrGNAKzQh4rjfCFOQfwHriyY/8eRayJYe6o7
Mvzt78XY2Jnl0aWEh5bsjuGhlCi8EYDOjyaCT1Rn69RE1+6mUabp+qD2Jd644h3pFYbYBGbVuvDf
zLLKEUsGkiHgklEwngatLMEBO1rrRCE/sk6zXRxTTTlLc+FmqdK+Bc8HdgBOtf8pOpXkmqxJpbuP
3tFbYlNuvM3P3diNP66GSvZd9P/eMFlDOEgVgFQg5Er7ZohweMH3rWrbW6vyg8LQv4+V1UfBWFG0
FSVtKMewLDQ+QTzLxqK9ZhgLamT3cxV8qYnC8Gh1UNLg1jbDKmb3QQM6PfGNiFfZA6BA0AXNyOPK
mPRrWA8WJY4L+5NsG9thRiLNuVmx1ZOV2LUpsBNB4CbYWd02SE8KGbQi7jPaCQfNcxbvHdyaOUPf
rYBMLSPrsOwyrbBsTseoGsCi8YEsuk6RA9GqJzvdK0PGcJLvb2+5rTmtZjNYEipaDoNlN2SPbh5A
AoVxjHnQ98ls2cghLgHEurB+mmxF6xyaUn9sEm6eoRX97aqg5dFxErMhxMOxrbOUn7ArqtgeyDb3
tqe16fA7W4XBwHa3GBPqUvHuZuGMR1+nEh68x1398I4JsTiXlHavtG1gDFG+brJTsUU8A7FXwq94
vEZ8u4BceaEfMlFbrGt1YeJEeFoqMIVKdzTCpAr/8bOYYsybAbQF1WKccn/XIT+iaITeqTX/D41e
d1spfMpHMbQSOH3vQJr7t9pksCHAFOacj3CdTH0QoWMcpIjkVjog8+CVveYW3VMByz/FZ+n7kOSg
3SXnZ6MDEK6EFQqAQzItwnExMKfstBQxAhQItEAaAoJBkV60HnsEoe2ly4o7AKotgXJi7dD1gd3g
Xnq2LOg49QCJ/R5DsSgCI0TWihODs+slHCSZvPOjVTQUgiPSBio6a5HvtPeE1XcbO4sAFmWrlGl1
mE/qr+4NiUtpxVASDBOoe9wQJz7Et7S64m3loV4h6GEemQ6TcuJmsqRMlFHTEviFsRn5CotiAMOc
hJpAuEu9wtk8K/ZSV1n90/JZ18vWbCHPZ9qZdBFMyruSknFv5ZW/LpwH60p+5sAPvHmY5nKjWV9O
UFDEKGgL0rimgtW63U5LUJTm2xGN3dVV5ltIUn2tgDvVV7RdGz8dIjDBDs6qTUKkRLuPVNVVeXrr
2hJlnUvDfIBZ6UPomPgyQ76L/bjR74Oz1Upt45R4ZKWtmBKCbpJWowBf5aA1RAMrACITdVnTFM5x
Wq4inHx3d+pRlMSgAEDwsvtbTrKklFnf7mMVvaEOt+0U1d43xhrHQu3sbbTrzB4K9syaL76ZiNw0
VF+Qg/tub3s7omCZJes+0Bc4/Xuzn4yOQ5DPwshAS+Yv8U5JAcx3xXZmvMs8Yw/mA5mR/6JemUq6
VzFddgyigubp9HvuIWrGY9Ivr0t3biqzSw4SjPpY38IGHTTSuGRTDkczAt1BumdESgJ1msKyIZiM
x/n0efybfO1TkgQxYQN4GmvOILdekLkUKnhdFKH45ZbwQto0hVbWBDKBN83iwIXBgxRMy/cPbkg0
Vwtpus8pCAJofMqkoLxOtv4L+UvzyKpMQIVLTxydWF4jQscUaZugUDluo93qZ/+KDaHDzMRENath
4MO+hbHXCUwfLXshfZ79Q2gX6+1AdGEJoURqIhiFXSz7suSpsO9ShBEi3mC+Lz2Nj3bphk9bDE13
+uYLzyfN5HiIiDiB1XxyCCjybJFluPbB2AFx19G8JwK2ha6NMXuP10nW/sfKubTsZLoErQweWdHV
z4pbzaU9C6DEJ3PhC1EuwD03DSgKOTn+vpRanIzsCEmUEKEE0F+bjpLztShg/iuKA7Xyalop/bfM
5bWkIQ6NohUizCAzUhZoV9+5YRnH3F4nFmfPanMw1KAIqQKfGWi8dS6S7km2jGfGf39k0KT2LIY8
a154kdTFNJxFW0+2B9RQ0N/htcbAeGWbT9XFLOrxhXW5rD0yxgW/5JCu5lkNd/4vZH9BbwlAx1s+
/KPvx2F0MYHuGXjoX/PHPqJLtvKrj4sR/gFjMssUL2EpCrNHomWShDQ9GVktcZd7pwIprb6b/noD
XkisjZ1npf2TzPCuN3LYhijs8zQpeFfb4CPhv2rWKOhnzniu6n2x4R1Gw2aVGexG3hXs2CL1xBSZ
R6+9kVWLBtY9C1sGg5PIO63Yoee3uJghmWMd+L39kRtYuTwZvQQPY3LHAA5dP2tvqjioBZrJEOsc
bTmXPQqVK16cHC/T6a8ON/0Y90Z8bufGcDJ3Nd4F81ULGiuRqlgER7XgmiBHtWTxbnY49sreXafR
6hztGezbFwtDC4enwavduPVTWOVVVoQKhzon522W2lmR+2a4BXkCbO5cmmodQiUxutYjKBDOojX9
pDZ3amPBvpZD+odAHwmRBa52T644zUSzNeyCHuidbk88yR9not1fK1gbHQr9fgM9LJhwTGUt4pnJ
crNAsFg51v1fR0pUt69tHbpuHauXTlvOqRgk3zhzONO1Vci8N/R7ES67EfpWs6VYRJmGTLfcQ+IB
7hve3m5RlvtsrOZYXmeYoaYpWbUiJas3N+lYz3PNPcZNKpkQjpON9jwEYfkMY/lHQzCdaEwZnjpj
Er4bRUojw02te2d8XzEditNhC4DSyCu5TInjYxegMSbjqfejri7/MNtmDfxwnE/9W1SfRoVhmyOK
DoOqemMDAe5XkiYOdZ9zG6YdDnUKVjWxHUzFV1To12mbTH/MPR9EmbhMYDCP74F/HPa2mnv73EGg
pX3UzoanyRgmB0TR9m/6dKQH2Yij885KsBG3DE+ans4mFrgjlvkOGFOc0TzdbmwKkT36R/Hc0/tt
mNQVYTmORgs1UIWEkOu/AO8IlMOFdtCKGDxpHGe0LesBKWMUYgCgNFvNgCwi2i7IeE1/Zo0Ua+QR
vMhk8dUdoTpYZb2yfdhscyR6QeDwMhcVJMcbOdcj19PZ2fhWV6+NwjxkqznLLCYGIrny5xxZxkGR
0yo2j1jXFKvILWePxhO/YWiHddZIWoOyT6FAAMUBiuNhZMu/6fmaYdG7eyJZcTCE9H92h7DvgBBI
q3XNrrCtiuPD4LlHDEeMvT7TPvS5pnaUydsRrZzE/QPjMKcPTEgzRhFxvrveNCNhkmhQHRgC6Dnl
5xKemmKaooqM30ccxrMO6NfiGFJuJOE2BXv3mKsN2dqYK0YVbjZWsHH0hOmzAWtJc1J/qombUZ7k
eQ2jJ5XeX0Y9c+AU82r5DG7byVfG84vy3+9e9aRLT8yMy+FYBgAYOKhYeeqRGJT/v7uEBoFiIfA7
yDT8dVpziGw8Sx0lAFWo231/1kOiHjJrgktiufPGe3/dJuV1mED9LvT9lXpWmFVI5btyVeh+IZ35
O/B/ItP3yDvFRF3OttKujb8P3CHMecAGvlC2QyVjW/DIJWuedpmmX4XjnXh3nILBlN8f3qvg3a+2
GrZihCHtUss/k+eWq3IzP/bJHo0rdMwSii1kp7m+oqKjqYAfZrqGaSDXahUabVFfbpnGofSXKUZA
VlGW8mwtVdTq2Y7p6HVjeaF/inI80vwUgMeNKvUWdzM/7UPvs8370i8gVhsOsIBn4c/Nn7cVnQ8d
mHGmo2zHRsrMVwpOSwnVfAnklpUFzbHYM6sOM8X31cwtG54eHwKnpCXxxwTPyV72hYu+dQQfZjZs
4cYGpNCZBBnkuLXvL+qGKJiUYcBvf7n7iL9OSqHJvGdb9H/yQ77qi9jUYjoAtgoPXO7e/19kXezx
3RHfAcLrDyqP0EnIqRL1/2qaXsgs8yKX1W5MggrTMU+8UH0BnCqNpGYJ3j4LDJGSYz0TQB9OadNv
2e1dR30BQGMnsXTt3lhZaHoD0UiDNgw6cPhiv3Yc8wKgLUZAVq7bi1AHNxhAemOyFGxYd3P+dquf
9vYgFCx3gRhHRcqxvKL9f6gVvk0LnR8dF45k67EVKZmQpMSo1gwP+wGfIMlfDM3QGtjE43x6oCyc
xUnFWBnkaA/T4A+kYhqNpbFO9260O1fdcpuED7ndkncsDkPAuk3aZJKiru3VIiLyfbDcZRdb4WIA
gkPxAWzLUL8RrlNw3hiuZMUGVpLcO4BU0kK9zYBijjYv2uibcWP/+WoQ+yPBdJk1cZByZLKoM3Qk
JblYwAfYBKPqe3NG59I/CWU6n2fowvdWBqUaIKdV95jpj0cpFxNPLDKt1iwptqwS3d8E1XsCyPyG
/BerMcmXtAqDkk9sZ1i0s5p+GacZ5zuVArGFSNKTWoCpB9wkOxurv2e5ErFwJ1//+H9NBTCkE85g
tHxfY03fHSy+bWqVqo+pxS7M302aHDkoBpxFVyvP26dgKu9LZe1gmzTc2RmmFnMVW9+RQQz1iZHR
IUBsZATdVjrCd9Kh4Gi2pCKMwS/PVexjiNtZy0BR7hqEqZ57WBfh9JhsDsXGpYChxEhjI/gtOvbp
f3iV8zzeRQeQvLTNWp18xuZW7B+mECkTnh2jeGB9DdI/bghMEOnSdP53NvRnT0DYn0rrp3Asqcv0
efuci0RDxHONQdV+oNTxni/kYV/VF8np+8zrE3t9bzC6TNfjZ8uEkmlS9ucvD+k753vhktlEy7f1
Wtf0KtiKASVFMZbfspfh6G7EL0v3Igxqgo9TyKFwmeAnu/L0y4G9NrTLPUhWnr3fVu+raqAVu1tx
VSPzXr51Ia35COqgH0tzVWGx78xXoPDLD2bjZlXvxBFDUiPyljbxaItdyP1mHZLGVwVQRQNiXhWd
/wiKoQ/R2a47K2SDIM3mS/P/uK+WlizwaISzw7Y0vsfNVNRF7505+3TD6NeuUUdTWd9A6Dn8Hw6O
yeFcnSw0wcxm0y+oqC8DeMX1GcwsCEy3lgEMKmTJ0IBM4yuxGUXsuQ7MXhN3ueVsAr+IXQpgfP4E
0CWbj49tjAf+QXCfSWuKA9Y+ciiSnMsOo8ZWkrisl8W1OjNoXC6MnsWveRB+lGyrcnK4sWKTF/sS
uCcO/mQKN7nfjqQsUaXpArWnzaZNQLHR2rExwrAXawBAEOnsBGxnUZE1OZNmv8C0Octsf3POB2MD
x/FJMHtQLOA8TUULXjJkc/C/Y/NmWv1TdS13f0zgdc9iEACd8vDUJ6sDeRehXd6Tg99qRhjehPSA
D9pgdLjIAcbSszMYGJwtnkHemjBgNZe//tRK+p8KriFlcl5lx45pm/sX+LVaKsF6jKLhUotkyqiP
hjsOGHFjF4Xf/GXYVnjsyS//wbpKTtZ05ozbkneEzVLpA9rHrTtIn6B6dWHXrs9YmNtDTKyEp+6o
w2lIrRPj3BAtXND5p47aBXNSyXVeE1rbXAhGWxHTF5GdIUWjXsBG0mAwER8FYeDpM9i0qOKyv1Or
JuQHGP5x5dkeWRuQCjbXnQ13KDahaEyXe0oj0CPVmjls7Ze2+z0uxj2PX0UR0A6LTrEWdcJE1l8D
3NHam8c50JZpxLDWVoTQdtg/S/YJasv1ktH/fPmI/6fSX45ZJ7Ep0TT3k+CIkZS96mM3rI6eCH/C
Ic3wnA0fjxn29YDmSrSfD+J333NTyLtv9p7bb96PTUQrtA+A3LdjjBEYlwOtlDsmpXu0OjvFbKCN
UWbqWrHBo7sUtD6JYI1ppV6SAIGJlFN4zbItyROc6PzlnUC3wy/ARBH9Sp8Qf/pnn2L2Uer1Ht6D
k4SjaSMdGr0dseZQLNNb9YWiTTdgMYB9/5ny+WfprrrSuHFqXV8ff1YGGR3hU1sd4DInGMeeS5d0
DlcdQEI46wbE05CFvFyWulDHGopekcPZxQdRSyh3AUxXhxWerxcRkcawBez+t0aaQELe61/D86c9
MKN+tKC14G1i28uvV0bmgTElKjX+SZRgEQUTZYIggJt7hmBApsE5BUI7zRnXIm6OKXgI65KmaPIZ
VCZ3xH48z+bqLXc5luguWtrJ1ncPflTwCpGFAM/lXxSbWBmoEwCRU2DK9H8E9y5FzVfkcNomr/Mm
idO+El2Ww2x1ydFlJkuB9Qy6GZlvwC0VDuUSLbNTrhp8knOAgJo3rtttTH9T4p0cmBSDUl7IVle2
WRpoWoSKv6PsiBSzuqlyOxDmM1gOme+eoQCpJpzCP1HoFPO2NrQDg9SQ0n/OKGdxTqYB6U4SQdm/
FNT/ahn6YpMlHVx1ZSDKcmoU8di4n36l9TRe0AjT7taBNfKdJH+XIR7Crsvcd2AStcV3P3w0/tDg
2pWTevQNlXEODiKo9WhsZzK11dhzab5xnTxaiJYaxgkHkOVx6QzO4Vp4E9fGMtk9UPEk3+WyaQ1R
RsihBFNG7mJ85cR+x8KG5loujj/hZ1o0ao/O/ymvtITEDsjEKAiHG1bHIb7Hehm3ePv+s/ppOD2R
WD1sCOg2vC9ks2DcIaNmZmDXfMHi9ATdLwhQm7GIMsheAolYAlOULkmuSQru7zlXKezLaQO3777x
vpTzpBamSkNkqLvdL7lTX4g8BeE4Mtq9+G5gc2YpZgc2CQHkNdFDoOoukrN/EwgyMliWnVtEDpWz
RYNtpfv5qIxfDTxRBX5c2lPXSwfuvs/t94vnX1d9yPc4bJ4vVA4ZJ0s8d3OeRWEjAj6VC+sYmGBF
YQ6yjYsvYxa3Qp2+txRt2M/4lOij9YQ3DAxIWNQ6afDd2T4XhBTOMM8ZKmmR+MTEWux8LMn00zvR
wrESdNykE79AXNgYm9wT0TQjpHWxlCFnwKjH5PIjc3ZJBI9QYdtAdP0osYCkMfw0PVvN5k1tqqNS
D2Q1uLFtfbZy84B/Nmwtv5KkJe3lJJxsrjn4PbRJqcl8kAS+zjqVzfhrSUguTz+lrIjhQZyYnnxm
8t/W6c/ToCMdCVLB36atA6RVVeXgqHfa8/2kxq9S7pFVqMhRWlAM2LD5C2usktFiGRZBSn1c4n//
AaRdxI18Bf0uGnUU7UU42sl0M70zZho661NPrdL3cLeGLqIBPZLaQBVCMHXAmhKYPsNxdYlKxOJO
xDqaZhbU6/PKlHR7a9YZ+Q4qeQrmhwhx+ofx0X25dNUjSwFs4qSaJPuv4bw1VH+wageWe7RHcKSi
3JAl+3Wc2sANLEq8w+jHIlnHbISssjF9l3YUglj4Myq+geMPheGRHyF9KVTJ4XQ44o8CfFXF+VXU
ha1kwzFZqVPjpBD7EKlT/6XQH4cZoC+167hGo0uT3AThnyv6Ylz2KGmHzy1qhCuP5QKozKV2J6TE
5eBkgtq1PFP/ElDFm3mZzIeX+VVC6YQ2Cfsfka8TuTOh++ewQAq6F4PVqZFxwt/s9gOTgqnk7Jnr
H8OYW8yhM22n2oy9Mj6/Hy55pcXjyGLMzPBh5hoVL57lfJ3uvpVN6pBWkYBjeBRjzubSeu6NBSL1
dF6HgYZPOB7Otc/nSzVbAR/2WazZsFReNEzL553yfBzvCA+M5Iv/WNest25dES95CeArMSPL2In3
Ubik9Dj5qe4uLASlWXHNTip28etL/ZgTLoJhuNmtjRwgSii/gFFhanC3XYp3XY7KSV2CoG/7ITkM
Ok1NTobj9l2l82w03ycy5TDUw5JA9c87QNV+gruO9lXS7qw3zWK8UM+AR45+RFlCkPXrMFmPeYPK
sAi7kyvRHdeeoReE4tsLViZSwq5ivhnAuCP+xmEGGouIdfDYY1xfJbGmZy557zokQvLx0Q0xZdP2
tEzc1bLBxkzY5/KhhC+KVC8GHUjZULUYgCtZ2AOrssII82yz3o85XpHieMRzwN7m997hiveg45KW
Y+nVpyMUklil+JQU4lLp+zsSnRUdXe8Lb6hTwXB9hq2JWWXAbinOJc28FBJ9W801bvCQ+OWuqTW9
+xPx93szOHa7he5Y8dmMj1RHzleN9S6NdfN+yU0DoGs2YMWoTKEXcA38MKTxSZ6BoiMp/gM66ND4
SWCG/lwXr6zSYATSLwfSFjdkcAlEbAwhoTj8bePQR8yuEvqQy8w1lDifx0b/zLESWDxBh5++IXs0
wJN3li8rgHIdptvzvKGINMPvWEA4fg8ftltso9b1ZVRgGQhxqsqDyfPObBrt5m+IbrBJZhLF65Uy
1Zu+EHMnQFS3i0LEr/cjAjI9JmVsV+gf5DY9/cmehPfA+gGJCRouUARC0vnz/hBGBanzkXpCiFEp
8xIv2UCk8xWchp35aw2hhTKhrsg79pmO7Cq1DvSRttGeRfyIM0acYsI/qqCpGQIHObG56pjYMTGg
B135AT/JZTWWnU8iXdPXGZrhMnhnCkbGeWskYRfK4QMTEGFEsPLIywMM3C9VmJ6fcd5NDM65L7ZF
BzAZ0+GLj6rcayLbMOlqXzAunvuGbUfJxA+g4CQ+ywLpTQoOcamdp7M+ak4E43s+KZighFm+e/jd
O7b6U1WIyxgrQ8hShoCW8noWIioOZ/GAd9sscov8Uzr97VxALxUoBy4Oul0svQ6kOimcIlsw7r5j
zP2Fg7uFHsOYzLtEfB5okxiqzHDwBkXjCMtsiap8oQGaeuQ8fqYsc79GJS/DxpToLsNHN6llsS+S
Xqe8uMuWnJ0IKLKZ3K66FJ9RiYadaFm1IMslLW8oiWZThc7KzLffIu0EZ31VF5jtB6sFzeQX29Yd
o9JHwt4EKYLdqPlbEGkQJ/z5SA6z6X3ptpb1fc4TJpMHzqwD6If+TSMAwq0pDJ2cXlOB3eLOi8mg
J0LkGDX1U5GbQZa1sZmKeEQrgAEG+LDe8HiPwjZTyZT/4BV6VfWHLdX42KEdnUTLQS8ZlM25gdAm
C76u0Sg+7NjdSHDSWonQ4MrEraZbhtGJOR4e1IFjR/meIg/G4hFNMlIcTXT12gQs51KGprtdmcLz
Fnv7K6s2mx1ZbqGt5Ra/3550l3TJ0VnQLP1lmI8k0Dzn+PRFAo5OT3Q7N7w/M9EouFQNmekdsrKd
ZwuemoFDiOd82LYnbquQaUjm6sv/I4h9UzoyhDlVtla56/piD1lRsqX7+kRFwUjO03XJSqgkI7Xc
8cpmGj6uRMAfpBqO+xbet3opBd/ACGlcbdlKfZbZLRSvhUGpUjBNYtLIfkTbkJFHg2wpNNvnX/Nv
U7JcrjAqm/oImXG3DwBpqkd8cVQ6cwa+1LCgDV+guWoCv4xIa1D52w2neLbjWOisVaUGvFzxi/M5
Jo4FAUODmaFnjrPqV6Rp1lOESYP+LN/J92a7mLUWtCth08b0GNlichC/diWXjplcWzeM+03aTFVl
D9pfX/qLhYnWyZNi5gG4W2cdC5R2CZaG48xpCau2DR5/oR6sPd0BCU2gO8AM6I/x+z7xx3YPLO3x
rBB0BNMnoQhic0ikS9ZpnWQs5Odg5r5CGcd/aNvEnTHCz1WVyCywQjiABRinLpkrw7cZPFHGIMno
6dHp7/SzjaLbDJrCUKdbDAEAk4MzYmkZHyaGFg+e74ScXP0XUD8VSjmTPdo/df6/p4ZFVuJbS4sT
BKSzsWTJK1wLfIsbMkG4U+Ef9sOc0mj2gutySSJRD5A1Frsyx9gRPugGg2KrBtT7eOkyLf/i1Rcz
zAhVqRT8HJuDkBzclLkfarhvhmJy3nwHScEjnlfJvSumYT5Xdga0OiJ7iW36IVXnfAXYbnHDrgqy
EaTEGu+ln5UpcQstXbKi43U4cPPmhO6NOe6SVownDqgBorFxOsFjk3poSfgILEKVFwM7A2ayMUNM
37ncf7QVf7t1ZGM1JOnvKG6wyi4NE5PJ7OXKTwgMVsTWW0qe8ORfvV0tqqBtFLbgk+fewCrgBr1E
wKQc/fA+Tv9g9RdMe9GRKinXYCCTqfbXyPPb9IfhGqzaSKhx7t3jeof02cDaqdfGKu+xXk9IC86L
vnaP+5j8OeX4tzXX17NulUf32KN0OYzIRAQusjco3T+p/d7mC5UoAYjlZQodIL430a1WF/r0yU2q
NIZ1s+eW5okoQ/KjXfl/D8jMwoG4IlwlN8oIRJwGvBHVhakzfZPrB6lX937k2EGkmXaAPzEmEs1J
DtA9WoW2Sdg1J6IR3Zi552TCUJtPMdo4WTqkN+pvONueiG+PoVqDPErhpO4i9XDK8vyyZBvtgHP7
sq2y3Vh3lZmTCDII5xhVGSmiYhoWz8AuFF/UgGmmoKlY6LUc0tcp4A7Qpja75cuNSeSBsZDdtGgB
CFNfr9OF/lh6dzZagT/wrcRsxteKvXvARhY/TwtS9cANz9SWwtvWVsh2PygPeRjQ0jbGLvWBgEHc
xVd4Gn5IgBzFDLnFZWz1y5Kgg8z9b66rNypVTRN7e89vxKuTLxFG+iI0OMZO6UXon6eUdzEmooqB
UOHNMQlNdysJr0NzLPy97f2d8SlGQDaWLO7t0f5C/XKEugMpXRMK6Geu7Li4AKsSpMn7F/X7NkhW
Xe7/IyIlYNHuc05S9Wr4b+E373gNK/tkb0zkhjjT17Z0Ac688zRQX6+L+hoCzv+QQrtOZMYimNdT
uNdJNnWM+MvY7PBZACwe8BmaMH0mvI/1BZsf8kzHM39T3vva5i63YNwkFQIpQNpCHPlm16tMbK5h
42hU8GbBNu5btRBoKJxATkJf3tdXHx5CPvRH1M9Pf2f+JcGrrLX1T//EwbW159CvuCAuwbqTe7Zj
r6PDM71kCKLVjnbi7uV6kBz/QiZBSAYY+ZPPYwh6+VIDgdLhykZvUv1m/xc9S3/VFRPOPKg0/EJf
ZGvyxqT36qM+b21VGsZDqq3zcCIZiY6wzSk7nxLy7JnYe/xYqsA2Lpj0U150MeiPJoY21j4eRml4
Vg0ZJSnm1xUE2F1DUvdtXaGL79KJk7bExeQpIl0SC3zefN5BEP1zah4cuVTuf486D/Tlya1WirSM
ewPIhdINg4EE0Ir2xqzTWpQZo4hIk2b94yuo9jUodiLky/lvMR+PkjLgTA2yqcc87PONoIZKqn+P
MwTfywh8bWg61QXvxLxrFzKBFjNjQjiWIWDFdPaDVERe4NgtcpLsZ+r/qgoHPYA+mGAy5KNmQfsq
pMhS/Nn5yucYkw/aaFKESfY2crrZp+/P17QR702ge9g0UBUrYpePO6LtLlp4sCLxgS9Q3fqm5Np/
9dLUUgASioOZd+lRRbBVhv+UJCzQlhzWiWey6lk/Wn1PtEaltfKt0vPmcopjLQdzBKWCd/A4vq6R
Dq+EwjfDivx0IhVZOfgpP0k8ABM0YsRY29GuoqHZxrMDLyHYAd4LFPln8hRxxSikRR95r7lz8uv9
YrKf63T08fh4nHm8UaVTisKVlSdxEy0fHHIKMQUygqq/NG8L6tL2dEuyloX7MAlp8C5Y3xh/bDVH
rfJRsvvnjV1S+FsTqu5nTQhVKUFlHIC6KesUZQIgxiNrY87YbuyDZEpE6TYpvOjP+2upECvVPkju
T11GwzYdcOhMyA2emGQy9U9gH+Y39qOxjPJpCQtyFb3bH8dQih5Qc7++RwQae+NgjE8whGZ89Jg8
OVs7mEIIIvXwrVhSGd00CrbwAm/AbdGPpx9cvx5Xm2ZYM1roNNawYWBtbtrai7rj85EFvtYEyALK
IqwGhN6Mbtjfcte2pMXW5+T1stQuQZ5M70UBBT//d6wmMnrHHkUWeW3YBjUp4L6+jQxfrE9a7CeJ
+SHxcuoxyUsY23xlKI+emvlHRnQvMxWwvwcjZ/QeN3G8cwdbnFwdOUX2LzUtMpLj0S6Ix3ngXFGW
sTyvX+pW6h7b8baFETjVZHY+OVS8Zm6mQLY70WK/MJOLFcqwk6xtbfVZUoYjxcikzCXfHMpPAKHa
hOCgUyW8DLpHIecqw+dQZpyrvondti2kO1XQrp6altTcy0tvT80rQqD2E++S/LD+WPgLzA8MxFI0
p6jAgrUSmPV6LL8OW1XHynbtw0nxtovml8bU0Evw1ciIS9rf9KxxHwwDCrwwL0R0SCcDil44hrFb
3683VNoKsBk8P7iCUh58a3VabdNp7jbFg7/NbamINnwXGvwoGdNi/U0F7NjCT02GPRlA4wKAmJTf
zRVVskAI1QVUHMa+49IbVedqhovoeTt+O6KbPTDgC8ojkZP5/QVGpoGaTIqfXl6ziqR9qpFtL7Ww
JqwwIUyUAP4GqgSUEfPnkkrZ7LMPTko5I3EYKCdjlVy33A6futcW+baCyQ3AzTjIMBKQJlk12eYC
NOIFlisClXGdSI7ZZv5Si8Ll1a+VGdHYxpLQn+fbMc7Ow9t12U0EX0z9/e7J3aPfnn4Ky+jzw6FQ
T8x0EmlP94ZuWEv+1l7LrRlKMAnYapuAgeqKDgSI5L4E5W6PYkJUiVRjpFChpSV9I3dJQ3O6HVIF
0rweFdVDf/xx7x/GGyiml1xerUHJyIYeBsvxEkznlC8ho16BsfqUtr1qMnale/COYpjmMhGHNPjO
ceLU7WiKbIHplxg+KR0xZxjJ8hw+31Lhlnn8+NwvxAyehVaSzvemhC7UkW1oMrhlIKhsaX84UK9x
VHLPopEuBP2AHWxkWNy+Flu7734X1wUZ/9TIqWp5MOOtOtTxJPBQhcIguEA0SjXgrRcrWXuEaW4a
keB7bm4kqhj4HeDYWpEAfsU7p67z7XMYJy9JFKSkqEogIAgcA4CUbmtw1gs83floV/TWBHvnAclS
sxe6qUgdzkzoHZrqS9KxhBthi0dUaENkPY2AR6ipTXYreb3jXNvzhT17MiBu0tlgscOv0X8oNorQ
Zzfti4fA3+agudnsofxW/wsnnCwT8Eh+CVG88W7nVndoLbtayZc9PPpkvIhyhElKgfXlEfOJkvhp
J8YI+EIctn4wgTp4OohhS1mT6MoqECf7xlcxccV0mYXKbuxjTIQLD2EgnBx00gFY5KDVONajQ+s2
rd2J8+U3jPRo0WZdVpuv3R+JiKYkivmwllSlKgiVDYp4n/U8G7eVa1BlKUryyK0L94srSL3KEDtJ
AMgcgxmyVUFpxgXCHlRrGWNDjRLxQo06Fd8pKfy0m6+4T7jeJEGS47QutEAQPyUv5sTNx9MxTPTM
AZcy2n6urIq+u2LB0g/nClDtQFVmga9T4Kv8R3ul8YmhN6wbWG+V0XeF0Cm9zRvwupsF4BKLD5j+
iD+EOLcbKQ+IyxRHML9VTyOBtgLMYWFl9mNLosqyVuNsqqxMzVXCt5WESzRK5pc9c4QX77gKgOaV
c28AHDgCZ43hg56RwlHbXu6oskuR31J7P9mqPbR/zuYmnVqjt0+QkvrVeGT389DMi0wp90OLjOmZ
Lv3tTBnFAF4xzGTbXoQtdxMZGfMSjlZBXM2jw5HhHnvxCdHXPmNx6YwSrVTymzMx2l3kAV35nsx7
il3r1Ct89WvnVN/Yjwz8fhIzTKZpeUo5eukwNP0N5LQWl9j6Q79DeexCLBTu3bEhR7WI14dVmdCH
OVc/NlTgRXv/HlNVdi5wm0p2WMr17fpCBDgMKOHVJ3EXedeHTJlRyjk6dn5dnAdx65jnMuoQYCnv
Wp6x1UnynyjQp/QaychP4DPY/stVViOUh9w7XPXq/x5eldki70Uy6i5/xw1RDb7r2E8VBI/0+NZp
wqmE8SShviAbheXS+8Lzj15T1rHaQs2Y8r/hgboBjUrshj9aQPs75+WYVxkcQVHbuG6jC0/Vd6FX
RC81zepzCE9VxHYpWI8c06hMqjhcCLneU/v65GTyETX6f/U3xZ1WS79nkOzh82WUzio5KRNQaCbW
YdNLiabl6EhTmuAs1+FU4W2vcOGDPC122MOp4mDJCmggRT2XYDl9GHkuRKf8vj0NPEvl7Ae6KJqf
2Y+ffPdUFj1yg0EEQFWLYmLk/r2fiU+ibK8pxDDTdoF4BaI1Owj7AO3eXzP0yLalN1NxN/cIeoLH
mZA8AVPxjvoiesxDdsYhYcAObDXDtolfJ4s94m9cb8dKNS/qBqcj/1MG12+OlN85m7l9cCUdgvn0
Up35LqunzRpSCNPnenwdJHGBrprWKeFqSQmp1co/7eatDqUua6eyJQqJMzE8PVp6NAWcfHpRMgYQ
0AE4pNNMXnV81ZK9OqOsgRrgeOGM4prOOukFNa3e3qE/b8Pvx7hm+GNFAqSLmH7FLtMZp1dnnDo+
vmUmMuUcbK6/4YhHOeqJLwmS78Tiw2k6hxwr5jfZnEbhTLmnitWKcvDMUWknmPhP6lQowxHQ8x7y
L6iz1dwsQjWI12wXXgP3bkbeKgvOvRxqjo7Fn/HT/xbl8Ui/S3fCD7wQzfc4Z26BKVF/X6G+6jih
ddTpyhZriOc2R/3trbcrqv+KR5nGQKyEtt7IPBdlE5QutJpYRxWko8a0bTp6Czkkap1UfzuFpvSB
R8DFfU/ZUAMpHWtHGl0LcY5P3IAYfdoIhDossHWiPPU4Z62Rjlh03s5yzVQIwTgEsXL15WuV6zzj
fWoeFhrpBoOX53+sgDWOY40z8U8Zw8GiyD5kbnihvFwPE3J+00Qxv0AXu3LYzr/eZ+ti4FO+L0Lr
5VH1W+pk2YGy56nquWnOBMlbUkc2YP4yz0f2xvvXx8UAiZNTOOWlCJbKKUTVUVk6a+u+blwUsIhh
qr3FoTtUICA4CSC0X59KDWE6/tl26Ncsx0uc2t4nbs57l9cG/4F3XVL9URt+HrjgZZa3FukfqVma
NiHU1OKH1SEAV1eC5VdyL1tOSbzsuh+qrCRfDnrlDbqz4WWVd4BwpRXrNBCCYrDUvEfV5iDFC36t
Uc0Hd0hxCfYLeF5dh0f86UdV1MB8cxd3+uD6QJavTqj4gufupJ3sOwNm6ZJQjHXC2IgD2EEdJDwp
rd0BlfA1qY1OI8sdiS0WcY2efRU0IlyJ/Q+CXNj/LqNrGqHcjaxXVfN4KPj/1jTUY8Usum4/qs5H
QMRyBP+OXHUxjslMi/tQ5Fca2EF6vHsQSOJACnWbJdL4cdppBNqXsQpVxS852rxxYFn7WWUcGXgt
pCU+6zm160gRc36LLZADl7e9deMcG8S5Lp7QBQpYK3i6AwjLtTttEolXHfGinWIa0WRL0eW3GNPd
OmBSn/czZ/nPk/vHBePCyK+YQBzHklRuZHE1bBcRsUlpzOKBQSLZvl17IiLPpBHJfygISIxH0kMI
6k1wpyHtngoRBjYeJEivG8fIhjDbxKiD0zRR5yhbozDouz10RXhX0sOqmlyqK0wK9tUY5i6UNJ7Y
2rbuZX7p0O+h4Vz33WYHtVx8mdwIsovkUcE91xv/n/td2UNN7hsR1d/ghGhvEZMUBRitHz3ugIqY
6rQlxq8nFGEJS6somjvsymG9hqAJBi9qi51pImVXBKxiQyCaUIBJhdKbGn2zf2nSQFT+pAZWSmKZ
mgG6kFUK05fGpae0jZNw4wLehCcKPAMF2T9hg22chH8owGhqov9MVqfKg05LXGL/bBTK5V5rnqXy
RnX9x8QNVxUGiX68o93GSZX3Y/1r7IGyZXj44nYLJVWO8Nls5G67LZUjEV6MMZIRGCQQenxkmFSJ
lb8a+gPZpM+tWVmde+hTIx+1yiN0g6OTvC59yaqskKcJzM0t0iRY8mwV1Z71ecnRor/pHkd1s6X3
knDP2qt2+zCxEwBKv0OhJ6B94Hs58feqypzCWniWgEK2kAzVVEnJld+dR+55fNUR+3SPyS5728Pz
LHJ68Hl4oSBFHggMG1eY72sHR+su6tgCbqKV4nRUzdVjo21isqu55FN4UeRvngDtl+ym361jRnMk
4x3WW6otH21P4qA/qTFJ8Kps0mH1KtovyW9p3IWHcdPjJkUOw70V+mu9t85AzhMvFYT17Oi17nTy
+nu2JCbY8Xt2VNaVEraxznWmg1li8jswu8W7S/unxTic5l3nhMA3WCyYnPBQuP5UYm0h9JYgEex6
QzuDto9Iyx+lvucF4sjSsf5yBlzIOHSZMmOlxBRELjdowWF2Q48Zc9n8GGn4CQsc1RkHC4DbTGwg
iwpgRI+5qcmDcfzQBIqCzcbi4gC9L/gPqIFqhyGbveP0VBq5bcmON+k8qHQ4CFSjzcI3ED+dEM9K
5uk/QnnmxLQ+gX+LDO7xvwQtYr217lpyClkL/lvTFEoJHDd7PVyhEBE+xuKEPsNhwv2u9h1M3v6a
sdOLEjWc48c9DpkE5oYb2sgGyFewfRi5/n3W9Yj2PlQMmriJsa5Spg/iC8wGtPlFjYvJ38bDKhY7
ORSxqkjktdE2wOiKP9ZtRih1q28dBmCltbUadM4SZZq0baldiNLcVrarB3c5/lZuSECPsdP+S3EH
8J067zbNNhY+ZxMAr9pWHYMbIF3tQ+1R9ngbHXT5A/6YLIKWZLYd52ve8VvFabyUOY/Qo5xaKWI2
S3Q3FBmZH2FbLx8PvG9El9GIt+cxN5SjNJIU3oMNoGT8EchVuLWsqSDhhTEE/O7WEINemDtTCOZQ
HSgtXKMln+LZoWpxs1UZWAmoXomKh+QkSRKD12jatwR+5lAzd/Yx7t9ZKmALWDBX93UV9K67AkgL
kwkYqFzQumN7ysANsNt9sKOG6ttBNKWdvsFyFX/6OVXuNLWt34jQm47jTY0V2f4Et0L2xn4ovHh/
XByArjuqM0g3cJHe7gWuM53hcmDbgWAZ83iuu/6daPj967a2vmkbYs21N19UPImv1eU3ole6kECs
Q36+3gsa25OgngULTw35VUnbbkKP2h6Qj/PwkmoK2oeC9egL9I0dYrfBLrF71Kiih3KdPWnethQi
fzG0v7Z+hHl5Xvo+o+nRpZ+lVMjKMut4vs3PK/C4JSDTp5XCEWvi6zdXyxAINCydLK4VzfSvnNDQ
G1JJwlF0N6l02jz7hwbAzxBpVwpk7Xw1+Qja7KvnIFTnGQTJaVleOmjONds8lp2AdbG10n0kAAgD
EsYBGmeML1bv8ncwl82+x3aGHPL6PRtqHqyqKdEMNrsJgbQ5vUDkMl6GyNUFTx05QbUrbdMgmkNJ
jsQA2TkEetGU0JH+3XlSfcCWNkds/CA5HtvAU549T7ApBr923FNEbt5fb9kTFWs0seQpx5fWUDQW
BegNPBUUwT4k4X7m34AP2/f5QgX0UgrnjttSZ3PXLaoMxXPRYFoDwT6kp4HLUfyNIN7J3mdlMBqU
kX+BX/KsxP4f6Fc/cneUQ7I2Q4RhUxzUpoJnCktJyLeIKIFFZPEBGn45DFlGZWIfTsI1ajWznaQF
V+bJ8Ihb6IzB2PZUszV9f/ceobqDWXHkgN/h5dRKCo1JC5Rh704K5RoWSbAzHbuv+yCXM0HHg5ZS
S7sb2G8DqdkHIH0ZFgC/63N6ooEbQtz7ySb8D+ZCscdoYhu6ab/qP1lR3IB8aLYOMuo0YU8uC4S9
6dhGB82My+XkAkPHGC8KEzql8MpQIGa8jLUPbu4DEhcM4hMI2jB4Vq7lEFxgrImy90q+BNsumEkY
rAPSbAt0NYPWcgez9mysiI6vvkUn6ioVyNfwaBKcvVKpa5HT7JoOf6n/UlOHUp11ccSeHYilVGZR
rZz/GiJrA0IVo+C9eaQYYiecZL4hrFA+tsJT964MfGannyup3rGwr451Bh54eemLCfSOR03cf8Yf
PUcIRMNmPX+djvsBGcyCTyNEj4yGCnFZgxCirhKO9IG+cdkF4REyK7ZbzTfysb22+Hn6RT/NzLeo
fq3CLPdKK5cdDYXZLV9IDZ90DsYs+/P3lA4WS4awz+hSY2/yAIgwhxFrtJrAmSRBgVMqfLox032/
1B6d4n5g10YIfJESPvu+cryRn639xzE8tbOp5BEuXKgWmkpg4MrnbbHtUDclKnZd7S7tHkT2CFEB
RCOXQG7ni+Lq6j07ykP6PtSIgIsk1cuGtCumigltVaWEv+bJk+K92LCRmRhTy4G2oz5gi+xvgDXm
HVGKrILFagmEPlTuIYCxGkRgHYx375XWdxbslN/llDyret0lKdr10+b52J/cIcGPfS/78kyZIPGM
CIzVeU+K4TI6OgcOidSXEWtJ7ESnWeAjkxC7+n52N8IMvVlU6XRo5x5WHP6jsbowt6c5i2YD+qfJ
6WARrPXNmZcyN24ppZGPhvRfStVhvW/T34A9sXVEvooKRJAJ/lwPGyK6BQB2a703aPIvJxeX1PGM
OAsxNQLQOAdel25Op9E8pFRl6e45aEG1WtLbG18D6QcLlbU4O7BgHL+/QlOOxC6Cz3dPc49+qZAn
pyvSGxoaqvNkX04x2RMRHo+xuUQGsBL+lS3ofHhBj2ITXCUTKTq1l/dGLhi1jLxPjAa27148pGFC
vx2x64NIbLrnPTLleXZSetEundDu+GlpNwab3mALIFSNTn1iAgLZFZvQQxGi7YOvw3PyfCI1Eq1G
xCe7RY3cnY9BX6R+9zZsDyMsEwjBaZ44aq2t+PwAiaa+UqfdCqU3Uxbs+OMlOvGUgPx2lqjZFblS
EyNInWjbYieSbySqfU9eFcqqIfAOKYEyhYdtkPFbc+19KTDVUqrzTEaoDauEfybTN0hkr7qrQe3f
qxXUsYffDilsN/bW4ioogcA5CIozCH4LkHI+ckhBks5Qd/VSbmBVsiSXutYYS4tUmCk8vPG7kuy6
RVgj/AQ0f77JoxNCdRQyTTuFMiATtr+LuCTdhbg9nMMZgMqs/WTxJk3RW7A6+2YDsNZRGtGPsMfv
soMS3SsLS2MwhRJyTYmQewpYs4Gm/HcE9qsWNWsGgzo26eo1dP+zVTvbb+N6EzXneJkPWBNfgqDH
fuVeNHD85wKDFR7B9kh5qgAjD/wjU+8XJtVVSoeEeU/oes935PyfxA40xGCTQHQI6DCqoho+TIFY
mB1JueozNihcZHHIRzLnps7knjnsRngGzkeGdteSGTWJjbZOkGsycPZVfUUXLq69a9LQMVkYR3CH
vH6MF1Df9W/UQa565PzRXhk8pTs6d85FE7Th2insJramrW6vsw9GK+JVEHGUxjj/jCWvsRVUJxpy
iOu9t3LwDKIqZvsoYlfNqEPt4zOVMpzHSQGKRM1UZCN1PbbY5WB4b2WgzXn1euQD3tDUa+0PHqW9
hih19cYNQvWqcUEG2OFqzmx7RhFRYW7Ryhy5z1yN1bBG7Ut4ui3SO6f6BVqtzE2dtoYbbanOkEzN
BLrjrOvthfElLFUx4kBfQr0O2gzxMkm236WsNYVZbotbVscbjICxeKrzrKjBu9rhO52e7FlRrEyP
brRVRffCP2Gwng8+vI0XmQOTCoapWegLlDgdcLjZtvSX0V57ImGaJxd13YTiYR8PuArCUSf5PxUc
1CGLgmI0tYiNq1LTZ6RbptdJdzoHC0HnzVeFQwZMy09l1/ED4/sDviPs04AQPoNDOCnpXA/qlKxs
cRTChEgVakUzgPdg8C2HOg8tvncB9MbWXnr4tBNaTcimHx/2gTPfafp2kKLAgCEndZ316+hW/HL6
W2AtAha/eZME3uciTnYNATXRP0aJYvOGixCXUEPZHNOloI+9oVpcvtBAZkxmdUkZtHdaGK8/7dff
27jPiJu+pNaYiE9l5GKHKl7F/ih3lXzGEKPmL1eTei0kZ4DJmEowJaoVhdhVYXrYzmyW24tP0xAj
d9QFtfdBRdvXY6wTNiGRHm/1RbDmTfSHF9hJpRBJMJvZ27ryVVbjHPh9bkBOBEUE+frYCWUMMSH9
ULaZtgF1IPBzckUmIg3+i+7Mdv908MQPrJY2erZkI8/ZRQYPb38eNicTgmO05FMmMNpjgxzG8uxS
AEzQO+7yLfqeNXmop5EtThU10kokp7BupfPC8x+h7LeT4sfNt85eWDSx/YTIbDReXu//wmF3phA6
pk5Za4YK1xtSpYFeNfAy8lW8fYAHGMXikl2WAV7dJ+cwZFpjMktySFIwSsMvg5y0gCeOk54eqVnq
tgEB+alz8su1uzWZ5WUuGggxfnea8Q5/BqeNK4Zgd3TOo63hjYrHK6e1QyGfhp8EoCYuEsSGws9/
+eMABahBw1sRTwol6IaVzIseYeqtc8IkKbMMCg1YzPuJffXiPmknOXXIfjfJDPEvEGHYw82jFX5f
9NVAPL4gYowb9UGezsvLv4+Ou+MoA3Yx+fWbd1FFDDKIBbCnJBMLre5LvGzwtYISo0MvzxKKi968
cEJ0PCIV5FWeVUYRBbdsbqDNcpDE8Pc0UFajfUMBtwnpYXip9k6dwuZajZdmYQVaywTQ2/caXQpJ
QAcyRF/9ZbWu2DSgJoYvZQHpIekQdsz3Gf0w6wXeU7rQaBbKjw9In3EWVi8+5jEkSN4XSiH1RJh6
bz2tKQJ6xs33FqhZJPlbMN1aW4wCSx16vAe1pZEhSgs1bwVjz7CVGSW4ScPZlc5yuz4ixxhW3p8o
JS11oShn0RIuW0MBZ5Cc6eZ8oTh9RaZpXnj77kedjlZw2C/BTtR0ATWH5PqjPLx9InfMPXXNj0Pa
1wwwkmGw0NqozFtaP34e5wmuhkveuP8UavYfYBMS75uh0J7/uFeNCJiTBOJ3RI0jibqxkfUWpbqd
A6PgAwdylRmUYK5Z/FufAcRyBpc07hXPGhN0l9uYO9mB+lrKojxJZ7S5zlagmRH0qQEFPuWlspop
BA/01bEpY/2hwqTROJvcmi5PnAVMICNEYq8wLeH3ANh7aBE3jm2nw6M6LNBjesqllgNC53A8dDSG
xllnhWXNPXAqGMD/OBTZC/YU06Mii02G/CmI1Ph4CT+UQUQ1gTht5aFptHp29efpaXVcU61Ncnis
0Kn1B0ZO4YXVoOUjhk1ChUqDK04Hl92HfmRWYXNYUkkjN9o/2wzPm1siB+oLcwKv1k4JeJ9AKzHc
YnhX+paPvAQlmVsa8uyu9x18tPcAp0jaRdkzj+4i1x8cWCqkGiPIw10hcV0ZmwRrx/Wyt9EbRU2k
xAExXx9gZMzLm9PEssTkL0VXXtoUFJy5ePVRK2gakJcuXlnAhdFfOpUyOu0iJ/EXaDH7XWiJauOR
uSiCEcHvmlCQIF0GCcJD9x6Uz17IjuYdQwmb9LGBz3fBKc6KlgUw5imKZAYS4zFbhUMH81w2l5td
9WFmDo/qMDmftIQVcQfOad42y2rs4yGzdQRO58K4Ezg7Yz6BkLZEJ/AHmWvsZEuLji1rLuob+8cp
1iqP0jBeC01X8tuT4ATlOyBPOcxmSRQRfkiMUs3GFMjjM8hqPJzAhGh8cHJEywRVWGXbpWFyXI6F
JBVjxT8UE7JBY2ALgbyaYv8VvQehTOLTwflcvC+forEqW9kLyf3U5kARK2oVsuPM5BWmrr4LxNKr
nkbgxYrxDH3rba133tVXYJYhbZGMv2sg1q3KW1llVYQFzBRHgjiHllQECZSLyp5JyvrpOcxEfRfr
+IFbKSFJc9hBBex4c+EqzRTQY0XkgDkTNEwwf5Jp6O0UFhdLCpTHKyGHZr6HfQgCEbCaNM8Etthz
hfFLM55pGXJSJJii5+uza5ekvH0I06iX90sT1f1M4nVrVF7VPOYRHF8P335hzGut+0HLaqo0Qr9O
JyeXBuqjHbtcd9ewCmIm9ehaPzRh+TXWksBrtXZsjK6VO7Q9zyXyEwhAjJYZEZqOL4i0m4hAailN
bSD6WhrUjYEvooVtbMLgi45c98gQtZG9yyGXYIOQJuZa8TsRR1ftFq/x2bhnx7JYoaG51g8NU/lq
YVErFEcQKaF4ZX3PKgeN7zv5ZBnA8KM7qSrqaOn0GISXSr9TGRVpSJ3lBFF3tWxHd6Nz/5ZqVQ4N
7RL/kDAv7gZG3WNbXGb0Bm+JbNqYpc8WDIySt0ARvTdyumwX9wl25uqVS195EoaTwN0HPFFDaiF6
JZsKuLRv0MYoh/NCgfsoSt64RGszmu26VwvTlmmvt36eKSMm4/QROwk3SCMHS8G87ooXhzj/PnO2
knXQGrhDphgdyvVHbubRu0VrqHGyJ+1us0+sM908oeX/Yt55B+6T5KN+iQ6cymPgQ2VN6ntH/Em8
Zke820g3HnS8vewSM98JVTBzRmVSy5U/xiP2sRl8HGXN1cB0GJXpq6xyuILiDKNBfRRxHi4QUvEP
oEjR+Cr0tjVWEre9efSrR0o1slHQ7ZVc3ChIwRBZbijPfeCweTb0ZMvz/3jpZCc1TZf1KWat/ACx
R9yPgmC7urYYzR3WC1hAp+9H/VD5k24DjqIKJGoAozXuANXbeTG+lmzraykol1GrIStDNNqN1ROO
kcvE81LNC6Egc5ykfwXPXxJbcnP1Rsa+f24syGgYxVWIBYc7QQjiTNEHasbuUCAq3Xt/a2kIeusK
UEKx9w6OEs9sNDaYCvJZdl5I/6YadH0tU8rgOODSQPa3GITdsfqYenJzI4lN0PMI8YBG0J0KELN7
j7JrhOVFUAKFu5M1U6oqrc9jUUk9Jh2Mj7j42uSMtPb0Zotm2vQ1veAf+2iuNYQ1AMHbX9BklPRS
6LzIKZv62FIQMO01xpvLwS/mY3dCuAhPbu0Fy0BR6pm3gisbOphPHnfM2/fKdm1X4nqMoV1aesW9
Fi5d44VZQvJLb/mXU5IBdWR1QqJem9HQyf9TC6PgE9sYwbodf/BqY22Zn2lLuULOC/x0Knlqj6iE
VaVUc+Yyv5ZdBUEIOTerXZ/r4UnnGfKK/QAKOMQgAb3WQAyGpPeuWnuXteDZsylz8Xpt4tO1kpDl
hK0sP0ghW3AMUk4pDYEBqPDqxOovi00PdhRFgOH/2wpyJ59MyeE4v0/m2ZFiFlkKCocPqZtVkJfD
a9wWGK/c8SgPE5JWlYehrCNAVkyyED6kPBKjc+YfuFcVcAsorWNvZ5tGUfyWaQhoYQp8a27UXW2n
sv+BbnP9BjMRBB0NmufGiVbL0UZNFfIxVYQD0g3eXU05nrmSA8a/4dz//TX2BCmXX1uAbZytHFDp
BXuCiPh3Jw4zCxf32DA9tI71zHTFmSTzAtL43i4LFOHIjsPP8540V1L9bFP+WeyIL36dPr9IGkC0
1Sh/8FYYlnffvl+5Wtx/FvJnJ1V86VuvXGubjJRannla7bhs1ueCYY0gBw5HhjLPk8EaBnDZDW39
OFZzTix5XgQfyaL2EJIAI81S76akw7nUqA87hXd2Rc0yl8W1NdWsytSqR8vdH4CwskqEo9hyW4bz
bYx1u4/yEL68TVzZ72FpVi8r0kNj0hOfcXO1sbACrIaKWmEaYB8+vRIm7Nd3N6Lx3otdcnFE1dXp
MtGPdp3L8wC+S8Sq9/YshA2wzALNnfhZ10+cvEzXmlmmujejzXFRXJY4GnSRiamz0pQ7Lm5cqhIY
PKG4IYDlf6t/ePBtzAOJEFKOO/jWJVjHB5FcM2T2mACNeC1Qm0Vbaxdn+gU5XtqQ250CZtvgNWlq
jvHWJlbCdPvS0r3qk0kFz9xgdVIl1XKkoN7jNXJcAUkyRNlVP1dj+OpjpsgrbcPygnCP2Jg4Y/7M
ufbP5hJ4KVgqJMd6hHTQQR9WhNVz/V1VMt1Zymak7yfQNQ8DyKtysgZTApBNgyiiajPhu9P0jaq2
p2KiBe03DJOzFUJrwnR3Rk46I/ITtS5McK1Ht/kumEc4NEcT618zUAb946i7fOqqtJUrKQwNfocS
mWjBC/mKieh3F9nVeecOb5x5Jq6IUlJO0oL132hKUeHrH94vE5s0Nz8RSclbh69JLWKMihCRcHC8
AAz1AvFfNO2kvwn0Aw6xnSlohmP9JffmnHq+yji4B0Smf+onXz+A/HNAbDUG1ATx7OcbUDPR/c9d
n0hn1ySubviE2h+JZbx43YVAdFPwohzP24C6EZaUyXiNG04MWDF1/an4LLq/+yOVU4plnUWT4sIe
ao1HR4jwmHzHPMxSx8PIppxwrCyDqrr1s+UugLE6m+lOBO48IRa3reJZ27zPBQ9DFfnKa351zYt4
bzwPL19Z+taDYUA6hOMm9+sxKCFqfvPgEucgqBRFSRp2DVdWV0PZCTBc0Csx/7iKbvBiGTWvX4Y8
2sGlviljwSlON+E/EV1gsmlaqXo3SGxpRGqUvWag+yKQZn/lTHghOupLgwTD0Rc2WRvJ6u7Uv7Br
EY2SmzQgwSDlP99VJkzlorZDB+JBTJS5Hz6saNPaY7RrQ2Wb20/m7hca7cmJgDyEyDkuGUYPXyz6
KWYkju1uL6JLCDh274eN4T9RKaugQrExqoEpE7n+xLHYc0UMahwSEBb7De4Ba3QBWuStrW9XCfE2
jzgnAK1UwuzUmHpyxaLBFD8rHCjoMkgFRRhvhseAQvyvB82FV9bzZQqsDyiO3HVVHnW7C+XpxVXI
1zg9t0BLO/DQJ48PK17Y5fZLr4XZ5D/qrHy2KZ7KEGUJOher4H64144zJRbvkc83pcL5NREJeKWv
pK7/QfE8x0d3dVtIr4a8ayOFSThDoA8I6wfVv6xMFQgnLwOsGZmDC/N/BqeZEF/JEVqFHzSa/gRK
YTZNvTETBPzP933xbD2jdbBqVkLh5Nn0MS/D1NIustRnGTGjLJcfOOWCxWqlvyJoC84/rGWtJgFw
+ZkqXBrf5JxPEGKc1K/hrVAMVSV4eIlNQ6xGG7ok0V11GcxJw9bnj+c7+N9z60ipqZrTbXXs2zFl
7Zd3Ly9EyBf5XiiGDP9JFxNsygK8uKfbU2moLU91yk3UNICDMTUe29sb/or2yTHoSbHEdGu0gY5Z
7XuT2HiOpRwR/7QzeO66fEslbqvmjAhe4ldWJrGUM25k6f+K39c/DRxmOtM4od/hCi9lf4bUfaIF
iY2mxhHb0fjulzEaPJPiAN/loKY8O3jSgnIoGxHIuIoUczFIylLzRxx0S2Bk0W7vjIoLWCcH5E50
n38S8fX5Uu9g4tU9/fxefUAPp3P1jJXOOfhOrGhBxIY7LCchSUHVwXIOdsRAitu2fYlX/ULbwERj
2vjIf09nOcE2T+nYY1ZJ+04v0KBlf2ugvcFcAUeL+koll22/f2RfMonmIgJXr0ve7gc6keETLRSK
p+lZPOFmAJvXwNL2fhXcfQfttzyh0hKcHPU2BljJlqgELR8+kL1hiGerX7r1SJqdvRb1oTtUeDZM
bAOC9s4jHoIi10pUtB1RGkhGoFbngEJ9lDf2mWFJmrRXiaw0WVvTpV26Aw5Ugx8xt3wxP0hX0hJr
PYiJHceVwV5yU46Un19C3KRmgK37+y76qZEsId0ASeL0Gb7yGHhNsy3j/VIGjli7cwDI5PYCgRHI
DRpKgxVWIxbpFT3HrbN8scWn3IvgfXkfUCmPxS2xye48k+F6865IsEfAKTiZMyOLpWK9YXY91ipa
MV3h3/cLQa5P+78eXSTumDCbuyY/x+W0UaJngPXULGEBI3PDu5qL33wq+G7w+bQKZ3JW7HhzT+xa
W5R8ACFp0vrTnc0jKiKXf6xWO5mvQLtKVT+TXwK7VOnoBTL+ojtopLDOvOGXPOgzaBST/daJYiJX
iycMc7DHaRuzv4QodFzRzFZ7ZUuReERaGVmV/G8Vy8oJVO6z+sdPA0NVnN5XL8oQ0w3zS9o5zpfq
XLdVEDT5X1aa6c6J2IGqVVWKgidS3kRgdfSXDBxJuMd0WbWELbuSV61tIo1uIwPs5IobWtsKC7ks
gZlTXFZMTxH8sLJErpjydbNn0oAGKw7s6r4egbDB3WALuVTtkO+Y4C0OdLXpMHjDqQF3ip4f9xnu
hrSfUCSrog/tIlIXKrAp93Yan29N7H1sFw/DVtJQNrlXoZlzUy8juS7Fio/q6cRtsjTMmSE7wW17
4hLroR8AvpKkieKgtvCW/7QFIj5GJD3Cs5Un0M8GvhUFiln4awcmWltQc1dExL3fGa83AkjlLgV6
6o+QIBAvgxqZPrq8d8FsYadFcpiLg4iIuCvNHXP2WLCbZ3krhNp4UhxTye0qTFMPc+Blz0k1E7KO
1mUJ/LH9vo+jQEAVaXFk966LLqIaOj/cXe5NnEkcXqTAZZy6nJ7taSl5LSwqOq4HQ5oMkqfN6QkK
n81rlb7ziafyKfpnFyFtUdz04qkm9sJgD1auXIS0jFd5P2Xkn3Rn8dpqJzxAdG0flFv8NR8IUchZ
+tOaKupgyzt5QudfYU9f4K0T6Rv/2GGyPVFXbUz1XK15lbEooPrleL/pxMMLapQ5cH3xV57l4f4g
7EE3Qw399l+dxFJys/II7KkLvYTwN3P3+lGezZZkMO6Uv6o3M4h38bncUycDOJcVhUT+5+QTQ/xF
I7qEym5816ezsV5dSUG/OIzMM61t/pw127No0Ly2B/JYz+nr6k85+cabWheVtAM6Ox3Qe1INuNJ4
ogfknS1yqxav0NZZLjgRqm5G0bOfzwI7EsjA8IzRCs2RN5iM58L/GKCsTibnkO9zlHK9iRUfg5nK
rMj97jtvIiMQYlWWHkLDDfqFDwv3xHyYVmNM/SZQyGSZSms/LJ7Op0eMaTzBchMxkrh2uudkd3v0
i8DFNiWLJYOf1AyKV6TdWEMRKNszjKK5H4mBW24cvhknMlyTM9lrMeD/KAMtAFvoROdneMmAh3UC
HKupsoO7zndlfG+2+RCN5BOXwq34AaL7FLfGkenjxIuzgMfdWzBqpSOgLr3srM2cwF0o1LxTrPDM
KdbQm+xkG4lEjctC0nAJ65p2J9Zbozp+qYA+z/0IUsXCApcBW1UAOBgCLlY/6EADJ47xHSeLokOj
wodbREzFlYWW4TXShQEH0p5Lp48xcUsNaYhqRvnYNv/TW0yY/oTWatJRhsTLE2twO8qTwxk4PZWW
tXW9/nfZ0vW5AplE5Y44kZZIVxlo+aZyolWUKm2K1Id0JS3H0PXAIhKnwu/hTIQQVX2bvg0ksPgm
K9eh7Nh1C2jN5gNTV/MjiI0pxQl+NAzo3/UH0qm2kdjRf33ilT5w8KJv83Xn4WORF6/DjaMa1fEC
YHYocQ5BKmCWF5VNn+ShoFuqPvRFEHg9w+ezno6ZJnLH0rW+I2+iDiXc3537EnHATKs2h6Id1ICG
EL9IyywvVNHQGrAYuFcqpoU4Hd4xy5L4CTL3T4dg4K0ClETmALInvkAvwtbmGv5UWzxzP9fX2c32
luXJr4w2sG7JZAldCShe//MR5AwNBuSQhxTN7rbKAc1Ps9V21xF3v5/WPThBDwamqFv//SsKtQO7
uSMpwp5EIY9PVNJXLsHMOWmm1V+w07HknY9VL9iXKMQIcAQB5KpyswgsqUuAsj4irgQ8JCdyW23b
h0O9U/x/5llkwY6By9T6Y7dTnwZgnkVmEi0i99rDyipQGrAV1wbJzIJPlz+xai0pA/5AYbXwELv/
U476pvjto4MslRg+lqD8LgwlbUEckJMlx2FpUHe3QVcAI5CGhMhJBg3P4wMimbIL9qWPVm2lxSqz
nSeRPmBCtyq5PnwNQRl1sPyY55U02viWYA+Ota3st1qa0BE8dOKBc7r5SbVtLaoPu3y2T3Dmf3D/
YXhfVbWi5mIEhKsc/7y//JE+Es/9/aT02rEx5qIZExthC6IiIVSrRL0nATgqYm6xUwg4VVw2MNDa
4FAEfeUvW2Qvgnl7Di7g0H1s6ysaCrEFxHpqnvI2fGpOOt9MDIozQWHn/spXgyUN995KItKLSyML
YdaJDaQNgkj/bcGIUKLsXU/HYZitMyUuXNblGFJw+gnjZ5DGdjIQG4SeeRV87lfviBDvwvDiyjCz
mPWBVRK1Y4d4O3y1t1Z652KL9fP5jRRqvaN+oFcdPleRppMGwK6gCDinvg3h+pPXqfKrFj8S+Mht
jIFirU9WzQblJamk661hKVqTvAzxHdwK3t8jmjgnerhvVsHUYHgA1khkdEfWAB99QvzAa/0e1NYO
bw4o/LmnC/Haf7h7rWSnZuCQiPxWmXAE9yQTGohHaUzL45J6NQUsSVodMV/fZxqk1FicwsbPlWya
aTDnh3UXnbOWOcVp6fC04+vre/bD1Z0YUzI4Q/bGcy5EHTmBC7zIIVF0f+eg6ac4XXAHpqKYKroo
d7FLc/3nLYCEg2oTFxkdiI3R2K/okgOys0Hw1j4BU/hgTxzEMNXE+rk38sjTbipjZv2fxvGe6GwA
WXOdGfzeIrVtOEoWwaUeP26DIT+tyO1xNffgI45pAR7k4UAQNYI+L4hWBG3Lu7zSDQeeS9puG16/
vJAW8UTMvn2PYVszZKICdGwiAhL4Wd1VkSyBO2H7hHkIbZMGzIZqgeqjd+ZMjYJ4YfGBQQoUAa07
uXaU4JcdICy2XL0oQdXdDRFtwhnl+cKwjY+CO+4wM2gCGvgneoPPwxPrTa7EiLTweiAWppZ2aQVg
5IAnvwuMfA8J2RoVAO3yDxbiGRyhKmwYiQCk7HNTbBK0ElAM6Po9SKInycAXnol0brpuUW7Ecn0f
Byfjje2U38GZRs0bUj/hF3ymIPPDOTcNRpZvGJtU3uZTfhXwyDyFkNXhk4kv1QMf6SgkJJxDdGrR
gMiSXj4K/q7Qdyla2iwyzozSrZki3OM1QDUt3ElLCF2Dsc/P+Ppex/aURg7HjiU4TsZZsQCG5HLj
Nds6EHrzfzW+7myNsNInz5prqOe+wbii6uQSHdrD9LhE7Bcpyu+gBYX087ivDiou4lczFacz0YpS
VCocFT0G6bNk8GzHAlSSlGHfpK8ExYshEy96GiaHpasLdM3g9I3ed0rx+LXzdUntR0fLYORaE3Ae
dEydgxRilmFlO4iVebN8rwT5+vf2W/jKv4r3MFJn1iEv6RlEJfT9ehY0yLx6+4Y6SctbUKyIv/N6
VfVnSY/cnXQQxjL0LzHzR6sZF6/QY8QhQxf8HBjIWf1sfODtFOMZd7zu+cq9ywsQZH4EG3w2J4LM
zRv8D1WwEXvNqPG1vshE//MpPVJPRNRK+9IKNtcgZwHe63ZFhsTVz/NfRRLwzU4g4kSzNGjoVC4n
AiUKAoexQG+3un4SgB713qOO3/g6KdGruXEvhywDMlle/ETqDsgDmM/+Iz3vZrB3bArTY/ZVyPia
DsW4GK2Q7U3/ro4Z/dY6AhIbveLNv3EWW6aW9B4EXyHLoPBKk2UOX+eLnJYUiObJzcyH0zVDdPuJ
ol3AWwDqqX3iofqabBjOFaW3WFoc5mchYFGw7FEI3833gK0QSa+0wGNRoK9711KwMOW6xaV8O+7H
Zd374o83BMEO5hyINu4MgQL1FPES2QcSi8Z24+ftiicYERBknd4JebdWjjrhkNncm1LnBhnwIcE3
GgS5PmMNngR/GpYUjO8mBOiXkefv19pRHEBx8uAXZFideOJ0LSaj3tdWnbrDv1DjeCCaCEAePqPe
XFMVUGuWpVLt0J4hA8vtagmyW7Nf2zyksyiAQeo1ip8mA97R6RUML15JAYCDjzk004R7zdwuD+4X
smrKm6e4b1VrnHbQOyQ2zuynyBHe3Q7PGaJ5kyeHJWdQZeUNGbw/ox44udPLlsPi6vOPRGtX68E2
VabZCqTS9NcjYGPwbo0DGgWK/9wcOqLtjJjORb2HLQclWfM3Hrc2ium3iE15tbLPObPIvZKCQpmx
/jbJ+XVCdCBv3BxkH2SuZLnqCU0/fIpN9pgzeyuRAId4nD0xjD9L0s3T6Gmlck3mOq467AZmfAaw
Ax/BvINaA/GPdwyj9LbJuNI8Z4xYVeoRARGeolOfHL5FCrOuZl1loRLo9f2wz1cHTCy43i1c6/77
48nqPStHb6ymkavE/NOJPVLFvXyU6zkSlJhM9Zrb9EsoYlonmQ9UzY16Nz+vGTcxxEuUS7oQXkBV
0SuzFjPiY0qIeh+FK2MMzFCG7zh8ogtcEeFhMQPB3dlJsdU2jc6iYbyvC1aE6bDQX9gw/ayHfcgq
7qVf0f0w18Vvf2UzLlKuGwh4lij9rAOCbJ8GhtYsf7tm266iQ9xqzW8ZM8Uv6rl0wmJB7Vd6QpoF
w0GLRnb80CN68Yk9ywk12MnS2pjAkxc7MVSwKXNghoHVnjyBmpBIAvEMoi/gzudrO3Q52YJiuR7b
9sBz7Dw5B7ECGe/5XSe/yjHPOFCjQUst36eiokABsexBYr/T2VBP4srUUY3wcFZHpGt6FkKdUdye
hSQ6409JOaJkFjrvhse/QEAs+vKP7T6tFVVlyttpaVfi0Taj3+zQMRU5VvSz1AEnZj3NuqymLQp1
yWMWDzWt7qMDo3kNSSeyrUqYsvX2IA1CiQiqCeBQAQDQyJDplPHclqIY1C0kj6DP3fnb7J+bEFXp
nygUxnYjtzMvf2DRHon+xlLMR1QbMeQSjbttaJDlnb3HCtt3IOj9peNPpbEH6hMmD0KQhME8pRlM
k84eMkc2tXKuwFXy5j2kMOkGDTuT6xq6a6N1LJ0oOuD/OR/e+CJLh7AxXqDnM+m/mYzyBNWp7J9i
AF55adFVVibo3t/CKGNh+qrGtydLg759q90EPh8DpFfZ6WBfrSKm6bSV2oP7HgnhUJ9kTP9KkF57
873ePuNikVrnxiamuQaxACG4c1XffEsRkIJI0oAvYHNTL0iToYdzriMWdhXBSPk1P+Gmu3nDxrP5
vRXP/pYQRPYwXHub2cPFHXTQMZaqkk27KLm3RyVACxaKEV/pU3AnBJAlU/PY8eYGpgPCm1tkBSPz
ZG1C/8Q3xGF5j8r3tyz3dIkyhG11iBoMkDSgko4RmsQk5YqQ/FT3sX0tv6y5IqY+TUDN7MYyYm1T
hx8aEu4ifQ61q7XE1CDKeZ/D/MA6DSYLqyfjVDPQVzYInyOtgEyorFl1710JIaV/dSdW+vIewzNp
wriSjy30KOygi+Uf7qUvH1PIk+twb55oCG5RUP2td7eNF2uANHF4N53RyQu6fabBuh0KSdoN+cuw
dXqPtVT7oEuBrn7LWcYKKYoZeU6DOh+eV5I5gTny1tASi21FHMYpFROIM/NrF1mwve1m6ygioAPx
UW9vpdwadGbZ8MpmTqIlRsISuybuQ487DNfIZCCRVi0e3ZUveN+9w7PFYRo68K6u1Rlew+0hhvyX
tkL9+oUhN7YrviugnzgHoG+iJngw8mX5tmlmjmXhdnFQT4G0GQNQ4p4mEJNHk6pNVt5C7K+ueO3o
0iEYU5ksoGbcIe4VJ6vvpknKMbT185wS0KhI51J+66C0svTV9GefN/5S+JoXVXeyqZaFRfX5k7kB
FNAHV1NgtuKZi0Ku5Ev+D7bN79XQ+Ilglz+/GcS1jD93ZLBcPqbhH7bI/tF3G7QPYMPy4CcBjo5d
yjq014Y8wo3OwBJtXC4axr8pD+KQU3dsDQx2BRRspsOLBekTzOrlcyKEB6awx1ijWT/j8hLmn7eW
Gfj5Fc3J/LTjlzcchUtBBQnMvn+iPqgC3lDYRkPoo8SmPwy0tZgu5DRN2TgO3hTICIVfSLvhRg4P
cebWr/sMvOhgBzadeOMfUASZiTmrnBQpDSvHXCRaIqI1wAxeEMV61S5Pfbf35hftrNnXHMT1Fz/O
YKqT5NuICBUDbZ61K15eBFFoPZT6mW51cid8t08uGKYlhNvsVOC3MRY4/2tX+CXah3Pa79g5b9gK
RpSvUzlkbpjKFfx2DzSYBZb2QFKmOunEqP6DVDxXEPPwZyEFsB2Md+gUuyb892kLBhmoKSaV0CvY
bb+AyddFdrH6kgr/J18PWz4W46RhQgCm/dwWhoE30u0ccsbmfZftvzGaU6SpCUbjw2IemBGG4svV
uS+EGkjob7fsY2LoL3lXMFHvsX3KwIdGqvfuaQlt+W+l0B33wOlczvxVe47KYV1vUymur6LBB+TQ
fx3pzgp/7AFcUProVzRq5IHQe+Lkr9Nv9799YTYKP1T8SUQCPFtrpY2C3XQk81fDwXrHF3ovvBXE
u1NKxKjebwSmQEOKRuf+mP1q+80BkYqkofgkZ7FBKc0x37euo7vkIsTtFlWLos+ySivxogc7sbkE
VHPy9zYJ4c1lqZ1q8ppU8P4EMQkbyaLiAXYYODx8pqIy2Ydwv+Zl3i18VVP4oEcDcVpTjVJTRjBU
WAIaDuWmqWCAkhdmuzYlNqiL+RDzc9uRMyFEahpAcyUTV9klWY0yKc8+d15bcnKvavjYSuurS8IX
bS2Jtof5n4wCVCJlBn6K82TuI5SLEFrHrsT2k5j/BXtzOT+qGZvDxWx4cozO3oIhkrJaA0hmHxwq
ig0ri8hXh5LRxE7E4bDFU1ZxfsfZImZtIUvBwpyy7T2bsUNqyQjZqdfYkN8GHeoSL5hq+8wsjF99
PRm9HORuH85tuv8vd4D4TgtwtLgl7AzC6hJ9Y4zJZTL0a+9vpc8zJ9nmg1Nvm24G8jmmYEPeaZ+u
YME1x6u4ljTTZWkBmZMSAyIGRJ47kCKHNP+vWXOTjjaiboX6TifpZyPdsnc9XdOEup80Rnen2khu
5kGxFT/QmABCoFV0NYhvYruB4lVXxYKoloFGst5EgiZUKhz9c59TX/tnlUCLifyKl7rrV6q49oox
zXVqD81cGmD6+N9mbxd+MPsYSmE/o2RLVsi3jtusx+ARfW9qJVQ5acJ5zrY2dPli1SEUj3qqfQfU
/a2wbrgdRTmE84v0IOoG3nOp/3j94Dm/Z9TbNmFJWTNHFsCt8dm4FYUjK2PbzbfOWhc7FZ88D9/h
5LURa69JcaBG1imxxqQGNEE9yIf3aGnUlMuJJcp2Gic2gLGc/tQLH30py4c71nkoOtpdJSi2NNMV
I8lem+OuL0SywO5ntrewaontfMdtrb2JdGLVjK61PJ2embCit5ZGX8YK5UXx7HWSdDbh6y1ygr39
izh9dDA6gTArW8rR4sqrYb5ptcXlq2RL2CfjNz+PR99feb+ql7s3NbmzIwhOTRu2C+l02nhYYh1K
BP71FXi1vCnau0EJrHbUusXIZZQr2lTau0yqp/65kahn4fEFkEbqc/Ao8LFgyO8muQzV8/npoaaY
D8P0x/ikPWAwshFfEK3LOPHGmC9lR6AcWYewNBcsLpnqDM0XcbKz1VghDJ7WF4RA91EjbdCk0o+L
iGI5+kAkqwbjjQ1CA19jHJg3Qe/9ctCovj2Te7ceyt+Y3TR6PDDKynLQ5EPCgo2FdNCcUdm7Xd+Q
xX/DdndCPtBEU3fb8agIcYmjhN4YN+PPCvCffCAF1al39WPMF6Tq+oPZRbvpHWwE73fnDr8mCdoo
yypAPInih0z02N24LSeoOjNaD2EnWqUIjB45nyZCG+Re3ugSgN77vJMaAHlIYO0NawQ+G7TUNMZL
+eEQ8yMWDWndqEe1uyxdel3LPs+WtLPwCAiZVGtqIzJMMC2hWTCTZYtdQ+TGHKsHcNCST6nnIFzp
89MT5MfVTNrv/L3HtsLzKr7tdJLz0eyvLrHCfGAWQ3wBQ5sU0hG+wwnV32ro+xEfdRHm3L5xQnlk
pMH1BnD0AQUR34UTgSIqyFUAAqedCDewrm6q1N4HP4GlhAscZklGubO4wBtInIK5RzWLvzJK13fY
XNEkzX+r1ZlUzi8PPNKzXPQBlyP6JrDdu65B9uphcju1J7+S4WFmJiU1qluSo2ttL22OlvmC5gmR
DP3pbxHXvlYyDsCatzM6RmrPZ4QBdqeI4C7ARKgQXUg/p9F3hl3QpoKfE+rZcaRA0gBrEfc9o8oR
E28ZATbrVFKxEE/OShvsVCyASdFNVbBkhaLLk9m/x/mZpNVqJKr+NmB2QyO+OP9pd2v5Q3rIbvk5
M7GmhNb+POwHIqA+714iqBh1LNBZW2BfHBiuYYJ5wna5//gozJtALTcVbxy3ZpLwKRa0WKp0Q3Xo
EesEe3s5z44RT9bd5FXCv6bR4bzfg8lN2inf1oS86sdzEpoALFJ1A757Ata0ApSjfKJjxMb/xuSh
O8bWvYA1Bce5AnMXYEm2ggpWdfeqXoNCON9KPRTzBD0b2jkrMTiOXqaCqhRL9sO0oqTPfEyD/hjj
yz0Y2C40xt8cop0dwCmCglWXws5Exf6O1it7w7HQ9qxlrox5oyoEt91V3PJOfUDl0FltpmdMOU+i
nJA3W6TPpAOQni1FvZXEydd+QqY9SspHhGUgE+9lPOxQG43z5IPGxWovwoNGYnZLccs2KpAfCPG6
Pv43FNu87HmfYv/MtlC9aNEZsoQf2TrSOpJLozThOCwoQFCSMBGk/8OezeMpdRU+VkiJe4BHy/Xy
OsReyXrn25ZVbF62sPyjB/R19VVvZej4DPi+M3K3X3zXsYh3fTg+YyWjQC6HcJDTSxQHpa/saVkf
Ns+kVuGny9Mqvr21FpNwegy9sa+7RU1Z+HmusizIwMHBIJBZ8mgBPNYPlchkf74ZQ1d/bvuRqWyn
0IVQ3UpWpPMYyQhCMb2A+FSiZE6urQ+46OJ8gXWMmvXPzTL1djZ33B+eLTy/VIrNP81pDU/y0aRV
XXiwbuc5Dp4rbcv6eRGklimBkFsEfapYxFEqD/l+qczL1DcUg9kR9u1wpvZsPfGUhyeP6Ngu+Ykt
EtVz4gfg0Z8Lcm+VqsnvW3d/mOk3qvmhGbCkQ/8fCogWoiIDpYkfxlV7hGqVqwBBJeo8yJquXQKl
TUUG87gwnn3chw1IWsNqHWhj5U3Bh7Z0Y+D3MRCQbghPg73LRxWXfBAW5XHlkB0Vy8yVAeLg/GAd
b3qTlAz5FU3vIqHPtEPYfLyGZQQACBV4cFKPI+3NxPprxBjVQ6zE2083zk2quH0w4W0T0Ee7puQB
qT1jf8HSbkcekL/GGQZngC7EyUTWPLBvdrF5FTkq1IsoN7nziJccXh2x132fpBiN94JK8CuzJhvI
NbBqxDZML/kymY/x5GUTMCLtlVpnR0Qymg/p0wyOseihYM1EhMgvzcWgTI73CLCPqjR63MunkDK2
mpTrOLsIzaMwgQAtGkmRuI1d2mwmkhan1QXM2+MbHfXZxK4kpwPzdPiJatxk9EqyM8GbHgtccH/5
QXqyjmmLANw6h00N2r6lk7PP7m6FT/DmQXK/LXQwTcD+ea7Lhowv3CvfwoDLmpTEx/TLuxVlnPrK
cem2GcOoJMlqmJpe29SUIe3CbJneXy6xnLCRuFvf0zq35+6NqGd75FG1rD9U56ETGzfkQMmrY/Db
I3LgagISmL9y27iyHXN0J/2/JrENrzhdgzogQMMkZ/ImQ+E8hFKgdulundvjFVWe6WKjYy+pq1rs
rqOtWQrafHYpOBumb/OHj0OwM/o9/fBvZB3hC92HCo4XBsnlx7+z2/DqR5Gs95VxEPU1B9Uil0e3
PzTafb2WL2CAkRhq8M1MZWw95MX8NEnO0IIcODr/urkffkB0hZlptSY6Bfpc85yirsYKc2uq9V4o
HHSDor1zpgFPFJC+tVoH27ZEO3OxMEWqEkp1IGpfJBS1p53hV8M4mjyz3cZe3/h/IiOgTdKGekk+
vW3PSSTC8VKSXqcvy99rgCksOgt1c1Yccpbz2FQpIWkGMkZ/MmuI1I21A3LPhjQNte482CYowmw0
ZSk6owHZ0YnMFnVqNZuoBxPBGicTKS52gg2qSfLfiNTHCqfoECCUC6WneKcU8prrXZgDgwqfSsmw
SCeEUDQMUovJy/Owy7Ar54GHNwpTxbaQ7OgjDWfCk+skW1ydCFoA528OcvQOXPEBEfgl7KR9M1r3
YODsa5xk9PhzL6mFy9xcNe+yMS+jAw4T9BWGYFguXiUsOrhl5qy4Zc4gMuu+wmf67zlRDqbkDk93
355BM7PH3MWwDZTxoI7aB7mGvUMlSVhYP+sevMk0Xk8nb5rESojl1HtkaYbGOiS7TB0liLg6m9L9
USV6cvJcdAkP9l8OHgNInGaGl4/XJP4REyX+VwobD23xOwF3dEQCM11NsR1cFDqlm9XwUBtbkILc
KDKuXwfC7BYqRkQ9+qNSTlOL8fbT2mkhHUduocjwgGUrPIbjOnXY+nPBnLVh31nnOS9W7MpVgkPj
9dJYkSsgzsiNpPigQzCfSHnW98MgxMrEQ5X3KmTf2MVErNhQCP3ct/tNH6LtXTTh5OW7yyL4D6ud
TZhOLsa2XG+KBepBKmDA/o3ILRgPT0VkwRNHKco9iDIIx6dpEC8dvbq1wngsQ0F3Hl7MeWN6rd9k
+P9xpuei2YvU7AWsczu/6qyJoaHlv9n4EVUV9cFj8TYuE87O2gts9P9Q+xeCdX8wFPh+3XMWi9pU
xNs2HUXCvCO9vfNckF5w5Fo63LtnWfZvaRRot4LepkZHg3w6DNcFbwsfOXpcCqCh0zseIe0ug2g/
mdpyjpDYGURjdja10YvdhbzhIX6dsThT0RpQZK4CBWE2yvSyl+IQLRE/lxkO/GU3XhQ/VPcBPzCg
I/HVMyUjAq5f9wPXwfSbbkFVQGKSmGw8I9D7Q3vGHIXik0V/QjJA4UTnJxATyYSeRuDpWE2Mo0te
HbqklkLmbAXg2U/Qrtv4pVcdp3Qh/erDvccwNpwj1i8pE+3vIS3JGROmgxtdtHZrUyZiRXIGoU/+
5WVlB0mHwl4Wqks2xX410q43U3C5h3K6RUj1vD/8794jK7lHxc2PIED13FPjMGsmLZdX7gLDnSLS
hkgR1nySgaha4b4bJkSUBfbKWZ8C4zq4I6vhSTK3teMYe9+aZfrMU+Grm2A8VUt1is0uKPRjiy5d
+0cWFUg3KX9tnETZxI+4g9n3c+ghD/Q/nNTIrEdiGmXM5b9/ozlcfO0a8yzZ2X7UKVQh9W0vwsAT
sfrbyu3J4CL7+HysbCS9zl25bsDdm2onVgPy+Lzv6kYLCmTvBVRwdSEj6SlrNLrS6LhcdmRQ7kJQ
Qe39Rk+hOloBNZuzBft8eUemmnbnunUXIdsgo8JJ3jhVlvUKVucjaqKhqHGvJmpw0y8LsqX9nNqh
xtUaByA9h0U3xvETXoQvD0VD/p8OCgjk1HqGGmiV84Oq9XLDfiP12BcMbmdl9BliPyMrsBzF6E41
jjmUDDDN/pQL7dRZVLe8XIDryUdNZdDCFB9vjXeAZkaVKFM/p1+ibZTafC6CBA9q5/fQVDN3yosz
NIP4mxSASO58WOE+yFANQkHdTzGZqoOs69Dj2yh2cv6Q3Ix1ke7JOuosbIkQ2XjSsFBtfuwbWqC9
TzDlxwOxIKA2SVUX5h7u5Ap2xlddKfe2tFgSgDi0LIVQ/K0KFh2LfU60rc48KlVylI/1GVep7Dkv
CNzIyjcQiNgJzCjFcAmxawnPATCNLnZM20Sa4fExmhjjHI8HQGrBIeQMme60HlHLm/3NSgWZ5f9H
VJk8Zyl1AVziB6/v+KSKAmumj2q5WrGvOCRuzHw8kZyOxXQ7BDyOWzAjuNhjgRRidVFsB/gJLi/S
+Ik7Zc5G6ayryE+48KozIFaI7Sqa81lLDNlo6/TS+6jkQOzyzd432SXAv8aaxZFS2CGHI3174+WX
8L1pXf2mMChk2xB3rnJ0NVLBdzkb053FAwxP+IiNUbNM4iIlhB3mCDAuAatB+K4C70rlOGuHVvHF
/o0PN3ubnPbE9IekbImGgijfq0DYe7KTrTCtvCdHv9Wy+K4ObQcLA0l2oLkCgTAZ2bSqcqSlgUyw
xmxHaa9kI7B2kyTzKcOYr2Ff+42Hn91cGpnIqNNwVyjro3uOEQ+oLmYYuNVTvcfNgqAL7VgLqIbK
PhOJ6BjWzMrsbVTODMR4Mi/gikFwAv1RGhtiS6hB53HtEQfDC52wYgs3Jd+Ij2oDHf6YtfAvcqOI
aDtN+VAg7W9Hs0RTN/OPyA7T3VzTvlOJ1qY62+yCqorEijGOqgqLfJpLcTqQxLGF80oDHTMdZ3ur
Z2zeDXASQMs200AkDEaH7xeY0LSJSnrI1TaIK1oH+eka41MoLroAJDeThXb/LUM1vGGbAJJYxqkf
Bp26ze3I1fYvSlzbUivlelnrWn/aaHTqqsKUSgYTvXhWJan4YuG/Zje5yYtrZzbJRhsDeWyjh/tJ
KhgoxXLrIqp9EiXzCXlab9LqjL7YFFcX4DLAfcIuSnBB9oftbENnOkPT0+4CxLuMjjtjItBmpsjh
1iVKfWPpu98zuJtenccwBvlpSi3PKDPeC53595DT32PgvIesvtmgYp+f3ImmvzW3i6MaKQ1QGie/
cMC1x3SBiO7Kl0lzQSFYSDslImj9BK7EeIZBs5ChWF03LoYplQVmdxfRNdoPkwQe4zn9y1VrgoIS
nD3kbE4LJd7ntUyE/S9LwfsF0OGgT47PBkcEDPo6eSG8q0MkNct9HXsiH8Y32QGsFsFpm/7dlH0b
IODzdCudq3UTKUq9HjjWmSVNhb0EcVuXKukx+rhByw8y4AuAh3gMv4cszg5rhWHBaiMO8kRi0MxA
xo6GEDBRTGUAw9k0H3afOFClPbrZv2vF3eTyOnEP59HjRulDIt08n4AHAIJ2LcNQJ7oc2OWDUHVz
wT/W7FxNRoCB5CGS6pIvmvM3qMnfxotVh5Epky9onscdX6bQpKDMy5yaDyNVizI1+QGUN3IMut1k
8m++6FuVJPswG7wo5LquWWZhfnNTAyaNcjgpzaIXSVA/o3QZfqOsnwnAwpqvnt/3BQflZrKH6n3X
kwtpKN1Lq5qzLJmwjXvWAgr1BlLk0WWzpmwE3cfQmPm0DnUBBBoH2BeE9WB3qaFWa9WRuI5mOh2d
1N9VuHTvH4XRkouEnGU6Ccj8VbS/ecQhMChy7g4iG0buBNalnR3tmsUWasiggaK+9Fi+JZDabnb6
TlIcWClAmHQOTNJYDsJboNuBRJyW8cMRxwQ6POY5Tyw+i5WRkvbsAH15FWRwQQfna6wlCUQ3ZW6W
FNs+YH3Aa4DezHxYcw9R7x2ePttTHe2pi+4XH+uQXpGbASC31CZ738VD7hNWt7+Ol++Uc4yOwkod
IgCXrBGu5sT6sdXfKCeBn17/LbKmtxNU4Z9F4qKhaAhAbGCF8b1ceESbQg37C4KmmSTLkYg1V7ys
8SsBx+M+I5BiVp4O/3kaHGGyzLix+po34fh7+Sv5p7kPVhbCrwIGYdCUytcVjwFvHhg8rfqZS/eM
UCWl4rgfTbmv5usJQK0sv0lA8DcUP1zMkgrLakG0uiR/cxBncW8pkkRPIuCZw7u6flYzYom1YrT+
SzskOhVz+WSjYvrT/ORoB03eDwK1C8j324KqWhB/LtcyBq+4Gb/hJ/1UdMjqB0i6S9jSozp6rWbc
rs4OKGlM7GwMG7RBB3+qZEIN00vWBuMnbsK9UlT9uED16d4fQqQno4zQWsPnhLRPgnCZLRl6zKRL
x9syXKWQ6h7xa3DukBuPvqXYJgfi80GtXvaNuydKlc5BmrWF89x/p9kLxnCHn8MVvcNGed1o3m+c
XlVBhjCFVC5OvLxr7noVDaFn/aAXeXh/Ysp8mD8WAurFtgpcqwbmdC16S+k2JUe0JFkp7aKGdpax
w+VH9gEoWRw/mosc+JEn0BP7U7hOK4CZ6mCyEy/We+6b4nNs6su69Q2cEwSqAmn6b/cMJBe7z/mf
gsqKEDVMC3eQ8MqKvfxqjssVP4iSEKTnmJ6+ymKUJHl5chz87FUDtcvhGVDBEjSJS9QlE0ePtn2/
pPVWCZyBdarXScBFVNTPDhmrBJF8PlfE9my00m7ZKWJfs8lSCBdou9UWk1He2jDSRCRagxlNFShP
J5/89U7NaaRVil5nLVLEHfZ0NPZQN9t6Sv6LIOKmn22HKsDQJ1jEmO2U43M82qjJcaLSLap6F0zM
ztdi+9312m+XB5pq49XkYv0ps8AT6Xt+DGM5hhVfO9kGSvujy+Snqse71I0HdtDy/TAThl3BW9fi
q8MLiaRJjxYjBMhHbU4kydWKa2COMPzX34cyoGCqj9wU4PcBIJ3uYxWdbE/cOpGDmUrB2Nu9ndXl
QTFcikK75XFRi6lShusP4NoWexP6pOs3z/uXAclMJVOnmTVd1S8BEngICvyw3ZSt6KBWnz3Db6fd
fmPpmMQjMyvedNxB7BHg/u39qVo2eKP4l2ssT6ISEYG9LJ+bhESpUhD/Kb7gqo1iSHMKOluAE8Sx
jD5Kxws7hqLJ2DfYhsksHfHx8X3kCCiE4YoaoexUc7P8JpalbrV6bCgjvbEKzVGBCmKOogaprzoK
nQ7otUKTJoX4Q1QIt2rtdgOjXOdTxOl/6AH9Wawz7KH2P7DsIczWJuhHW7WitcYLRgKCer8uClqC
VEQ6jGp3vVlHkr1eIFGRVaT27CSUyRPnI9m56NpItXwWsRfh/Wtz/nridcGf8V697OXmecNEDC5E
v7XWtc4wylrvaK1M7wDBfb+WfL2pGpRfqRGd6rPLZ2HU/qkpTtvijE3UsrMRCLUrIKlLco6jQR5e
e/3eHRJKpR6mQOugaLxdc11GhgTldehm34WshI2DKwS6E3j8eGq5V+ODhcfC112vXPn/OfHigZFE
hn9em2i+yTologTgunNN3tpVqdXaT0uHT9AnCW+Z5YlhNoIr1vVXyD0rvoKIJDxW5rWSRFjxovTs
yZfnBQRSuWdXmU0Lcdkp038IbOU9I2xVZqiLMxfGtCWzhoNrrm3WXuNnlgOdSO45ZODl9XSA6AcZ
Wuda8tEVK9UrM8W3Ge2rriomNmiRI972+rXzTssDU+CY+5HwPMAm/c3t4RGmIluRZy/96xPKIIQ2
NSybqodGfSxs++8hH7JPYq9exHV3S65C2d8XnM2upPG0+VxWGqOon+kC1NFPD/4O3Wq44IIB8MMf
U+8/HpruLBa6AvS9tDhGs3af24YfHbZ4DTYL3abuGP+BPeFhQXaHTDVbbhgN9m5sOSOPykwQyoMT
DB+pQjIFSIzdqYIN+JvfbfFj1xZ3S7xSGTbjc6UO32ziuWhxQAofKDoOy3q7L8FyhYWO0JhNrEtG
aqPN7GpCb6qAUMIhsBd9YWAwUG/KygNkcvVPV4VfSC+/vus8y7lZzOy2gyeVHW8hgqqqFmo1aBIK
nX1Nc7NX/jZiVF/hPm+t0uzBLdyWdbC2ewr2XqWe+Gsqgb+sHuvthD4KJZOYxWJaoqNtvGvetfCI
CpghmR+l7QDr3Shkx+iSMPRQxnEXu43q+6ofnBbhwE/padp1abs5rdPeUbWl5YmxtIFHZAjXnH6u
kHYllILKVXbidh6vD2GmhHzlZtURbRZRpGATiFmDAHGUAHMvcq9FFBskHoEmxtsRCGNi5rhTimiz
XDDr6D+pZEnm0U0kxRWSyDc2PI3y7rbq++TUFycaHe26kAxd7oIMbtdneI97QQf9Qdp4lxEa/WF3
+6hL6+6DZGCNqxUxYICvEjSn/eEoCviUWuyAQ38oCfclbC0FqV93mMz5YW8eeUxKstHhoSARrARm
5ijeRjZukJx9xHPSXW7/E/nvkqqbkGMAMyAhw6Nanq8n7OMw1eMcFqj2r8B7cxsnL6aE4h982o74
Put51GT46XG7tEI+2iILasSIrcskXQIti+M3T2SzZIZdCTL+TMoupR6BgcN3JEAB1mP+2PWiezRq
vqFO9Lm8W0JEYHDfTHLJUKJa0LFyz4kYVm/mtwA93pHysZRqN6cq6jgzKleNCa5tvwE9KxWl7MU3
J7e9G16tXKIhYJVCF8TZnQG/0Tl3XUrJ3XHGSrXmMNeSg9cBYRH7kiOnJ4eA+DyaaypaNJkhw2gv
CamHLe7NhYX6nNgN21lYHesWV60JmhUkcMaOduIpWlRBJUXkXuR1pebJmh7gdCNyfxigp47zs/g5
K9W9pFXGQzChLTQSfnePK3gW70j8F6FQNvYmFzrAgz0Bi4DOEZNvxHgIFllMCwpcvl6NG9gmD+r2
5OBIlIgmfpn0O2isSgE3kwS1G0MucASSXVxL/yo5ctZyMDyWoD88UPVUl/8X4YnuMGl+qJZQDSUd
Pvq3p9cruEsqT7mjHSlMt6V7FsDxqiuERPezs+PGuj+QOlam2S8eqr9OXdXnFGKuM+p6z0A5DsfC
+2g1GeacW7deJ/Ik86iDsK8p/FQ3X0e1aqTyLO9xX2nzBkH4HFPBUfbc4v1DMdPqS6LlEL6jraRv
0Lop8SO6sfNqf3Gmhkh6d3Ti9qpVoCrSsElTIA2oUQHVUlj82y5eqWqn33svTZFyGrAiaBmzwhk1
Gx6Q0GlK9ETU91ePhfVCzZO4+vlbAdZRbSI+4DogA1FfAI46oQZisgo0NYoKbN8Lkr9APfuS9KiL
x+yZ2Sh+V+GagRedx2Wsxu2Eprth6w+DNh+DwnsboBKvSJ2ScSBFWxgapa7SAiGr5HS27vfg0hUp
G7EARzwtSOAFXXRv4OPybcpws+52tVcBI8YHV2tVQVzkyag7pwLuXasOUq0QuKnpZPuht1iTK3hJ
doS2k1wahQJ6zeMtCUJiQIIyop/tYNSbrYrqZu8KQZksRxDVvG9DG6QxIN6o2k4/bAKdg8ccy1Z2
2hjMiH9sDjGsVOLZQdzCf5UsEQy4oCdm83mJFP/wbWrY/JspL3aX7T2J9NoNdwM50hXGugV6BVwk
pQr2d9ufOzHJAgeBZjH9z5Eg8qoS1hKbriZ10Vcs1eepEkVX1CKj9lj7Ynifgj+7GD2MyAs59fZh
O+JH8wRMVGnGCKZvprwiPGkjyYMBfduIz4YNfZUlAjgEMZ9GQ8Aslei3C5xXZDFJtNCCq07bB2uY
VX4nntSL8mYy/KDLeEgonZqjMJZ8bHG5OAC3aeowXNUsJA/Nq7zjWqqyhLZe09N/dRCk/4of0RW1
+D2QnUL1OWaMzlx5otIc9344V4OIZa5fkSFWMpNQk49delAGfZebC4OeogWIIF8Ze/zhpJsCRFCr
p6uPfZMSpn/+bs5vYfUH/u/KskuB5IoFPezt3hyjrG//sKWfDjCGAGXqhCtPFe6hxCEzYDPFLh6K
jWEmdOeDVRWQ7U9o3HWYM4lPBkujkey9LPZngE3tkwFR4sR//+wihwpQmncFh5mgBmmrzN+PTg4a
ilDBnpOl1l8T4+n714Da7V2JaQeVqAJvZ2fkX/dKsF+EMR8vGMPhOjqkWS/7SFKho21a7E6RVW6B
bNYNF/SfhPmvYSbbHI/s7VziYDdEOisrsSqkpqwNKRNC4KfHf5JOAya/e4BGwBzO7qMnfWD7D8Pk
Fut4hhNGkME45l9ZPSqDrNBlJ6NI/u0W9gRj/x5pl3F+9BZw0I+CWmwg2RornncRc3qHeYB8wOUD
m0AQLlPfQKytmXtUlqqB19zlJEikjls2Ro4gPT39gSAEdJiIp//gK1iBV65Cd6xOpQAGOaJ03HHu
rGWuKkgMQ9d8HsntULtfLwkVY+NBi7JIaI+3qRKAQbrgPBz4dx6Qtvl3aBm3WKVc7swF8myD69j+
2xc2QeYqGYJDlGTk0uV+eFj7aYC5mkgjm4kYTxs0MkxIjr/70DhY12Ubx8dlZi75Uy+Pn9nD2FGy
f54p7OK94/iR+FCkPANYCVDeExPsE2GbBkMDWy0ETQweaO8I/PSlg6lRDCdaDbL5DxIoPLrk1n6M
BLT/EQTUBt2WJ+hOe9RUVFmLTpgCeIk4vkFer4AXW3mLY1c3FW0F1F0KD/afILkLH2ke9syZaRdE
T39Hvxq/aABFNzadYIwRaaZboy49CfwPC8jK+XDzfleVp3RRhUxvRaiyK9TkZXnKEunqQr56bHMt
yxgX4EGOmSDEB0dOL5ic9dN91kMDI8tGocEjEcmA0iACT5ThcX93KjWixYEenym/MGPH5EPyqHfW
IHZsIeyaRncgYliDuxR/bDWa2H8JGbC/uW2V0IVWEd8p/K7wpj/XbiCfMAXjgNzjmeAGzYKEEcq0
F3coc+vEgHyY740oWHNBVVKpUokr/GIaTzbnxpHLdmMw/T2Cs2sPssJ+tM0qQ0gyATiac4AUGqiy
ryeJ/ArrRr52EhiaXQW4sOA8/M9y4nlh66A15oK25Cqt5y9egI8Sg/Y3eK8jpBboiTYtbfM7GUvN
5GjqGGeglMDmN3QZ6fElYN/0jpkUmC1TzpFNdjwdHsFs+vMwiKWJSfMLUha2QUOhtq67xs4ZECsk
OTIhsbejCIXTW8oE9Q+x7tcoOdgaNgz9+0mP3nvruZafGc9Zf6PSoF9rWVjkZ26bydFA+OeEiV77
Jx6YhmHdpiVoo3SeMCUhd2DPJLrlh7Yw844NhHK3FMSU4MPgs9v/BzpIy+g6Eaqkfijls+hqnk/K
MVEr1KTFNjKQCdmmpMWnsjGoLXG4IsqX4HooR1eldk71XnhkJ9DFq2RXqkF9XEmHvjPuBfReCPCw
jRa7fWjJBQAchDLB+fEuLaOpOICltac3a8GGvw0VgFBU1mVDyDClkTsz9FhlJBEFzJ9nE1OTao0T
hm/rtwTDgZ62dFA1BKJoWKtC+U8wKY75uBXp5AYYEla37cNqRPbYRazrZBlh0XXCcETa2yBtmj4R
UMKfIFnYyLgiY9dFfFdw64LxDTclqdqvCzvFFhomSm4UOeUQto9LLZor++GFSAwMfJx2/F0T35qC
+Pj6UcO38zFd2lmw3nhAsRrA1wTOyrm25zbHHorbEnezU1J0f3/qimCQzlPi1eR0QqcUh4O+uiZO
rDdqRVAdg8IhxrqD50tr0jJ0gR75zqV9m5fXZEug2qNw04wHWzXApIhkOruuD3jITWZkILQASnZy
f/ORXSCPfL84TfX/z5sVy/60ZEnpXUgiSTj8Rz6w7FB7hMBDCPcoWq+MXicwQHK1CgvjvPopo5OL
8+30KgoLU3k05B5EVO9/+5P5qOd5YXuPDuOOA1c18+DyY+QttwbhKXTt5fm6UNrwcB1enUiqyVoe
VHTHPH6Jr9/sIQxfH6zMDIXxhCagQdUm4oLH8Ll8McT1wbWLn99YOb/U/5u7Hl5wXHHm27DMWRTn
wVMYbqV3BBYaKmnnVK1WO1Md5NwgnmeQWzyjAIzXXiiIP71spwHV4xzRDl1IvOtavBZE0M0GN146
6jGW/rPdDiPMKsmBRTJdnz3xyaWrWT7fcXL3hbP8D3PQ+whEE9ze7MQXdcgeTP5Qj6Di43Se+S9m
bAduQl2w2gwgZAs4HoDk/bM32H0rGOlo+TgrlknVRYsq7OLDhQ65u/rDd9+XWu5lfEZe3IugLeNC
h9QkZwvnspU04z1k3x/MkUgFCUJ5SB6Sl7PofPxQSEJQs9pQemmZrXMgD8lB+d2pwcX4jnd3pXYm
qiaO0s5O+XIQ6KqDgvxWKbiaMCBp7SrlOXKZBjgBNeXdrtAixyO5pkTt4p7UrXrs1KPxJ4Rrj0on
vmxl+dZwyNF6vSfk+lnPwXlEfeHYHJ8VgKJuogCxfZ8cYQH42dX+gqNPRJTaWOMYDaBthCf59UGg
vFU51RLWCZ1b4lVdLoKV8at0DfDdcnQGwkR2WsfXBjoBo5SbG5yR0jaVLHeDI8GVQZ/Dc+rRRKhB
h1jNH+1rj9rn12iCiNexiDyo6UoiObU79yZ3tcGjmAR+D2XhX1u+DC0QLBL1mhd3a+injmq3mMU3
anyoWZEYl+lsGfjUe0TiDk9xwbhojfZgH+pn1UunJDeT9WhRZGlyFSX7/zcQgF/Y+8Cjp/Erkw72
9rLZueCewg54JELsYuCrLQfvIQiJQ8wEpCvmDOvFdLVhAPeZOd0HQrTOoXXSkHO83FdcfBBmoRxc
hJIeUxCo66w/coBmdk7mO1e1ceRw763oIWNX81L0N6Q1oXUV/3buOGmEVY4sNihR/Mb+t7/b5K1A
5fkv4uoSlW+uUhSJ58x/vb2cUsJXSfaRymxAyfFU+pJTn+DetdcIzyWRBBxQQSF9Q10dOwhq2ior
uR9gy6cfthppJzCKHubHfHVi431Pg09JznVkzupSUI0mrOKQ0AavLRY/gkUnuJ9xl5gFUZyhzI+H
NXr6e2SdBNohJEa21j5Re8g5JDe80cEDx49xT95vdgVO8uPkortWt3XgS8jWimJogWYHvGss1KPg
xlNQ+K/d44z/Fq30vTM+eHymjWgqcGNPx2q9aThgi6pTIe5IkDmqIu6L404kRn4C5drn9mr51EHr
K/GSAzoQStv3JoLPuGD6JxgQKaisE8s39XyBDl1CDd+5pcIHNEE1nV4VFDo7mrUJBGZ7RRUuA+MC
Jw4RDpnS8MmoGoFC//XI6W1rgpUh5CqhAp01HdENh3sTbu9Ua5UizXZh7I1GeYDkIxbwbdLjiyxw
kdbCuoIaw7WL+qVv50KsZdsht3nS0GTl06PKy4963HSiNNSz2rAZJhT2xfQptD9W3AdOW+H9ymzX
EqGe2UUmY7q6gHyaM/K/ScocEkayHUTzo29hj4IfHCD4u7t/+tkyvjTowovVx16NurNOTHeMseeG
L9PR4CrQ78252IXEQ4XZ43xVEtxXoHhgaJxTU3JUKfjSuzitMB8TzAKTiJcsV5fPXJpNdGkjc3FN
/MhejyYBLmLiYfSPFOla2fa2P7/qULbVAkvH+WU4WtNvPvfapOkVVtVt9mQXPH+A7uIoPRxxD18Z
2e4swRuN4Id9jD4SxBmi6N9d8i1XpLv2UsWIfZRXvCp3PmKdmO5UnpZ5zNI0DncJmi0E2sjOy7cR
OA46fItytkAnU1Z2+CJf4EKi+ZN8tyiw1EoWno4n27h7hKvqtXeo3xO+Zyso9OjcO1+0HDanr1ii
mJVRjzfF5qJFw+p7m81oNRO8C4oLPQRh2UyZ41WAT4M4M8Lgntl9YuwvP+H8h0jPdYcgdPIZGH8d
BLwn30yuCnRbdZGsl8tenGKIOzc3WuJn6ntC3dsP01irE63xK8Ogv42yCCuaQsSFaT/N0amaDqza
cPjkbFodpoieTrJ/9xZjqABM++QexjhNrNowhLTGUeN+PXwW+xI9WU7Vala9X4ILaQfaG+x4n9Ly
SOSHL+M5OZ9Vh6H5WUtzaaHxC1FEtzN+aoeiNzs1tqyLFYk6mOux4GmQHTGkzGcTEv6JeJ1Ct7f2
3rtEHOV+ptjdIOyJz41UXiNITxATIQ5QAkbBETXEThtxsbrFzHcYFZiDoKfutmEg1JGd8c3dVUM8
FHpS12xDvlfV96SQbmtBSKMtxj2by8PHZC2cx0vJjIyiY2mpos5ZVRwo2csc9ESvVG+2d77MUkHg
f4/MhmsJwiP+NWfZngJBZuyyi1rei4W5UKu9RMI76RiHt/iJaPDTIKBCbznjiim3E345INfV9fyT
NdTg+IoIKGLkoM/q7kikMm7dFoCMi+dVmtvii4afc6QFuwKktcxY0/tHbbfog4qs6cHN4MuSQX5W
OQnrzmDtpecwSK4S/6QQBSHsYOLpTKdZpwFuhn1LNole0DqTwiOvZYLn0sjSxiDtug/yuZWmEbWI
eEyCoynFn3GuTZWkewvSaN2mdYNVuN3fihwh92vfWN4FVzwZlOBuPKdY/EeauzDNPvSj9KiM7VPQ
RQK2ECFktFjpWyzUmhwD1tibWzlCofvJQ+A7X4iBBfW4qhIU14GWAKa62OgcSieyQJ7mXABWkaGF
pkhEzlcbEp7Mt3tme6o0ONsg+TK2TB1OLxWo53REXVhBWmnbObyipSuVpdree9R2Tky+W9V4X43i
540vsOI30EBwQKdAqts6qwPTIQSAj8eZSYA1YcXdOFxrI6Y/0UaIt9bY5/w+YE+2hJ13BZ3yLpN/
gksMoX3E9lObpD25RFDN6QPaIOw9WNupetneWndUkXimW0A5wgwSmOeC9x0a0xwUPQUr+Su61WTB
c6e+/HFyVTNegXKFI6E6zSmIg/DMlIGUGT5gQ53iSWqcaVb0EQbrK4m7EoA9dpIQhf0pux/xHHmb
kM7vtydobxq8KwfUC4K4f/J4nIlw1KCYKJFYvobSUnOPQkdOazL9LiUCT0f2MLSvhApaiDR8g9cI
a51JV487I5bt0KtLzHjCddp9huZshwFcXM41aQq2xB5Ft63WUq0jYSa6XjgRBnPlzdA+Uh2oJWxV
UIZp5rxDlF5dkBiKTRrdSWxedkUToeSHHfUGe5raIMPkm/CeeVfqQUYGwUSy72VjOHQqUe3dUZp3
J8AVfj+JQZPvhs8IustEt/7FTnxiL+4lO6z3GzoaaNIdjSt9su8ytOCviyNr71W2C4D56hL6kwYF
QR1DkqoST2IyEZPs9aZ1q3EFWrpOWQqUgRmZEgD9tLFWPQ7B33vUOZLD8kwuAQLqvQ/HvKcLS165
zHJmV7GDHzqq09gGeBvpHyys3TAoGRcUa9shtbaIT8c6s08Zw+YiJAgIasdoSGjSxG+m4w2QPlc0
+AqZWhAGLl6/C1sLYSqbmAa5HnpazbW5rt/w46lYy5qPyofooMzw4QKKzN6MGGRqYQT+JvbICmnR
xfakEUDDrmWLZhqaPQinsjhWXF1NdrtXkIiPD66rkoG2gvn2761arI2+DYC9010SWj0oU0253wuX
v4ZSB+9c5yPO5g0KRpyforu/aCIZOlNWZuIQDumer6rmCJml/+xRHvsGRrv1NQej3ZiDQeXolICL
JMVbVTyukcV/YnoVxnIH7HnQxOp6w0Nl2SEVLmAC1dc9gX88JsSZGfrA/DgXqOsKgrcEpn2XrBFD
4ueatqhdtb1ISwaMgJUQjD2m+GrnNrmf8uk4/5MdDJK+Fs/f32FcFd9sLVOGR3ADyb6uCB10ZM6a
tseiMq0qabkTdS9hsBCy8jhXo2LJjZRnnObZ6gA/cZbL3W+CB9iapBS62Ru70mDlMLWjnUAqjHKL
2mrpbK9gOtHY1XRzCmpsUs8TFXNZUdOc8bOVJ0voRnAn4RB+Hm+J9TeyETTwJV+AM6H8c7hlXU8j
YO9xe/PgNpkuF+bsVHeKGYkU+fExQWrNMNGEWeHuGOcNcP96jAne2AoNXJNIUz9pw4oT3IQkoV4z
pQMp3m99mCsyucFsBTEc56WLkvkEfpSOumlh7F9CcKlZfYoQj6ssmg5lZ2tQqomm12yao30L8U0T
9piyaMgeuix4lfoTjH5Gmv1zux+GPScXrFF7qkeVCThjWtE4tmXob+Y9dNEFjEcx96Nx8YGLb9wo
7DQHOD59xYJxaguDCBSf/OMJ7MfvxOFuCUpcLNl5Bkh8OhwhX1r2FhV1pJYXwYNfMoDEOc2cnzKF
LdCggWFw/MoCtXhwJ4XH5RjkwdGrSVJS7vrz6FxtDWnWV/JOTvo2DA2Lvf1p+oNI58LElbjs90HQ
EfaI8bst7Def9fTshel6z1aevtVWJmOcBRkGLxF8ufW7zLGgDHIyZATkxrYns/bepYe8OITPcN/2
ab/gbHMbZzr7MEI1AFb2w2m4sNX9za9Niy9n238176CQGAOhNeVVJ52L7yLSTwNFgWpLyM6lWwRH
pvFP2bflELTqCsp8Y4p2PgbfbJRqQzbpQY1eAHPEpLkCIxqNxrhldd94P5CjoZmKAA2HJh5Ibis6
NtpUk7/Gia+t472gKjHNIasdmHWvKbeYtzorCsxGOJHuj/7PV5p+DXf0ijcU8BFUCvvz8OkDM1JW
pn5I+ac6iEP8M0HJTyWQ37tSEiFJ8s1cDzEMo6giIpbJtGFzVGqGRfAPl4i3/H81Aal/1Q/64dsv
IQfwODFLPuIXt037SK3/5SHbGGjFk8TIOyUNf7oBS6wQExwb2ZqjfHR9Ey3ZaU7o2nE84nM5/1mU
4fYeuYV5DTbgvrw5GAKUBxw1QfPMXLvSc+695rv4GZthXK1sheuhMk6EJLq4NSZKkYS15SQJ+IJD
iaslKU9jF0hBQT/acec0fszfaVFz+a9pzCQcc4Jq37d8M0fSX2KkvlF0XzlA5NtPfr26UIJaB5XD
22l/TvdM+nJoAut3FmEkKp8uCmZ5DolxpeiP/yglezhlT+Dt7KRSIz9iI+GzlAEuBOCu8Xhbonj6
eA7lFBspv177p0V54DKSgjxG/5QYSyOej8SNfz7YM2gR45P3NBTFRD1JysBweWK489eeCnSfzsvE
wSBL5/k1jd1AU+FkOTVVyAk5mg5T57AhRVDSFfuf1vgKZ9GLaXpfDO4ekWAs3Z5f/KoJ7USYN30U
Wl9oCD1vNUMZVlFMYraclJM0ZfKmzFliOyT3E8C5WV8rfQ5sZtz+v8zUCYv3U3CzC0mbWlYZKL9r
Umpyle8uHXyl79jjQ6YjI6JO1MDlgGAdJQd5B6ovoTbmFg9j8uRTIrxWdk4C5k5cgpgHOGjHahma
hZNRQyjX7GyT6dbfFWJch4RtEcJUFK6NeGRor2+URAjh1KLQWREGl2E+hTerM9/z6F+druktTUN3
q0qBI3mqqSZu0emJaIVlIgGapKHMrK6Juz+SGn3F8b7Ozse4SMhiW4XawEJ0UC/+peYJptqdL99e
ANVzI+wJw4HPY51+uS7XLesICaSG904vnwOv6CDJm8nXj4MzE66bZr5a8H5iYiHFqXfULdxhRNTy
QvR5UU6RAgZpYsuBEgYGTmXLh9Nrr8AitHiJ24XKs0rrj+E4JZdBMu7IHPD72Ns1AQz8T6YZW8AB
gLPc1JsexdiApKoyCD7ucX7kR4PgOlXTPfhPjnb4Zd+UAI/eLUGOjXRVRwwoAOaEdkLbqdxXRJCg
6LrWFfZuyrEH3/CeFB1GGPOHktHRL0SSOMuASWzrjcEW/87qldPv/jetpujY8OwdxkDPpE1vng+C
dEoUq3yxfvRmhH4s2hPO6yw4mQeVgorGwquon/bFdaQag4pPfAvIQokcXidvNC7EfHQY+DK1fKKu
vjbJ1Y+XW6L7cP+56Wr9K7JRAREnUftI2YYRiTVfsmwtYZTSsyFf4IcFoxuvEKD/lDrCxtt4BRaD
fXIqrQTQcW0t23uyQkAy/vN0Tkqp2Zqt0RQCes69JWmxbIYYcFNouqhQOhEjKBCXDM5K5WFKlyeH
9motzvimcTBsGtZ5QLguea1BhWsLXryhD2nc5vPlbd7KA9cHnGURTzQYbELMng3ycFHj2zmrNZdO
iKjxAtttfqeXTmDza+7h6TR/pYbRpklKL9bE9f8EhB6FZuoorlM/vLofwqmyqNmOjUX0hv4diCQ9
MWjdMXfsCOUCTCkKVpd8oNXI6aZFdylbCcKhtBfsWWE/GxL1dgLs4DmJAaO9JSD4+ezt1m9bfnb5
jHAGbbEPdmML6Cx2WZhbgjM6HnMCJrEpWDEO70H5M9awyyanZGJStX9UJCuJEmxSMaMtNFmXyjG9
8VHHpiSNdAeroB06mT//G+i0kTMHlDVYbAfToTQUFVIuBqUA93J9jYX3CGJFej/58pbPBn5cW+ZE
WXdjLNTETseGKK36Lw9hmHY7t5IOAQXRrn0evw4yakafhrPaFnOeZS/GLyaErX06Vl3IWIzWrjbm
tIjo7TGrnMOM2acpYYKIzmWGrq7bWlK0C4n9T498mcVJ2Aq0jHEDYB4QUlRTjBtNgeEm07+qf71D
gtIqiRBjXy2MbBQfyql4chpdqOYwdU2bbQ/GdpBKCkcsV6RQhR55MOuibwbD+jppHs16YjOf14kk
FZym5QBBfD6PorgYF810uDqxKJao3VcWRvdwUSqugzumyDWMd1WKg5SV984d/jg1h21zytPQZnkd
15NT20A0AGZI2ihW9NNfvvdETJ6W4tMDagSndUz5FsNpnLwRHZxX4C7yec0hxZlsQncnjzD3bKiK
K3nh43WX7qoaA+1DC3skx6KG+09IlBjd8ldJxwJgG6ZSoGFZm+NuQ3zw2cBHjZUKcVIVAlqansfV
LpgpEkZo+g7nv1yUA8VBaB+BLP9R4aSF7d2QbMoOj2oUFT0sX5ihAQ05EtyFdjQAcQttFXc58fGY
ttsV1QJPehhS5AP0qDcfg2Duy2KMwA4SbvEtLz2id+WPMVYlovp+WJKFhVaKSeg7Ff+5+Bf05dJT
QfITccMZJdhhQY2Sx7V9bNiZQitUhsYVN6JSiUXgYi+8qBYDbQWGfrfoS81CT5kAs+5IoVc0PvAk
2pNYPRdOgWPGLfocxTy8kgdiVt7JZqayEkh6bA6iiqa6H1alRlpNLonK9e7WHIsXylOVS5GOA+fs
HoqQG7RDoKBt/EMOg6uLdI9k07yY4ZhXSeC/eDLCwMzGkVpKriDCBVyBlx8XT1iWUOPqZW2EW3sx
LwY8O7qjno0f2PU2EhubEKqiPdVOrKxuld7Z0qINvnxrHs/DBk91yUTZe0PSaaGM3hCoNfoVgBHa
2UynIVy+m3eDZN94w6Iqxfu4zekHNNAs+c1qM/5uiziXxrw5UM1y1KI9Wd/iFhhJORRvGgaRz5kz
X9XrLB/p8j1z8ubFzzySUOaShI20Mt46LtzZ6hOfiV+Elp4RPrrid5zS4cTunRtX/G+x7pTWaNSS
Xjeg6Ss16waBO7bIOs8Aisu6kDMZxboM0jzLcmeetbtKsmmMsAvvUvrZCe9juzLZ9duXbGhNOzuo
yzmSv1dlipC9V3c1p475mI4jzBtnQHQYBXP2Wz93Xk8Cw5zU7sGUVYzd7OjBujsymXIjawmU3CJU
bYI/tvGWPjohqvWyBwI0I8m/scUjenRNqfuSrnBztfPUZrrD87jtDZaanygLBVtxpxjV/+Sv3/Jm
4eWXMM1sjra5gmSwuTpaceYRzdFf2I+uRBtHt63oUczg717wtZH90ylot47FzizYS6KNeY/oNwx4
4UFOxMhAvTnN9wc7yxOPPZiKbgwVydTn40QksWf9qf2usWHI/kP/RZfD24Yq1DqScyiHP30U7Oqc
mTFHA/V5naDXuVPk2LkGIK4xqo8YAziNfDVecz6VYvl8B1WyP2bIkXMUyq0KCpp/DFpk/aiCYn4m
tFrKIWYGTtmCM4/UErk9rXohVWZ5vOub0aGWyhxU5k+lXuo5UuBgl7X/58y8xEoLjK54Q6hfLRwA
9QabGsGNgl1VKQ+AYDkRLuGJT32DACilx1TP5Qk8QIePOxpqs4/r5GTAvV2LIjoXJ6JLW/nQ+L51
T90/KY5DtmyU/uoW5WLx+fCuWaamprkjozHWs/fzcQesGFTNRDn6MMfqh4gwbpvHSEcH5CdFzggs
OjDSDGPW+p44OQmYyaRzIMxYCqZOHMQhGMGr7oCVtSp45xlGFjOSSgxvoL7b0D56fjZgi7kUalYi
qwbVx7WZKbZFB4wWT852RAaE3B2YzM/EB8JRJpAcnKTKu+vMquFVgC5MrTOV1hMGpwdKZaNhqXBO
Uotjb4BnusaNeTwvrdq9YKQ3MuLBezgEYQb8/SlK9t9CX3uDicjUa7bC1yWc8MSFQC15pNg/qhks
fXI4wNxWg7fjUzQwg7q7WxJjf2uoCtbpoGnHhhn6ajTQqWA87Ary2hPvbDy0aXgpFPoJbRG+6ily
50cxfbbxbvvmoQcwGP+NdcvmAXP3cxrYVClINaXP6coQMw3YzwkkeTRWJpL1uEHGDVBqxotS37kZ
RZ2iujEPar24nvGtSYk5CVZ0t46ishyFhPETUljqh5JezSFDZgwHV8PaddiSiJ+dN52YlRg8vtyq
tdrB2FtgIVR/B3NkXPVUjyUMSgC4xU6OZMlxWHIrr7NrYlkhoH8HcgoAkjSYFRaxG5zKBZIHXfQz
sXACbV3fUVCS0t+kyuSBVpNt12VmjTVlIl55+NrQnU7OtSaLduzAszDbdYvCg7tNf29HnnDYz3s8
U0iQX7I3IilS1t4IPHLTsat0iUDUfFFl80mBPp+JSFnn8s8gx9oeFrnTeCjIRSvon3LSF/KffjZ8
iTZf097RzvRrpBRZJycZxO0KfA/gA8f2uxPOCmGCefLSG9WR6zSk6XijCkceZ4ZNf+77HY8AuEDQ
Su/83a6JUUYArunl3kXKdEcZC0FUzP+T4elbT7OERlgbML8T6PDVMqe7ts3vbpkfH//ABqW1Bt3X
e5zB5hMrCU5GRAc0q7ga0+a7kYgst/oP/qiJ+Gwwdc6K0PPP1cGyrrR7i8Db1ZMldLBKpyyl5Y+B
oAQv+4O7dBGxkVHMqOAcuAh/NzOq8j0UU6OmSwP+Bo+wJ3YGZR0SgrsnieTMm3R9CfkWC2/UOCqT
y4DrDLpL7iFmtQpStJq8MQpkVHd4h4jNy0dsknzx24U2shJLUUuikapt1fH7gYJeX9o/ZPJobn86
ZUWT5Dk6bLZ6nDiHi/fNxFMP1ZtvYmiY4H802enMPFFPl6Sq8Ao9580jrjm4DhXFE7DYzyci71Rf
9w85VjLt13e0Ct/5233b80AohulVM1Ak+WziaYi3A9jRsKihvZoj+3VjSGH2CAbvISTgBQi6CmPR
LcQYX2E+2pKBlCNLUMDYRBkDhqbJxWoYLbGJTTySPJMBm0ZY+QUnCvEfypLPWakZasBkHsS351k/
BwBjv+O2LsOeVhauhf0Q470fYzrl0FyVymFMonvj3JPfs83k2ON2PQ2pWgtvEf366Jhq5ipb69Fh
z1emPhu3B6kcD8P2NE/9zFTRh2mtLIpT315qiA3MuNeuYffPcBlqdEEGJEOaF0y/p/vnvVZfkOlW
bWB5rSADe2iYVD9dOtD5HMO2ZaLLMN9MruV8UtOqKt7qbmwaSpqPKMvipreMBLmbswykXIagUrAu
0AHv5dCtN1fYlGG9S/O06bfiSs4FTZOQ7L5U8cjZnEzfStS5USOO2AEe9RfmkzbUXyqkQwQLWEq0
cl/OXpppsabsXItmfAy2giWFoLwLHA1CtY4CnKAxmaMMnK7jPnHWoZ0qWWcLsqgq6oI2Fu4gWtC4
NzvlNffjL4gNJG5ODsjyawv1CT2ohseADVktTwWZ02hDRX44N3zjlZFBr38ARR4sBhMjhcwpM8Nq
IU1gGjKUpjl8CjkSyToTH946KBhbqhKsAZ3B04sztLiFxQ0noh6WolBE5HdV1Ut3oBnZp2kREf37
cDJuIk1fqyvpG4lxMdyG0CTJH4q+eaoKU1IQaK2Hvzie0gQvYe7p1o7lgeF0i+Mz+6FipW/YkLUt
3K/FipR40ditoiMEjFh5KfPv91lAKC1gZPZKUNgkPL8dMbtdOJX5w3ubv5+e59psJ0O+8I8Xm61P
b2t+YR8hqjIkpRfU7zKaLpfxOp7w7S/JELcT9RB9sn1/+hit/F7fKta13QNpteWuJwOm7omgy/m6
bs+zYFmZjK9Ze6m6ejBq6Out9Vpcq9RFLvesZKeYNdChdkUJPwPgOd5ZqSZ5O/pEC7Tgz1EyLq7F
pnO58O1ANl3gjZA7bi5CfEJOd9/cBjvzjJxbvLYkDOiSG0UTqP/KyEJSeOP3j5fTvMe53C78K2Ea
qzsFAgn3EBlQ894cL9eGC4gF25ZpLkdUtvBwdNt3Ovm7jIU8yZtFzdkawNI0LgMKtlDkUzt+z1CY
vxQftkPWrrLl0M44ghdc2kM+J8ARaUmTimQcgrB19UrkQCh0FizDrqmi7TQJ796nBu0T9JleekOA
CFwgvsEq/fqp+9xhGB9chRCWzgTPAM+ge8HsNvuJeT0NnUpZSWBTd6ebEbr3PnSQkKo4XwnSeXvz
Eq2dZCh+uM5V+H/LR9kwM1g1WXFdnjttJY0Ssn4cbZaqNVGqAQ/cRrCIzknujCR8qPPmllUCcCoJ
ybMTZzwCiFiAfCsQdzkl9PO+LFpXisb5Ijx1tcIQuJJnEJ/mklFgtJCDksM9w1YAgfKyQqGKsmFX
jIjKB2j/kLsZAvjQMlRWUVfY6X1ED+b1VZ1vVl+In0G8pngWRisG8xJfZ9xH7svOOS2rGP7gc6pd
xtCc1HJtlhLd2/5PzFRYntHE/ml1ICU/HPKEydnVE7tHI/WvMeNI+yNwtCcfRioZ9W8nxhcBEaIH
d9RGC/7paNAs5U9I93pJilJL49GNt3PEhW3HcnU3a3mlTNASIsR+bFzaND9ZI1mFz1xBQlKONDwt
+T78DoHpayxJBW0Hx0AYb2K43APle03vcOtEgfwWvIedywzE+q85DX6eauIIwDwlHkpYoOGzLjlr
bGhu5Kz/TGkzEfovEYQ5rA/qrVyh7LHR/tuGn+MQ/TMo6kv6TFPzy9dnFcLa/Px5dZU4/10gPhm8
36O7v196Eq1tfq4lAH4nARH0oc6bAyiIehoVKmd9j3TokZrJIt9xrZCvAbNAVYoyMzmlccmAxi7t
HbrpDFCbddh/Cb2wA0ItPdzv/lJ1ce8532f69dBd/pMdvirbl+dQ+4qt7i52tWqRrRLR2thH1giA
Dhfc0RB3o/HAfomXC55Ir/2Nkmlbvgr4zSrxg51Ma9zjRpwK4aKq+3Ko41hqWPSyZ7Ps+aMqir23
kGdMVHaLk2hDiwZYmoWBCk9pQ754TQAtHDLKl51zgeHBJ58PfjpL9ALPp4A5NCEYQmju0uwui+7h
kPYT9gXuZC8JERb15anRZbMtpglNHDH3thiaqg0K44VRLg+uDvNigFovPwPZ2Gm8L2AjmjVccjgl
IF1u9U7uU/ZhzPXwDFQCf/g/ANDLukA1porbqwHlek2ZL0zpzT5UiCoQM+brtdfLBaTrLnA8E8M6
bDF3sqqIesMbSLK7/zdXmNLESQWxaPZPNHXiOrguMTfT2m2mEGEvTrtQ0GKblRdHRKASHK9OVdFi
7UW8b6zLZk/Txx0x7/0ppUpwHz5aEPkOcpgS296ddj6CJLqbXKF4wAoisL2j8QfvctSWbMuQjVjy
mzlgDA2/2iGKIq2KT+fnqajcKmb56uelF4wsXDyo0d+pCNy8kj13F19oxHr1+4ybpBwEeVbMM9j1
6WDpXUE3FO5+udEP5RtqCBwB8+qb+/ei9y+qeQm26LwLh2aNjKEzW24V70sePSRrGNqeFiBcW2mK
PKnFkQWO5WvKdYUZJk6QWq0ilAAptePFumJml0tsoXZtmwFKDmavstHnANmVvofTC8IL9g++vFEy
K0rJ2y10+IZnoo+cNy7bTEpPKWP2oVKN0kdP9zY1JZFJDhoBba4vevkOiXGkX0TgHm+R4qC3cp9L
UPdScI9DfrCKSJQBEWbyJrrKkepZfO5MBFQQ0Q/YOeKRV4iL5xsduTbnj8yYDcy/1eb3qJfEkSfc
19CXjiPJ6MPat+4DwckcXZ6e9tatEUbyAR1HpxTkxn06sEM+eOZYIbc3iQiW+qewnrUG0o8P/fhB
KnkBekKse9cpeUwK5eIADAXqndgg45wlu/MRpToKr6J3OBtXh4d22PVijnbzpmKsGV5dGQVTcVVH
TwLXNAgqJ1WeiVzrlhcQutXeNeC9qrOZGZllPLISdo+DJNQcb0Hm9jbf7CGJJKqOYCH4eLKWbLtH
jn1tjndyFYZuTOf60e8l4IACYt1cndUlSB8JzZDK9wN8PlOrw6/4IW7bOHhiwki3N3OLhx3wxXU2
SYyOxztVZyacuJfW8GjKtW1EDFkXgJINFpQbITZVpFrUaciMAG+35t1JS1PO+xU4RScMohVUtZ5g
/xit6mU4bvrzJTZhIPeD28p4D2EpdtPPb951Mp0kX1hnIRknNTuP16SDGglPktFk08fx74T40xC0
xbqKfF6mfUcwb1CZucRMe0ILI3k4FTHZmAEVdv3RNztwQnXMseGDsANRC0/2Nqti4AJ9wiLND6JG
j2gcE9CZgEH6QlKv8jt2ec1cmd+rOfNQll0nMylkNGfCj/tUcDm81xK6GutYza0sedA7fxBFJYNM
5bz+6126kfSS0WBeOk6lkFhOh9vZbpwzowutLkl86vKAGMW7GuQOr9kk51Afpd29r028Cil0MjV5
xcYrOnd1z3rcOnTIv4t7HtKDhnB69QCsnoa9ojuhWY9BzVjda+Pzd5bquljcMmPF7J88PTtcMIgq
syulDB42ZqNva+ba1q1O8KD/NKdGs6HKegfxf5ed8sjhgpxCfFNivi5fmt5SuuzWsOrBIAOzL6Ij
jeme8H0iF9o86z3UGBKdDnIb2vJyttQOXTCCcooY32/zwIhI7Mh/Ap3Hm170uj4gt6YhPuXe61u0
uXcVr05U8hANdTIbRNKqEpnv2pZZiea8JcgiVfgjTSzJWw+k/EO87/Ok3g4GsiW7OYHwUDjgDv37
PWmZdJdajfG9E6s5D45EyIj9c1g26f4kdrRMdMAnF7hskbRoOLc7uiDIwkU/TzK9jc+dzyEofzyc
WLMLhQLIYfxaO13VBPxW0iWctyGQTzpz+ztURYmuoZwUSWzx/rQFg+q3LfMF9HBWjxj/bC8cyICS
z5WvD9N2tuE6uEiRsCQshQmkMG+bLDh1Zn394af8JJ7U5R+Y3se/rQ6CGnmjMaBjmxO+VCV43O8h
XT0EgePND1h70/PVAPXIQMAvsPuUUo1PlTMRaGgeXU9DCcisYBs738MSLiC+3GRz9I1YBgrCWqKO
Zr2D4zxaVDkJLQTrHQpE5I9wREfKrOB16EPn7jaR3kUi8h9NOhAXz12KUxpV5PM+lh7eUNUkU25S
TCXCjq9U0s21VJ234tFBZGX7NSIHho0XdvieZ+wHZgZ902jKiXuwacXBN2llhVhJUrlamHPP2NCY
9Y6G+QnJdEnK2iuM9IZrda9lqa06O/tAG9RkOMkLBBN8yTUXOggCbjgtir9WcUuzOu1kOIhRtIFA
gtIAbzbvKt5If0yV/TN5GzGU82/uK1N0Jg0qKRzRf0gjXMleBDVEYAfixMGFYyapB2uqAedP0g9U
lsqFc2lbMCf1TWDLdq8+hDtkP1k12nEN6WpD4LCHxMaUSwiSIfmKZMngA6Mirp1h3OomWo2I+wL2
z88Ym93GU7VpBjmcY8HJTnGNoJvrLEfVh/pEsYsZAXPyDeF2U136Ie5CBUKK7mu7PVLu5zybi9xF
pi8nXjwWX4C630qRSTN0O3bJFGD7d8NgI1BTfdjwPjqAYMq9S/t6nikdI9524/6RKZHXSlhwMZXO
eemMVll3N3UHSSKG4Lg4mFxHcW7yYk2wjJD5G5yu5FRr25uNKr5Z025Hq/7NrDzpxczr3ECQAOSn
Okemsl+EtKciy1PeZI8wVeZ1bQ0kOpxzgy4qi/prIQuITy22ZLNV5IBv2HQ98Gz2ogBB1wHvuWDi
PgcKrscIoAZJNedXY6VyhD8jWZr53/rk/nJv1cQn74UoFMxJW5Pl+U3J+dkVLzQHloV/5WfVqqJE
nJIRicYX1eIRuOsKvue+kWMdk1uL7Q2RP18+1CTK2Yd6OTuLlbWuZCQl/jTq6yJWsLg96GAIMHc7
X6/u2WbYiniwm9UP/x0L8JiTbB7f+4uAUVXo+ZuE6v17aJ0cu5+XlOflksmT4ZfD4/pMRnqpI2/e
Azk5ruFr7vswOv6TjrPp9zIAgPoqKe2Mlb6HPhtaN0Q++LkCSITLlKpp1Inx8hkmb+GF5cT3021Z
xIxWrNYQqrK6se/yec3QXOn6BxZ2rhwNqxj1WFus3y8mqPvjmz3O8a9zO4me7jcOUOvJS+5vP++a
RbF2GSNoMrj7qYx6kU6JH/qVvNHt7f9LYaCuQonHIRWXmpisDFYsP2CXXZPEOwcmTwvEjCR3Rme2
b9JNpDNK5XkuNKHsTjIq1ftOnx3S+B71qZSFnXIPKRFZsDbPqvsqJQHG18ccGXCG2wGOzHDtZTwR
tgy3pgocNoNZZBRPL2CMewaSM707fJrKP3kXhwbyfcGRCn/G9XBfxbHpcGgPU5go5J7ZsSsisj73
OqyLn9MAxZ1W/UdCLv/2xsV6q//xpKv0IIB95AL/PWSM8UrRHTBVHNQ8gXEoNUGM1CVvr9J/BpgJ
n1q/790P/PcwxDlRa2nzIaRGtiWimD3Fedu2xlQol3hUzerrnhZ5LoZuM+A0pqyv+EvX9n/KthY4
I/aPD7iMKd8fOWX+eRnQBHriJs44Ls1fpIYGvuc4Oq/pbC6A/6zAfBPROlkQsxnFk93zAqeqdOL0
YYfMLmvrqYD90SOhh1A/SWQgRIHrO7+ZdBnT4EltSB0ULo9fABe0V2kVHVk09Hw/ASD5rod1lgWO
jYKcS7PamivEJ261cHpHZ6bg4XTbYV8+YNhj3z5+pVYHTKbQ6ReTIq25k5A+7MPZaEQyy+g3PrBy
9GtY1mDJY0iLYnAxJmYJyeY6BzQFXCAkhjQuxRcna0XcvOZ29d6EXupvsR9WJGgAqrjg8l8zccR8
o7BaWTtYsx5J+f+SQWPGFqbqeptICg3UAv1MlRad9pSW+nGvRJJJ3VuAwYMTkSSMWdPQvTG/mS0W
pz8neyJioEL5X3mDCvSZv3ydw5pqbKkOrXw5tvTGsLlut9zKYTObxCHYVTZ5cudFyVan/lWwu0QU
+/T1s2OxLkBXbp/+A5EWC8JMpLijSjcCBC+EZIMSCIwiyXlKAGqsjNkyR2qQ6pS054j48eF8Kk19
Z5vQqi6HGuPFEyWgPxfwwds2OQCbFirYZrOkHtAgk+us/8HcadgLTZ6QzCU37WKPhP5UKtt2Ys0P
5S3AFV5gEwcZpoqC2hT8tPrtyh6VjhPcMKNHSJIo1HcqilUyqzlEGNWctbbknZRsnZuxHUGpY/IM
CXpEG9MoVW7GUUGDQsG+/kuK+JSkOBQhLThTD+LsVcAXs94BTfGy8ET+szN5IXyDkPL4OJVIUv5w
WeWImZ2b0rwv4H4BZDQPrm87YTH8B0c4KN3T4thNLwo4PCfyitN4CClXLPKj+XUUEVkV/LHDmoHN
63+Ugn0iOXeHXviDcxv2AepyEKjxM8+90tsuRqOSX3knrX+shhvteBNZh4i9nXjYeZ+c2o2vMQIX
MzXNuK0JJfSmzo96mvbgZpNfjYWoMXvDt5ViQ7KXA69elqC8gB3z4+6vShhET/iffnv5PeYVKt2g
CCepfbb52NBFyjwJ5t1XpbKf7R6UC61SG+APYhfOZN4JI0VgkMNyvUF2WnAmp89KglafSxRl/qCh
QbTw1YBcecbTadBlOzQvxVCF1KtLcpPQiVvZ4xe38GPE3zb3wvfIRN5ntWw/qAxf4Naj+QTwY5rh
FgfOrgETYpby5a+t2qMDZt8hdpTwMVtpIxm8uKY9Hn7sL0yl43pwG/nBZoxK0aMCh/GTo7ku00SU
+WMUBkOUmrrtdVTla4WaarsYqJ7J0OD003aY3XOSyvjilMsnugkmWhhlfTL/2lBjiXEK3pbMAc8F
TbqlyGrV5fduB6KxG4neoEzGpq3Mdpbm8cqDIayirgAPaU75tFwVGal4x1c6TZgsX2cLqyeKPxo0
umInFNUzbAVQg6xaV0xaimhr2JPbfUx6Jx/7a2QnTqMgH4xaIEBY8hfcu9yxUYhNiLO8Be6wswFt
chgwCqw6ov/AYxHxyXFrkO7+wNu3GId1ERHKiiD+AETINY+/D8chy2k2KidiyJ6lEiQKguoZjD0B
a1+69iGFAWz78sue7RMcuVjz4YGXmnPEOBVNM7pA2rXMvRzb5F19tykgwyiHw8SMz965qe78Quu0
ISjOwI2md5VsxSsBTeKqcTdRbetivuZZT823Bzhs1aOfFuAs1C3jyT/2BTg+SfZImK9Lr+2b1cFg
gOeSBzee/zJOqHdRnZDSETgEoQqCPwFV2nb5mpMywvAbS5lJthy17GqavUbq1cs1eCNNuP6GySMm
r8gQLlKWyLltnHuNCZQD+7JJaPiRnTEEsyGZYXmLtjB4Cdvh1w+x0ZEc01MScO9Wag7Ry5skThWL
ZCk9B1xKdaRm3p+L9oNSi/XgqSa1kHlD2EbpQ+zlXptDP/DWwKgy1BpxunkiIkrlMC7m1lLFcqQG
uFctbsSoGAAcmUa6hPMzz2f3oHKMbkf7a84qpHBEXu1QCUn1bhyowyuO4TFI/sWQ+2yawb6G+MyB
FpcH7WLpsZt4eN+xx1+0Bs4AQqEBVsMQSFZ+1jwOod+ShMxtkPEj05aNhvnIRB1WSMtsicXcCCVY
Snp3neCK6LnmetM3cZZg+Y6GJl/30Ax2qc+g/tDiVUf59QmNLeBzkAcTjWRMWMvN5lizPV0J2pqU
Ec/wFZEtLz10eUmHrgrYar+Bt0Z3bWnMtPlGdwNhlxieis+KapQe5G2b3EXWb/nIfrIhXtsrGZbO
HhYA/32nvSPBVwxiusjQ5kEtbeeBiZxJuX8NqdN5fcEV86cwEbdqKbaungjFIFxbY6a8i4t8/3Up
IXZbO/lmviGWV2eisiPddt4UUZTX3HsFtENxeGF05M+gef5iB5tw/KNl6XSkSlu1XHpLtMd8DrN4
1fX9MWKg91LMWshgCNuYTlNWppYW7PkEvJd5PHwtcvnGM+z3w9DZZg4A0LZD4Si3Typ4A4yd9YvA
96cRTXCSO+4J4EBrkSyPV8Tcx5wITfFjZ8CVkb9MvEHrVUUQtJpcQGY9k4BjG6S2tA1y8/CqHNCU
2Io30OsyAz9SdQ9liiDYZVVmOyPDT5cayq9aJEh48H/C12+F2kX+jBLH0VjkbAz+LSNL3NEKueL6
vLLKKCLFpUUvqoJ9WGrD72i0oZqIiRMsh+zsWfm0q9CJ0TYyEyjsR7ZmUTcyXb/t6RxU3CtoTK0w
hWoJEK4v6Z2UhyJjkLliyGZwZuR029hGAALBdp3qgwcD32OoD53a7lKvHsWzbSghVNnhGpdH0g+l
1u1oLWPmN19q2h+IajtB3MLG6kJYPuVbebkt8r3guFsWwDt1kTqUqJPD7nldoKWECNU3sXJe3bGN
tTczf6qyllbLDLiv3CJmA0FgGwHVTfCCI3pnHsdAULAWdNZEqQoS/Pswgu5SSN7gwyGpWnmw3ltF
7LNjeOAy5PtyROINqbQwDSlBPwXyKzv1Hv5IIsJzDokNe4r8O86ZGq3ZDgSArM0FrTFg18reLiCO
qMfsdjEeZSDaiZpQd2nw5et4e2vKOf2yrGl3Tx6C+w5yl/z6lkYaytVVyRC4AVaa6sLRpoH1XnAv
MBQzF77AisZ2faSfB7S6Dihk1Scyg6UMn3bNQ8oDQr3rLkihRV7BCeLOJ0AJsEmUIrLQUmS7MxXC
Lg47B78AzFwqFsImYQJjXv84ZDao+/Cl0DcymPIraCqJEF2khUC06Qb1N0wC5chmMGmLEYzBoKG8
ZEL2r9jkZwFaSMW0BdyqpMeZoon9rfZ0Q7qZmlsxUBe7ErbfVYzNoL0owGry30HsfbDNoC+wrilJ
ec1affQGDvJB4OxnVAUOF3Z6Olamt8AHAWuuSirlsN+NxJ703k/4DKffL5TkTV89uMSRkNcBs27E
TCTFlXAwW8KcLUB63xU/F5AZa7SJ+Rk2CRwLcQ+8ksdfiuxb9X6xZhq+Tkn7n2Kp2BMTdB3yJjgN
auQENoTvpeSt3PqkEEL6oMrYorZZcCRrs34ECQgA/6FmQM63LEQRSCFicvX8HhrtcTgk7e1U8Svu
ywWvLaViT+yxaGrNJ36a6Fh+m02wuMbu+07T3PCQfqTB4c1yLMcz0vUcBDrzR/yPl/OjdPPRWpsc
Xh2bmNsFrXZyy/6fNv0+4KOQnaS8YSc3jwa6AX8m78xFkXJ7fv7XLkrVywryJva7EJaaFhC0S0uC
sL8wx6ZCqHC1ImbWzC06bdGdcgc2+HfNzcMc9p548QfKveJU5bcszMwYnqrb9jhwWMwiwytdLRvn
xy3mLdlt3rbMsJv/fRC3s4tN+8pZlYrl1uDG0LhUedFefhaQd1kHe+5PDgnA6UchuRIu5k1LGDxl
hp80IwOD8rO78L3O71NwZGOi52FcyK1QIP8Amnswg/hztg/hFD3iTTa+yFWKoQMAnx5hJ+1Fw1es
bQoEXdz4wW3VqyXvTsS5Tto9IxH1SSJSh5UtD7mpY7kDzw6H5uR6CFmHuYi+1l/uOTIvavsgotyY
IfbFDZd1taKRGnzYG+yuGWpsVTcUMYK3iMWmeTsl5eRzIbZDz6UAML2ED+jSc0bwVzvYHHLcKy3p
7r1jg+cX3fVPdARpJ3LnRfuCXv/G1418xk6jVlc6SoYOZr01blzBkNlII2yPhxFHcv5MxgftKasw
FiaD1A5xn63hmkiK+s++uwRhsqFpqtSw8xa8g6bcpClka1aKl7ywvuXIE6wsoagRILHqJZ8tQwqH
yA2so7fbVJtHhHzbwoE/R5yGtmyF+fvdEvUGBKEUBDZGRh19s5QvUntt3UHDvFE5LbOhkYcfSA5y
Wl8ijIvHqU9FoxtG8OoVcMXyMfGxRGg2x0VCIvVNf/TCjhm7qn2WjcBEOa7sMCdEmMan+PIF1L7L
WhmLIAdRAXS3JGwZ619nowjAb/yNU1MoQ1NVSgTCW0jMH2/1ObsEyCo9YKW9QG2WPTh43wqpyDj9
Fb3SslHqlun1oZ3c9jIdoO48A1F0QJ3gUPTpvg7MuxsWX/4s8hj9OukhN51Ltx4HPKsmYboUHQla
pDf/2UeyNM0waH8ny3VR60J/bwMub0nZleJ5T7jD+9L02TV/tAHuQS9QJgLzvXxNm75nElxQCwgd
/rBEYGjspg84GMdc/VUmPqYTkQULoSy0dlWb+Fg+tTRiHttu2dUcriMRaPyVtPT3A72FtleE0sal
olofANDlwx2ft3WZX43HTCzIh6G9V4G3Ik87hWZiKJf6Q+DlvTEHdOzroFvEYqHN45mi+Oo93nXh
FSywatI8fZYz6DKqT6WsmosJUpTbCaM5vBej1EG3+tKUvig3vCwrkIEnorFtXglM6c1OwLq5g1WC
FirhHBJ2q9Uc4x6OplL5MMwHXUJU2O5kbKQrOyMzTVZgf46TUvOYF4Q8+PZQJduwoLKVyfqbBZfI
acy7B2o1rvwI1M7YzfFUO/9ZdKFPnptcmruYZaC+tN1Ss0K1Po3MkX42eIBxSRSjkd+h1ThAs+rH
DCUd2buyRXOSm1qyOt/0p05Br9AZbI/m3KgiZ+Vb5C4I9/gYgdduDis2XcLp5J3+ZWwGcFe7jBr/
VSMAOSibs7gt4iyk+7GIl3YYo1m9LO+DtmnUPe4i9pBzV5R0Hb2fiJY/me3rdnIJXwevra/kc87e
+lO7ThQxLAPm8PdAXyoyYGT5isSA+lWPIoLVHF3ECaunfxF8EAc7DY1kmlv11MbOiSL3wQLij+jn
M5fiHMoxP7mMk8iT9fYAFa4fZgmRyehQ6Z11eipTfR9VzOuUzi/20dzOIuanAHMl0eZJU0i45ZvS
BHsfkVXVaQgGSCPQnLlIk54jihm7BrF+4NWeFl4lQc7uH8WQO0APOPtAaCXhKIUfZB+O6s4xVB+2
WfYYrebJQnaOBxkxkzfXbKtDYl/I7pRMd2x27YxgHgrSxl8b+VqeT8wZ4utu5MVf8Un/5RgBbv2Q
qWq/fUpAihrR/svjMYIPCpp0n14OQJKIvVwnQ/yfUx28Rh/SEpmbWwShrJV1TCs9VlrvXGU95+Dn
xfcX/b+WbLQgO3gzVQx4YF2kTTFOttg9BgDDYkAXQewIMp+bY0LRjtYCHvsfLWiIt7NBpXh+hUwf
BAp8doqg0KTK7p7en9jS88PMvB4ArsRxVkl0Ahdej9Iuuja0eeP4HuTgocR5QHjTGrzDpQIlWf1V
plPd1cxO5Ko9mntnbLD7AOtd+Th0QG0Dzrp49nzsA/xxb8F41pBLhU/h2eXJbTE1CDvtOBtPSdVV
Bg2unUxegWX6mtx2v5qj6P+csGu9pfoxDi05OOQklTMtWWUTSxCNn0WmQtkvfQptcIKKn76j3b5L
RVVv/lBRmmaGiZV55q7Q7cLNz9LOJPO4HbzMBpJe2C8vkNGtGCARylHaFGhYkDkcYNMC6aMwn/Ey
vRpyXLycQzE50ceVq0JuTPxnYWBR1v5kLIimcaF4zjECQX4boZPrPsz8RNi2OxdMGQQPPw3/PkM9
ya2AtjffjtVcVMCJvGIAsP4zBwEyMU58K52ST7+J+iC5RYEAwRQKHqam4vfd0qwR85/Zx3UBK52P
PNgRKInn+L2Og1R32IcrqJZOPPBi6oxBRs6BJUx4YSX3cfHb9X8tZ1FPJkeMx+O8GbJGXB5+ytOW
XTiIiCIExql3Tjl9rDBC6YVrWLWNhtSvLSjMzE6pCMJta/3to5HibODiX1CBbj8TI9EPFZSoL62o
bt2lKpFt8hcTWTBY2DBpdgsYcaj8nZOAiYFNHlEKjEnaURKx4YPUtRJUhzkkJqU3zSjSPfi7AjWg
DxyvF59OowrT5WYOI3YmJa04GqiNay4/yBkosKqLpy874lHdExoboxw3i/tPvcx4hXhtD3TQzrZR
BT3gmT9jkeLorLEfxPr20Hag53YW4Kpr9jEzJevzXB5GaXyadBgL130AdMRqIb1BdsOICig9GCFr
eihx8zyUK7EKtRsXk3RfqPOf1yjFcZtcreYEF/VFQS7zXzdz3Ko+TPeNCp6SRckBZ3lOzpo1o00P
9V6eKVJaNf//C5Kq632IxGnfd8zRUk2g5plOKUkMTdJWTpE1fOk7GvUoKyo/i39TWnqzbCEJfJiQ
spvaL/qy70fFD6m9dWY/gnR5SB0Ei81RmMr8lWptCUtroUn/OoLI8Ty7E9Fb96ou5yLCVbrlg5Cb
ILjRsXkYvrhOB/BASZc/LwNV+uxuIX+0ovke7etWNQy5/2AyaTgq/4wCUcZTdzAzaLmNECymCeJs
F8Nw0Lyw4DveKKM8vBRQdH9/9CRTV6GLzgbiBO58ITdQg8c9VJciLMnaDlI7oHBfGar0QwhflNyU
SiwFgdu8wImQDUh294SbsQr1meDA7LE80Zn561jJKzEw/MSbXxwrOI5tC3XACi1XSWYCR0AHb3cJ
sjTlKxSxNvA5acA63hycFuUwvl4oOSeV8Qls2iuWE6TOXzvDv20bZ5ecQpBmBmlCWmViZQBqRAbx
7pVU2vnnND3CVuxG+Q4HxEsrOIkmuqxxZAVdk02HHgW7TFMN1EXvJD1qYwM/sbG5rqDDLY/3FTyi
3uCamr5S01g7ZJmGjs5yqpyyQPUXXdxfhut1zYk5dbpkoi3p522I3enSnOYaq+rPZla1aiBiVwoe
bDVzCSm7oD2iTAyVz4o1jN8Ne3fUnrHBW2WJgbfEXsMI80GHEbU4M2z5cpU38aj3y5gXoLoCd2YF
EdqbE0q/UxACwIJ7h5b1ZrKczU0mCU5478zXskj648V+V6vvP7Ad4Ej/8zuHyd0RuHHXkldZzdEc
jYVcBLXTTrdLa3uKMcV3l7EhMMcFCCZXBqES+erYZRBLascEBtjir3tb/NgTbX1XuBa7G0N3mhM7
PEskLCqIi/SxZTfHPzyY6gZfYAy/b2XcCZ6MiCrNv1o7TyasbwldxAC1zadvv3aaouND3dcMXnf6
EEONNvFRRhIqtCdKLLnYSwQWxlg4uklAKpS7k2GNEM23l/WZV+hXNuXojhgSzlXUmMIfCDM8/qEj
JC0l/Cbk6xduH9WUFIN4g8hB9MI4bbsUVq5GrwPqOWRuvrSFoETEA7qMoTMwDZv763wYb7DkmzC6
2goBnav+VzLmSouJDgsTCaZGKC+IFnu7NrIW1ZAOj9upRFcpXscDrRgpGwvBCfEHWP7sksSAde3N
p2boI4GOmrGi1fH1mgPFK4FkdCO8NlFAN3SWsRtq/H9oFM6SV+/OTgP8Jj4RIHbmj9q1Ho5d57Uv
C9dDa0X8qL9ght+fHyjJlDsbRZSOtJhQB1P8f1KhBLEqJfrNv0YDPMmZJeYnQ3dflLEN8/yyR6dp
BbqkS8obf8XxAFwkPt+xqa0T0tIFIjUkvqf1tI7SQZgzZHq6lAi54AtF6ZUPilM/3OxjFcMKVs15
yCSfD33NbvlQA4CktK3E+vsE0tgKveVSsXJ4K0H2OfFTmAkrrUgKFx4d1lBJQ6NCT9S+XsHhp5Dl
S5mTYxtwHKsNLZyHneCEUVxUMNsK9jrBb/9LhY2zem9jCocLiUhh03KQZwXFoRCcrSeTdgJ78zfz
tWDIcKZ2Qujx7ibukZWeRYIbAycfxPpQdxNEsxYUrUZWb+3Q5UVCi5E2181LaM9JcK4rKDgsZTTc
Cj5XGfXrXS/NaGW7frzqNOJ80IcIXjj4HtqdOtW+EHBa0e4eMzNPv/oHjTmDJ2FqOnqkqyULI+2d
OGTIcDz/4spXRu/IIYzjCw5vRy47xvIcU2Vt5C510p84IrbKafPDsboLIj0q9urEBmFb/+8Fj7P4
4WvaifrLxD3jJIZd81x4U/uJj77N2sPFlOto+atOnbmjVttzpL4DiuLQ9EpYIjFGi+S6myNKNTPL
Z4OcdsCzq9t9o5nu4YnrED9ut2ow4O1BosGnuCKRTIyetT8lFFge+EaVaBMtiUE7jWxg9/9HoFKH
bjSqsoD8GP7CDfMNL3Y2OBWEOcgZwE7Z62yFn4X4pum4K9HUM7NHHrOfK1gABPgd9xmL7JvQMqS/
XOxdAxMVXuvCyMd3iker3RklDEjexTq3gW8sSMIHT4V7bVvd96PMhp5BcmQ87laxRtMj+/fYeSpd
PmMY41NFIhDkM7pmrzuk4R5Kq0qyoIhcJlwMybU3zZKgHgRPnS3gxbbYaYecGLzGxWlbYV/d4Atd
CX1lJI1u/4eCU6b72T23urYIBk4J6iKryC97tSggQaG4pGsQt62YHojXV5Ps3SmmmVWARXVhY0Rq
QBvbWgh3SWtqgVA3tsC9Z2I0Bkyt/Z+KfYmufwboGoQw/3xxdYs6nppGFL4tGVfgkRYpGhXKSYqZ
Ldk2f+3nE57mFJ7999to5NLZ135wv7QLmcIxShmG8llOd3kDYiDd7insP3N22iKj8VVysvoNZ5jB
6sn2rEg34phclf3u7KtkEEc4do2oHKB3VIA/+NHWNkftImomrJ5M1o/u51gTIx0XOkAfLxBKXBul
19Cr84mmaLAdlgnS/GHzlks4ih+sJkVLPuAp4SqP8jOKap5eUDGLa2FsGUXb+vvJum9hfWpjkD26
BtoZF77EGz64sfah8gpVpSy3riBUPXKKZjdKzpx1NVi63v/woPXRoJqhgUzij6q9PH3ltvXUDgYy
gVebRFWqISpvH0xsrT18LnJ1Obzr0JFHOQrcupBwspkKsM4BrT343KUDFdWJAaInJmt06BsO0o5x
FUJZv1xiFQW9ovbsw5URj1TDGpMtIgHCOWH+L4UJXAxltpn5WBfJc49hvx4QBDXphq4XalNxSbW4
Qj7cOHlC5aehUgOpBlGly8JZKYMU1ndHH/uvant0g/5275MyqYgyKeK9OwAjgU4jRvih7PTALQ9F
MCBeXbOo8vJqzrrQApaTRUdTT80kcmxQOOPF8wQQVdAqczvJFLUtXqR2ocjZiGrwm8NzT4SAtuzZ
6CY8FVCEP4uI9p6mjYgXna6mY4ERoE5f+C5UGAIan+xc5PcRWdnOaauhpjHEa2Vtf/gNi9dyjuHH
+pZUTA8x6lHLDtlMTGT7/IocMDl4EIxUlk3bCouoobbPfauoD2hw9n0LLRoN1FNex6SgMdOX5Etk
0TxspCdz43Dle+Bdcslis/nVnB8btpXh0c9pkVDp++ENBHPjPzlE6ObUUJrjFklpVT4pAiKdJlWx
drOQqxRoHjfA420dWtJwNpYdm+g60Va2+OO/yUqrCrnxbHdTP1AV/GQCYL7+1m65baPye0cQeK/2
xKnaGkWGN6AwE7BNL0x5BWXNsKAhy6BLeQVWdWD0JcIc4zNnyBcYxaNhECs0kpJFpnIrF1QSNV3m
jWhO02x6Tb4xPxJ5nYJ9TvcJzkTX+w48nuHBDCByjCQaTR4U1/q7CnNw+ou198s4tMXiVacY8z9Y
AKlc7s4hPu2jQPnNemgIlB/eP/4nCzSrES+1fEHJhp9BEkbHZeG2xPr0hy+JnjkBBJxl9O3nYCgl
2d4pkd9Bx9dftWK0PZ9GBwehm21ulbp9kA2Ue1pwxw4nhf6YPuOCVPvTQW2h5SEdwzd9wopf1o5v
9jvNjy7eAi926ZznHBhLarwLqHQO39wrOB0j44Sp6cVszYuvkzCZw5njqmnneJqo7sxNJ8mbIcNW
5KHWXsgWgQRK/OWuljCgjnT/f8vfcsAcoYjBTLMCd06CvcWhi7RJ2QbQkF8QlVjw051RHCetsr6R
xzaWb8uYuMbh9Tdo9O1E01Ho7MlR7+06OXi+FPQ5ZJD1UqSEwjm62l0VSVYAoT26iY+xucZ3oCd+
nRm4lMQINdpK0kGci6/uNeRgwgdFlufE1nm+oq0sCx1ct9RIsQ6zMRpfgQ/9556jv9ogVwUInFDk
7m7gl3lVLKtqozCDzPr/sbOBVroNJc3ouXH7RpE86rLVDgSTwM7PcNqdVqtpCsLxiWTds/AJjdjh
PVimqhhFGGejgRCYJVUkzTegGJZFL/gFxrVxhnIzUbfk+nRlkGstCWO7C76rMyyTYxUHAua3pecL
nhqwF2QVCMY6xslXNWfutG+EmKnQthQ7Y984AlJplNe1ab3qCYru4v60+M1Way5thHXv/dBb8+6z
W5m3u6im7BVai5yDvVUxCjhAt4q4P0bLPmDMExPPrwrpFsMnyYyyjVgKa+P3Js3M1vZ1NeN/nOsa
WOC2ILbqmk5GYIFiMdEG66BOiONBR7CX9koVaISLBjp2xLLuLpWtK8+i47GuWY+wivmLbnAevkDf
GuRW53anoby6PMmrTdo9zhPP8vOG2xkecNjIVeQvP1tx1G7cCSwkr8WWHE7d/X4TviEFSQdFHeZN
gye8VXsSqGOCi2/7Tz9Jj3X/IDQnbIZIcjmNJF4G+P92Vtqw+vB/G0hUIZMazUv8BcAj7P591m++
tg05/rAVA5quGazH95rTjwAcINkeIN8Fjk6pOQjdBrHMZ+Bpq2Shh29ZDFdMcbztcX5ylo89MKIc
j5SHcb9mW8qEptAVhg6wm6Sw3mLim34rocz8iSmlCWun/h6sUyIkgpF21nYpFaIAEvWn8bcB2BQA
FgZo+jUCRsFqdpJpsjawvng6hcLW+kpseUD/s1ewTneg3BM+FpMW4h+F/OZc6sDhqv+eXG0dwHva
oYdAvI9Q//RE9kGVij3PlIfwRlkrSV8H3ac0CixYcnzuAt5BAB9Vaa4++cCVIYTdcVlwjZbrp0Ex
6dSSPsonMwMNHZgcFnWQVYzBUOVigAYVsfoHYNewqycQBehle72woAwb6uuDS+B5xUkYupfO5urA
Xwp6PKIVySqPnjozdheWR0tcn+eq6f8+Uu/TqjHujEywehFvb6EiBBhydd+mU4/3rmRZzFT+ZkNP
R+mHSDoSxOXiIBUZb7tVa9M/Nvmtbr47nDUNFuqVVloM7CIz1/+XmROmaz16xnKN1uD24WmPpBME
/h3FEoZOAABiFLj4SFfucf1vB+KFKDKlWfqBMJ64KGQmg9YvQyEQ9RlKSv1reduFlOza4FDEQ3Oa
qt4U7zV00LPlq6l8TzOcR16Xz36tz78fRoWCVDxYorfZ0gE2awc1lBMzbM5eTZteSRD70FJNqR50
FaMoSeE+R/STY95WLJG4xABmCyTNLIEjv+DDaVxibvHI2TuL9jgx5OvrTslUS6G9OrTkQhggvgNU
dwqyo9rf891Vc/SgrtcRlnMVtn+U26P41cPNrhXM7fO4C0yxfPq64s8DLHrNFhnLCBd4bTq7gEYq
esv+yTYYEEkqvxFeAnX1RQK0J85f7stsGQYTdwGVYOyrgFTS4NqQkTphWnyF0oyd7nvjduyIoKLp
pvp8B0K2gPIbWEOPySAbvSFTgxXaaQPzL9+xR994MV7j6xCZoOsRv4s0gBKN/+gO6g3UlsIq05Jv
+1wIYiCdXw16izZlXRD5D3XxnFbofSkdIUQj5dlyo9FsAsulY2TurXT9wCDo2TyNNTEVckLVG9mG
wj2IpsPiQVWVQU07Fph6XENyrKes1m7cC+6VECOesn8+BRY3p/D/BK2Y7foW/MDhoIFCs5ZsiCxN
L2dmK4QmdKX+9E6aupT9kvpqF1/r7LhZ52YkRW1hlMGY4mT4SPlCV81OCw3bc1vItYgVrc58xpTe
kJQ5zs7PS1IkVajhs2gi/60Wpl83jDfDqNoTvkb/FkY3zLzIjgIiOykS0LSQHHisq2SaMvUzGBam
led30VP9E+lkAYg/3QD+jemRljTLv9cVMPuC6/8I3E8Cpu2JTCqaqQ///C8byZmEeZ3xnmMbjtJd
k5aTOjKmzCeawu8spypGbDgYykIw8b1pOHXkFzyP9FL7UwnQfiOMSProPJaZ24Sg5lpEAUVVfWyx
E+teqbo+IOQC5qtDI+0U7l6dzWYxDlcqXq3go5sVGGBiirz0dzhwob4yPtYKUcxwyiwd1krUKr9u
JUFUnqrjzEFNAtC6Tp8TPudPwGJdiZw4L0bioW2F+JAkmx4FLsb6lieOsRVLpA6IT37+yizqAM9w
D9E5c3m5SCF2yfcc/PA3a+hUqlWrQ+uZF2b+RKGd+Yzpud6sPahxdtUewoNJnZbetEhyIYkBBEVb
k0rr2HsyDbydy1GUYEJqwu1mO7esSLtrEmm38DZjVobsUXxorNgh+0rFeAKYrIBUVYI387oIbq1v
Al5rYFhHp97RrXh6qdRBKnWTjV9eNqYxTYzKET9oCZ1IpJi4xB2IbiI+Tj4FaKqXcwOfwh5CfZ70
UCenNaYNj3VTPX/pkccgmLrBrF3wym0y+jCxGIF5u8J1nu1VXVQ5yMa1d0uL5ycb7bt6PkPeq6s1
09wth6IPaGAL8mcuqRTGc3BVbqN4z1HKPNlpl1oHtM9+RF7MsF7JIyZGOaLFZW1YPq1ym4WYKnl1
xKC+DWV45BhGc9c3+QFpiNaw+t8E13TJHdFHiJDmQQcPahwoEiW+T3+vDlLBKCLufppQgBOl0b87
l/DGKCu2K1YH942ZA/FrEyA0I1vGkP0qBH+1Zkj4ff6SwL4IvfqS0A8CsrAbgWRdWvyu5BD+ClD6
AfXCVCrdO6ZOUgwY7MyEZ0SuPm6lg/PcCYaFC/jjVY9xrqhUiu+CEEwaqH+RDPFsALx9q05+VMN9
zP7BQM+7xcK09s+DI/EZnqLgaC45Es26Q421PMovl/ZOhjnQXGpci1+Ei34QNeV2Wp+kFfTTfNPC
jm9A6UUI4zytaAT4Pwpl5zqOQ06n0LtIFAHhBcvP/PnSpxroFEGqmSHFiQMHkYjvDHIsmA9+jqBM
TB/2FsoDf4zNc+HJp6fw8g910Lq/I/ytotLfYd9rrtPe9dNFYmAtVYh8ivPJu1wb39meFBL6Q5m2
f9dU7ES1Hh3RS+ZKLCvBhTMwKqKHS3UzxnF62O6geCFPAWIlkedr0PrTkIJhH/qaI+XxIxXmvdwz
0ZWXZwqQWLtsfvOS1L9NJm6UCxTIMMiNzITvR8T44+VmQJDr7N3e3IHmIusIF4wl8kbeUY7l7OvC
PINp5fjenYzktHNJU+hBZxqB5F/xEcfj86jiAYGygmdT7rfKTCu0EFUDH88TS6A6ReZwqD52sHnD
9nUpHamhE5R7Y2hGWs3Vhw2P3H6BBn+ncsGBGFM1bkZVab2WBCFLSgNLHcLLES9Y00yfnwFLNhWr
M31FCbo/mdWaCLxz7ZfIJX3Y+/aICv+I9Tzwnr/vF/q7azwTGJ0yJ9dZYpTyoa0HcfzSsDGocOcv
W9CkW/Xe8GuV5npD85rlFY3x1CScofAkTXuCGS7GXDWsCuGo76ego8Y7NxgmUBP01kxrDGZFZn2D
RKUeQcfISrWPComuKpNBl9qjrC93eGZUzLyw/SY3vYKC07XrclUUXMTMIQDsroS/Bj6ynvKtZozu
M7+xk01nYnqiz/UUpPnJlqbb9dzyURLPZ57LhbFqeni5qXL9zy7nlCB4Q2UpAUR0il/3Q25X4Epr
bloozSRLeqgZScOff01Z3WE17xw6m9WlmAaXOOhFC42Sujuep44Vfa7JmN3zNKTJ1TsncHvwHTIg
XKm2lJM++rAdQm5MRhZSV4BUNUhzd9V+183pT8RJ9eLb9d+R8mkZ5gk5qVmvIzoL8KBTogfnBrQp
xVVPR7ABcB93CgmTVTW/2/RKJ/WdtBrwIC6g4+HlXjFzqrxoIpT0foXHFIGOb4ZcpdcajHB65J5p
GnchdNjWdsDkc6vyViqfMJyoqfHdqqfzE26p74Y+CSHvs+Aq4mEUiqM30iVsIFhQusKNOeGc8gZf
+N9mEpH285vs3gvwLqF9eBkCBkLNq8BGDwEmSmS0FdIydF5vHhB8FyKAXgub3Df4damtB438MG32
7fIxSbRziUELzGDdBH41GxR0A/AyBLaHMHJZnoktOgfxDPGBWTqVfYIQv0y+hWQbhlKgq1DxreQW
v9mxoE0VGt9gJbo52F74ec2kWzR667hexL0iOSjSohqIqGJb/pTBxcCgU3q8UyjLWQdxOUetQxTj
HYlClINSJQIriAmncYYUm+oad7IpPDEsdxVeT5kURxGeMxlEFVL4EPM+iptgzF38mVATg5kpWHs4
uxm3oFg33oFaFKyhwjPVqppzZkpia2XNlgeU2fEjIn6EiTflF8c9a1uE4jke6SJaNPJ4/fIbxxWx
j0D4Q4TSMnXhsF30kkLA/CRT7fMr9s0Ha/xKByO7hpEpjAItPzoO7Ki/uYEuVkWM+PD8WdnoBIKW
sJ1yUoB5adg1zYvnaLIp7UQeK9TWWfNCiOjURolvYIEaTXnRMC35cUEbyPUe2HHxg2paKwCMHzZo
pOC0Vm5ELSr0pZZhcUaZk40Z+TNKkf1Utq7H7y/yRpOXHE1T4uUrKbw2nXoMDDri4lE/Y5IoKIok
QdM1qbJV7/uCT2Hm4UC7MiFgetbA+qaL3ztwk0zyjkBfypiha7FVdYIk5T4HyUO9RxOIduauVAxy
QdezcLB9RGTNqQO7nsbq08lhymmS5GjzKRRlqSEzfUGhPeDWYARVsn6WfbKR4OPVl2r438w+W8KN
fowedm3c7Kov9JqVgZ5Zv6B5rTM7iCjpQLkzu06j9j1bHlk526vcwlYjwItc2utZ09PTM4V3iGQT
QBktyeCmabK3vQXmkG2MXG99DAjenUQ/qKWdl2FwAMafaB2ELU7KYBXScSg3J5ra+tQmWN6KCFE9
CAp3NGh5SHW+hX/iV2lHjRsxoZCOt7dc3etHVXwRVOFcp4QxWnb3tef1TLDUfpBR4IcpST1Xjnn5
FRLSqkURVTwWjUdVlwbiwtLV7IDJB7mkIrg5bXjarvoKDmZ+6KwoFdc6WgVOSmkH8C1hV8XsTl1Q
zclH3/jCL8FO/q/QYZPW5jvtKUzuRKNVs030sgLouzJg+jUJkqq3tt2vTcg3RV23MUaUMVcqUwHn
7Quv5JjhejL1KvA+YVR2Q2RiNVf/+sTQXO1lwK7BXmmIIt0nXLMjcr2OOnjEdzf6ALIMwEcKp/tU
Q4M77qQixkoN1afx6PP7TyrNir0bj5Ewh17EdJbKIswKTlqKNDpluWFNShHoHZyijw6SO6eAeGpS
0f+6MJEqRIxzeoLlkVn7HGiyf/gIdQ0OsbzTWho9Yjq3hRQ8kFHwYDOkDEmS8VIqJfyRIDZYXxkt
Azzt2t9LmO3q1TeLJhaR4j7QrjmUBdmXRznimaRGsRVmlWNHI96OGPJHHUyN8077dhzrLRCRFa89
VDtD8KAI8NTJj0THRwwkXFd8tciQaAtgv9Uk+IZZjptaIOwUlW2gCfbrL05aU0IuJXYtdtIYhBSU
uSTF42jyIuiI0KRpCY1XzG4bijt0M8HIQtLlP8MJDwYARLTokboacx/RrhUSM96RwOVkJTXyhjeS
JmJM51JkhboE7JG+vO7QCachWzATYHzzCG9DPUeXEl8Y2JjcBQLJlu8SmWCAZn+vLJcVy5Oq0/Zp
mEYyMXFVn3ad9lhh+LAG09zhb31qEyzfQxQKzbV5xERg5Txj8ZAanURWMkD2im1vcxxV3OyQFYnK
C2g2OxxOpmnF7WJjYLHT3nGB1rc5u2YFihptC8B1YBWln12Ew7JLUm3lQo2DjaX7AjDShqAiPoqe
wzOkDwIBa1YDpGTEb+MIXLe7ZC3IA4U6iWP19fxDPHKMTZlSHDG5S4pJW2hgFy8momOhdJOS7ZDS
iA4drxSamjAu8dPpxqyCaPOsoSoMxcAAEtf0NxfJ5ujNa31X4fmj50B8rY/tNochRR4Yo0ZlsJ5/
1hELwIrw5CWz+YI09skylJUucr1RhHlBiKUUZ4B4hrg47RiY8JFIKEf3Gy7Q3lRUG++BnWDjclZD
WA94XLvuryh+JPh6AdCFW3PpFPdzjg+EMrLqJ32FFWlwtEKODmQ6DUGi3WwA8wL5ZDUYsyPKIBfh
Qhd4bY1mTzFu1oXEgtz3sk2izQMs3RaRQFICWOJVJq/ZcNQYfodwA2W550C9q1otdOWQoCw1+iNd
urzgyS0YSSo002nLtZWqw1NtyVO7JKrlU1Tq6KldoPrpdI8J6f0qXG3LDa5B0HcIJS+kxU0zShyB
tK/3xmX2u/ERxhChzUJ1qCsULzBIbfFo7znJrb+2BoDiPFpZ+23Ab1sAzxWE4NNyHSHzbcV/lwAT
c5oDB4TeCjXkzpZYmGYnuVOoMc+N4eXNXFEwof86l134Gq8J1IHcLQW86gihmtajHBeV1L0vydMq
Di9iqLSMCzTXE5m5lQl2E1tKxTW+KRPmZzFxOLbdwlfcKRm7c5iyhLpJia3EU0RJs/rvRdlNOe+t
qBAOTeQ1fVkWz+6kiaWWI4RTTtevteNGZggL0PLonLbY1ksiMWwxCz0R1YAqBHFA9Gz7wKcbwDlB
fUoS3hlr/Wy96Olpt1aiMl6QG4uvjnBawU1mq1abmOxH31JmMIpJqFdt+SQJLJlfp7ZmAVc0ddHX
GWeb/uACOjMfJMpUa6Us0finGNtpwBmIhfTFWdj/k4lGrWCdA2InP0H1TZn5TnP+DTQFJCf3Cpd2
onyn7/VTzBfGGWOPruuG65lZf6aLIlYqG6c2K6jN1K7PiZ+u7L8b1Z50fvMnEd8LAjE5omZe+ZU6
oVRcvmRL9J2WRsFMnqy7lgUsqeiC27D5F9D7NSPzCl9mlvbsOB/UXwSAHKb4C+AhV9CtU/mYuTpW
V+LcKkAfa0cG4HHbK9pDQXXb/4XulXWDUKa71irDg4Rs+DoNspX9oonEqGaWXclJV4z903TEKdtA
KeNtrv4DvPUQ9mjKzOGv989QuRAcF+2jXNMQXsREwUf0roocufWTTQc+NdaYVaywwbIWgTRvzvSs
PiFq1ABZQkThbBplmvyb2NAaWci+GGmZ3niCfgPuEJSG7xtyDCMivhrK4Bz8MSjHawpvbTiy4z6P
D0jtMJ8q5LgcY3eldohAHe1kRYuH7VbOa7l5FoP/frJgai3uz7dDozGy8axTvRn9LoySjXOgfl/Z
bg6iuG4liqqQIn5zoQVIqTARTIhzcLGvVrqzjqAognzm0zGg/l1AMczGeM4jQ3hKJbbc0W9KtL44
fffD4xJxY0A/s241lraQLC9Mix+T1y5i+BDb1EXrhfYTy16F/F6Q4aCMv4RcBWxqPK7QWMfTsV7L
QXrC/z/u3g2zxMAcB3fpNaPkBf2iSs5x2XSwm4U+EtSp9dfhIGiqlpKjyX6AT4lgnxM9eBK3DF/l
DbKwg8CkD5z80kF9uLawbU7BGL3BIIxmK+GK/wxF0LTqDaupp1D5aiw6yCOQpjdqVXQc2lwlriDh
l1PDCw64CAu52T8UDHirdJrmGUzqkmS0WSeBOZoxzyuqzSSWC3ES4LrfODn22Lzptx2hqTmUZrdN
YQ6sFj6dFMU+Quh4TunbFSmx6fVAIO2mq3X5OKQKLaYtZ+kyz+RXP43rg8nAXVNkvJ8jbPGSgfrh
gChFUqfRE0Mg2LlCkQ0gKtYSu4Z+lG/fcu8hRFyRIoog2Feb08xc3icPcTxyR5BDUzOQsz+GJx8u
c5aPvKhr5W70zDJohB70ueQFNvELeApJpbyWXYA0SX6XraSEBFgLq26beeEoRKyXKkBcCJljfzxb
TLB89sPVKQemG6ngisIWFNzifxTyC/vqAGab0CmoVN096ZfqICnZXw/Q/UW+PCxnAwrx20MZ9wQr
inS3b+aOmHhpzyb7F5TZ0NBnlRCnwuislE2RMHiIcNN9CCPnEN5z4ivIfxPMEVHJfAXSh1XVHsBN
43JJT9kASHIJHRcWVQet3Rpl9MBKygTfKdDQGzxqCk7oFsiH+aVdthst8om4kS7b7MK8RhWmGAqh
CBpQX/pEKhHhyrcVNnvxfxkG0iKx/euacVQGfaf6DTY3L6AcwJGwGVasTebX/iFfT1zlnmIRfzvM
cJ6PxgzW+4gxxM7SLUu+Ul4gGDwJ/rxqVOapq0lg69NmIvPEY6nIizWxqWmmYwxPsSNu3n8UGghM
k52GNAP9DQSkxI3HRdL7bZ+19JmGLfgu0ltzdDPvmHNkI10gH+T7oKZo1l+T+bInrkSsvm/c2ogE
eK3OVNBGOEOrD4y86iRw77Zxqi/mhsem+1Gu3OaxWaHDxn3qmG5mKBYFbNBuuC2JfbbbPOSAIMzC
pxJiLwKqeeMcnXSFsCcG5qr+L9aXHaH8Wr0f9KCtu98uXHWkceXvbbuGCGpf5YnC9WVQys6H8899
uoP2R18tIf8wHnE+y6btnsfeELEvtrEEVdykoiczoCzrvhQP5tNkSVQNRcjpfdcryA5zbPbrnFHz
niev4Joo03CYJLEkDm0SCFUKxOGMrJMs3aCOCNedHd+O5G9sAY7+kZcShHyOhd4H6NpUu9MABu/N
83J0SdB6wbULLRsypPSc4KOnzqvhy4/Cc7rePON4dtaRgbd9uhmtUVu6llYA2fQvb9Nj2KfP3RTE
ky+gMa0HUy9zl9qg5d8KKOqOG2jwgDADEB3+Q08towlWg15qgmzSWDnXIkR3aMb3yXTksjgBLF+A
SfJsq0niE+Lc1eb7WZpK9w8vhkBfrO9fAkvvJSB66DoxGSLWRTO/sHOB8h9/osPZFPwqEa7Zmzx2
gyJIvOQfsO14rYT/zRoi2FO6AZeRqUG64kVv8Ujnti9+fKZEvAgPQ/h2Q1bVTaEyMIpNrkZCno8C
RkHwIyXozXqyX/K2UJLUsJagSK1E3w3dmhQYWTO0E0ZMYzVMrAquEd7AZZVtj7HrFTmjJaoFr5oZ
Ran6e3iOz8nvT4qcLpzFIScVAIoo/U21EVc7DJeKPwuJa/R2PAXLKatiImMRcn3JqCmZy31c0qqn
aupAae7regZ0iggi21hpt1pq50bIeLvRvn/3FdOTaK6dvKSmwmYb6+uV0tyPDuF8+/w8jgliqSVQ
QlP+djaAbGJuvgQYZ3EHWsGE2L5YLNGgsvPzvMWqog77YvlJV1QLv5PYnHNFVYXG/tdK8onQDcnC
xbkHN4Y0rM0hFxPUpWxFBJwgmzvoNpcmk0eBP+8uVjH8Evqx+mPXeom/Vn0LO2Fhl45JyUwkshIy
yyPTiDfFVgtM3Wp9cJ7k6IblCrh72a5WLpEkO1+TDQMnJpbgdIKWEcjd8SF2cn9LgMme7TMViuDB
y/G2nJlrYhLODQIBsKb+TyMpWQJEdwMfw531d4kezZbNp2Gn6651paKUohF+/bH/mXE1QdlOerRN
81npumAhoN3Yx95fOB2R85MrGOUPekIM8zLyGIrEBwWOvERqaBNU+XLrz0d5BJZWbJegUw/I0Kal
2wrpOvzXE4I9OpDkcujngNHo4t8XnHfjOPkviPv/+MSK6qpLmYlK3XGQGFCQXgdZa8C6rYacGE8n
RaEgEvKV31FGCtEa7gkGKwzGAMo88dT+u9qpg6647opu04LxG9aAgOxjFzk1qgvXRjKezGsyizwO
KOI3f9JqSQzjysrO43isN8AbIgymRBaz6l2iiQZSlzzFeRQBT72t+Cp2wAF9tuDyrysfoSreHAYs
cLXBoFT4SGlI4dSDI9kfD7F/9GzeN8wsIIEnID2qy9eXlPxo3vZoRMhQmRNRor/M+ws3NK+TlMvT
lf0oeEFrp6eA0vxSn0q3U93br5yMUpzVEvBQPb1YznmBjqn6NnZ1JCdDh5cfDqT2TVRtM1zWbQre
leG7E+YZznA58BSfZTwv+YJ17Q8Zed5wWFYz9xI1E5j+I6bknj0k2rM7qaxJyOJ89wkKTJv2Nnel
QJwgJ0wYCyWUEmtrhtHDlsgNaAq7AXnmATxMe/X/C1TQ0UjxaAgn/+fAENXMkuSSptBkyrohoryq
9PNiephyTjflA08yO4D9UAvsw2ak6e49BvPU4v4ZB9Xt0/3TMjw1w63oVCp8whg0trPYcnHRM3gU
VgT0kDr/GbHUK9wX3wOgDVhvym0UeppC8d/zIcbKquhKp4s9xfaU5ne11Ny0it9ArygJ0z53U6Ch
BqxhzDZhQACYUv5F3LlHE6KqasNgeW00lbablRl7+mBYyqnalchJbPDPgFboG5KmzcSWWHpkxNVV
Xs43GtRrUO9HaLpGLufBOZlypj+QOFeybUVpMixpkM6RcNzhlu1YnJJwWtgJ+Kf7ZHECAHCnG5pK
lNLXtejmDF+zeAiK0Q1TxTwKvyEayBrUWEG53Q6Obbz3aE3sYzsWZubTdqhdax0cSQ7mEN672RtG
LXB4PZ491EDUYu4ceXSKqo4awkONaEo8/wlydRP6TsK4b8j0JbssgXaYHPZAzWjLZbSHyrBJj3Zw
KHreRWyDvs0AmQ9UJ7QM9Z0hf3+RRhpRShETs083YNiz+a4Uma1S7dPjsQrXHwmI7dEoRWT2J0aR
iI1cz6pYAA4dStINwq/hv5vr0OOiLIWVAfodrtaHY5tMnYChOz/LAd61m1ezLV1ERW0z/8Lrj6Z0
JTp8dOEWDpvMNhLm7LViT1+kcKcLateJflUCdsuP/ZTT8eSSXrwM/Vt3oITU6AFHlIg1tfrzAgWq
6t4/tCNWvNSow5RHz0GhArrEQ2XQefAhGJGTaYrs7A0/x26axA5jGoaBBf6ao4GsyqUjw8Mr3eGk
9bOc0PDoR77ZVG3OlVCnW5Yh6mlA5kUuxLtCtjka3jwcmoc7C9fYH1NuNRHWk5kfSM2PvKzWRXIy
U2Naswj/EG++9gLllgc1X+Njzhyw3ccBKo39BwiknH/lOCNpNfILwGbXnJQlYfSqPwvTtXzZcOtt
HzSq2CQh0H/dRwOLRuXsax9eI+VhDdLhAKNFFMMsz8RB1QSku+qku9YcrVw0EPDmhCQFibMtvr/m
WKbpM4GdFWyJAgwzT+VhsUOXjDt8gOGe30l5S2S8teClz7gGJjHzKkQqAXL/6lfilN7gzouqLr3Z
7gg437p3U3097zdm+K5I1NfeqwS1ei50lRqXc3+h/Xg8veMvUR4eHGUOkGdLu6CfglXyiZsu5g/W
lgcqbGTzNv9xqfB3w8tOd+kfz6bpWbPlVb7p+P2kOZc6hAP56ttJ1f5ztmLwy1Gp6rXaWhgkyUKC
R3M5ca15ADtRJ6aQLXoxcffk8yEzHJiSi9qGyUJH92vnNlvfE5yUcrwJory8LYu5F7mZJttlxzid
M/dlUjDhO1NJvv56VutbuxNhoiHw+Zs9quFHlWZJ8VFu2wiCBY/9CeSMa2vnKO2EX8eC7DSy+wzf
QmKanyCcWy6A/b4eiO9kYwtEEqH43KT/5Pcf9rRgOtYeoUTbM72A66s2J2MKsSrw6DFDjnXWagKG
zmh+HQXFUt7fDq10hIPfIySjIQNZOpzP4W2bpWo97g6jq0Z/X0BwE1AwTmYtroBOdiX8pg+Nwxeo
OykibG1AQJEfEdSxbE7/mbvrtcAvodK0Enp/HoFFIroBRhKQoDJy32jUSp2T5JnIyktsnbcEcdqw
D7ssvOkOaT9J7xZ0xU75hvudaeFAgiO+zeSF51GqlcfJz3ZIyxtwKMjr4lk/AWwIgpSrDWKKiCFu
adnoYVX8zLdMi/koeyffCfhkQdiovwNF7qGcmcGl3l5en/Gff+ICe37aUISe8LUUYZvMnje6bwpm
gXgPm34OMVVwfUDy/Vo4twAQAzv5DcEDhVLzBCBprGeVZ3RwKAqWsb/6Bx/jn66cUFWaKKKskM0y
h+ov8ORLrqzI+fEkH8aF95NW6Db1VEFIUwh6Qjlshvels/8u0eYEqarmEzDmsh3GLs83244L2Lqn
MtEN6y6w1TufthsS0557OIgHzvNPCm7Fdknox/IuvhyN6QG+f/PJICwd4Z5lR+lZKiiM3lSacfGP
xS8CJoVy0ETYusbXqIZB8xi0BA0wAYt4WAS2sfhlaPahAogvUcjzhE37vwvK4GOVMb5N7VOqizCT
vZgz2fRDrbTt9qWOqlylTeJTOlD4QM2oboXxHt3jtmg6L/lwUsCAp+3kQMiS5A1Q6MGibYOQcsoy
Njfuk5hjCKma7eGu7U0PJboS/NWRBRsLDftOvphJgeOmCqxuCZSGw3EzWI12RqXMih30x1pbclp6
u5pDm+gDAnvAT+0AxuM7gbzsrTby5kfHGUDkqVhg2uHN5UiZHbJH+WtGQC4v8nIZYS9unme5s9Gn
Dl6YEIPQV9j8HkBHYN5R40c2LLKJ/jd5B07uy38FbhjE4IrdwANODnEbLUiFwMWVYNcIS3hAgR9B
OIHH0boeGGH2ANiTFJao5yzfPqC3QeRyks5Ogq2ENSKS4SOQYNqR8N08631n4zGQMAUZnEPiF76E
pFiVqoSCAg7WaqKP2SowH/kzVT9jf8nW6J2ep1h9EKXJ0vhS7kf/6u+ytzjIG2XwCe7f2rNPt4Za
J6dapLG7zG2/GxyuIv6nNgqazFZgZswniMey1SrDfLs1/9psaijlv5Bm8RLMchygFxW6qYaU8Q0Z
JDYK+69T5elnGIAwaspLsRXAbXTZAk9t6pR4Xrb2fLSuh2X0K0jq2ThLPUkXwDVEHsSXhv5k9Qsq
M3gCrliv6N+vt6qcXNayJBFKag9qQfm/o1H4Z8eadqjSDG5Dek7I0pCqcjC71RXFr656ofxpdLKc
/wTUhMrQRT/zzr31qwfJcAB77iDiJd5sUyCReLT4mVFqqqdB56g60boUAzgELKGvXYZWZUjm3kCe
ZJBNa2kcPaoxd8YrplNMxhvBiTp9LTnYDHoNb54jXOiIoRmTHagwDVSxYKu0pTmadYloU8mf4HK+
VvgVz9eWds1j3s1h+d0fbJDjtpPxW8XcN0H9dTIelpNXHOn5tJawn0JVyh2s0mjRCiApEvVuSObd
28BurQwsLf97HtbLKnAc80+wzFVv+t4v6VAqsfwb+7AYDby3EYx3MWhODeGUrPPzOcKdqB7iqElR
LpBuQV3tQPTeOiU5SLeeG6PyayOQUNGW1lYdcvfAlWeWTiy8b/aElzraU3t9h05eZglY+kV0TPmR
7gtHsC2ru04A3a3GCHbG/WlEv+VV88P6IZ10R5DX+2LACKyPSn0kHsqpb/8hbhEbxyfy1C871YtW
z7lY5zQT4DFgnwtlAp9g1DwnZXaiaSX3czg3PzzRerpvu0KZtcYUxvHLqkPYX1f4MaPkUcxpatxe
sk6DN/Q2Xi6V9u2suOTq+jflUlQjzCV6ZCpprV31byjbaKiMV1vcG25xSFcLMoMnxpebN/YQ5YsS
KHl3wY1khm229ptw/ZSJ0dnXbIUaE5A8qe2cOQ+FPxB9fv49K+AFhm++GbmRvSs7c/deEjMSnrnu
Xgu9LPXcSRjAYg5Pay3Q5PbeKuYlQxdw0uO8IHGjWQDzMCY3qhZy0nGAkhGbxDuz9b5kSJm7oESC
mu7FbcqSfmVDCOLxS/oOdVQ88vkM9/vdrpAh5aPd/QavVRkc4o8+cn0SUIva+7ASAwlP34EZPFCO
VnEiVC+q4qeC92KrAH67fYLoglgDcO9WlM2A54xmPhGpsb8hh2Z3lDnPHCzqruDDRnoOUDcnFxKB
bj05KR61IABxaP+IUAmnC5+v2F2d6p7eT+1ONx4QIT5cEAWv5VRAFh7i9S143QOKdgePl7au5E2i
/WYKUmN7DswVg9y8cs54brLCLztxJcqgLenCk7+jLoKtKDLzzqjWkg9Wlxxh7m5EsZGUz/Gf5omf
4A5WL/xYQuIEskqPuSYznkd27vFM/j239NGbu6MEthNeXbXTmbDSjPSmoFYqzYRrrCj1KNYANWvU
WUqyKcR0zpfoj1MWL/lKu7RW2H1YF2LRumZctpwfNOZCw5JNUzoBlBDE+CSqKBOfeHjYPvJU9WP4
GEHJNPAzZMxCfNJp7KYINISKTZTiH7iNhZlxuX2R5GUPVMvZ/cNf0IC2oRxAsn8ey8q16WzzUL47
oj1JXr692tY/b1bDfMX2F7cZODRXnduzrkyUD1nEBSM7rI7XH6FA4EIABwiAa2Dj/xaP4uXDEDqX
ZTxsTWlcDJKn1iQCJW571a7jFiDwtbeVN9PargWSafcnj2R1nU7sUZf10hqk86Sc0WpaqdoTi+BP
E4rrmnRxhLXWKD1MPeBESw7rFBTJp+mAZwb4baLuD2BahgEEmRkF8ketil4L1btYUVG6W3vRnWXb
Y4pTWaQEGPyjbIlmP4xQMVJ0yReVxwCJvGQix3d/tdf66dqFoxcvbxPdkixwo6tqaO8ebxlvxui2
mhh1BesNy2zKlP0n51K+RIQR7HGmeFKUn6K8bpTk0exM7uODo+1hKiTx/4PL0JozO8HYBxIeYXb9
92btAZKMX0KUI6IjhPZ8dkAJvC/nECxZgOlOkLgE9dcFiQ/zgt74+cf56EvbhIVKpvuB09U3pM+P
KUpMG2gKi0RsFYnWZlB9Z238333H+37EOZb4b8sztO0A40RahHd8qnVHa79AJQc57nB/i0h2R6kV
TbSFyeXJYGj9gkDpmhz0nPCpGX7bn9khpkfD8WqK11iJ2kOZyysZVm5RpXMuht3ZovYLR2ZJPZOg
JoA39YkWCt9a+VfGnIfe4zBUDBUBxiQNFkJBk1vfvzTFdJQrDnpy0rMajYxeqNYyVM0mqBXMKjPY
jeo7ES+0ghVvaSYESxOLV6qu9UsVpceAXO/VI6pzDnwvgCWE+o3ewdaJVEp/z1KutceytQ+hW0Gn
u7k1UwBgY1XyhfQZR/7nMIQGy1mS3z7gjvqh6/4hmuFGa+bb4CsODKzv8kByVtYqnzycvfrrCNnd
ygKKYrCpdPJQg9kEW8iEChjDmYomGbIeZiOqKYDC3aZOFY2hRna+Nu1M2DzbDNdCbsKgcJgeSEpW
QPc79mGxEWwJfDU2y3LfeJOqV4jxXIf4HFFoY6gUOv4I/shb2t1x1aPbS0LQhKNfCiARBEO3oTsW
ZrBzP6yagZeLzu1hGfQ29VB+xE0i5kpJIMhZrrVrJ/OzYcd+Eg0CwG2dTU6+m/21WjFMrZb2FwJt
4/y8FnO7EPfFcyc8ETLzQHKXo7FiFV0DrlxTeOHehqgJmv48WG234WpfvuFR5//28JxWysIHbWrP
aeO6BruVCvMLVHWimuxOsxe0aiECBzI0qE9xQjNsz7j2wl0am51S7A5HFPYWSfG23PmddBtSHDkm
A+JJmukkYsgnWr5VrfL/Zalp4vaLfJpOj/42XzT9e4Wh4PiYUuoStqO0swHOnHJVdG9hvzuI3kme
2zvArQ3tXXogSzI+2Usd1BFk9gW6SxqI6K7qjLOrO1LHpJ8bZAIUGyoAQNOJXCv5KowOHqQPmUbV
S+zBdVapyZuwRf8h1rz+v2vDY9uVSudW9/VIDR3XVf5L0BnE7Cpsz1KN9zb18tRQcsfx9l9jpyhD
99LjLa7SEohcIGZ8w/68lV1BU6ZG0Kk3upHlXpJ2ZMRp07oaeXFh5+LmJsB1Vvxx35kBApjevcu0
q1GklalR5+vtTR8C62o2h++fv89GjhMPDPOXCknYMfBkPZNbMx552jaq/EnGuY9Z6amKuj4Wosz8
ilQVejwh+MXsSUlKIVWT6RLx8OmPzq/wkKnCfOfNDfwJRNflhfrObrVD3QUZut0yD7gnDsN+3BUg
FyumO64d5pjioKyCjIX8Fmr+kL5+WG13sHCsVlkcaqyrtsISJvm1riGhjSWdvLaCz8CdZqndnw2u
j7Z9geQccQfEeGVGHWYGEIT5s8XW3mH4ba9KuqgO/UxtSdzUyviAmmPTnLAuPWFQqRGe1m9gFHx8
R0tJZdmDzwlkxndUrT77L91fZuOqfkd4xLW8xfEoGmJ1+8Cra74FMP59PZWYAkCiKHiRflIIaWhv
aSzrQP+dzizvrfUINlVmg2NNib+y5NjGOFcD/wZGXrQggGb3MLOepZtQJtiHhcm090JQ8R2zWYt1
OtpEM4+DiC1N26mvLto5tGSweUy3mvWoXRE8o1YT4KDeKSORNYikIyU81miuu18tSvwaBXtQyo43
KPIoJTXgEcR86TWl+euhevBLEID57T9vb3kfBGhwLqLTz0Yt+4wwMNTmvnrCbpJnKfii2Sbi+ui6
5HErX17k0FlNAHGVs6Qkrz9tuh8UTkJ6qzzCmcVw/NZzqxRjAUW8dCP1Ve9VAeECZF8x/s0JCLku
T4csuSu7KvcCX88ReNguIAZX759TayfUUy73B/2kMCepGVMUqT8Use9yUtc6yXZUhD5kEalOEttr
5M6vGiPU5f4VmbEHDnzGo7zxjemhtJqXtaXq1oJfdxhseeee2Qq9hwY2L0UOhMMvXq1NBT7dPBX5
0PXtcDVg3/VGZ3DA2Hg3eCykgi6tKIHVZx8A7h7Y+wNMoSaaAxjjwCJ2pnxedMWZNybntKT+PHyS
bp51rk3ZmDh4S2NSRdwQEK42IcxDcm8itzmepQj+qeIAoRbdeWdKcxNwSVaXOv8a5txh1uhZ3zdU
DkloRCe6a/lt/zbfaJkxHZu2P+KNfUDZ4gprBBwoS2y/hyB9hl2qd4aa1JWBo31ZX7uRMgM5Z393
7G/yhwsEnSSUk0Hj9d+BzOhR9zZkQuQNJujJ2Hus7en9aMs/YjTM/wEP96CS/mb84h1T4wG4GJFE
PZgCjMxUGQvhsIdg9QMmjAIysnI4vC1KktoGsblIcFz4Y3CvMtW/1awgiiYil4nq6hOQbtNJiqgY
k6ffPIMpZ2zhm251cRtW2Cc9rcj6wPkQzxOiEPhPOehkWX1ado13PDwYLhbbK7dqkFGDuTrOb+p4
TyuXZ3wAJLeHb54Z/arifnGT8vJ2Tpg2YXbESyzuGWYh3Mx0xOOy63fm5HDyjJbpTkPzCsQBbDNY
9YDCb1tY9pevQkV0So+qRLLb2TcsOqWQA6qes1CvPFachyv0pLZEQCgVBfsEL/Rc8Cr6ZUY9FZiX
51rfnGzitlknX4pxJCLR7fNzcLviy4eMiy6RP4a64Uux6GwN6eNALCcQH0vBTZHPRQZAF8uxZOtp
y6nR5OeP53rViOBx2he06yBQW+Yb2urIErlaixK8dqmHne27ZQ0//Q1c3j4plj8bp+UOk6Ffr2eL
BVfl4itjz6lYohumSAcEdZYaDSM3Oy2LQwINPOMj7o6ITaVABLreA9UpumiwvrCkEj0ou4xa4DLD
ud/2VktxWIgBVc1/0ZJRrh8P5Vz8jkWd8pidfLThB7e5zT3Jl7u1OWRmqf75KP8kA1K/4y6p9sL2
yBwltdZp3b12nw0fM81uzLgFGC7jVh8s/76RjPCdIuW7vnn4wL6IsPPK6/mWENP1EYUh/oe65/5M
VszJfgJ6lZLivdTFvzzT01mRmV8xXQBRP//W8c07tTMGHN+8F5cVpviL9F5vb+UV5S1r8GKTv/NH
DX9yjigCH2w4NxMmn6hu27ICI/ujuMLqclPGuDHP+DbIeM2SPAfW0JVp0IsZ1yj1YfdiiqFA5s1f
YT1mCYUqH0Ka9ewByRphIiXOY4sTfgWVzCGRnUhXj73sXtX1iJiNAbLUZ1KA3+rhDviKhJvU5E3U
+FMXCYjFNyn4Nrni2ijjK6x88g2B9CtNoPZ+XJY13c3rb7dIJlLPUv5GgwzII/eFk/4wp3WhJo6h
lyWuDcqsSd7WPq+tvWkTfXDfh58fLYRVGAbsUvDA7knm/Gfzt0D8XYxdixappSJRkjBErYIXPvwZ
uRuZTvrY97dujwt/hKZqizQhWtmtScSRlmc8uus6z6uEGLKOe1LEDAqPPw84a/jphCVr5lT1XV52
ePuZf9IKs3ZbarDTYlo6zVtOFjAPaC2bygTcqZctYfuEkNoVCL2jmSQtfee4y2tYcyrBkDOvGKyL
9K9HqkyfcOCTflVW8hxcPNm8WLXMnllfzT15g8+4/pNfQvsfaKIgaekq869scKpPtP06Poehvg/x
E6nLLrxHWomK98QdJ8Ue/p3tUu+l/p0Ep6JNmBY2ORk99M/htIT9e/ZOX7G9N8sP6N8U0YHwffYp
zg5+mBjSo4hj8Vc6Sz8P+Pehz94DgivfA6JEl2h0zP43IpYN80FyaHDL7G/ES+GuzcMRnmUICsxH
FeYHwSTxabdylMo9H1epZKKKHBq4ujnStCEHOjG7D2D6LhoS9JhdI1YyrVwpdM/a9tz2uXPQ5pbQ
UDYS63p78SyZtERyx1UvPwHrG0zT9fwMWRtJnMw0AkNuHidlmOMRRAUW47zOixOMgyijcNO7xQNY
jJp6NrVwC89nLd3pZjE3TakyMqCt7i+sVysLU6KbOGyWaT+moG3OHGwfI04oYZmgVG9StZiCi0gQ
mHyidHeAGsz9eBZd2Qc0WZ8Mw6cfINjgVSJaosBgZ3HQHqYjttmWhjAOntOUlUMYNy9XjrVMfeSN
z3b0MaOsl7qL2wW5I6UpYJ9b+x1V0HihXh+5PfUaNI6BOrn3tAU64B2Zp7wzHj/X35rkVrEQdB5h
lgGj3UCEWmXV9JnvnwTWCWIdPSfx1cQstrQ8AD+yijWcFHnXj/4TSuOAZGk0d1ZyFxic/DFH5GdQ
Fk6sMRTjkexc6otWf8Zn/biWetDTVSR+DzGQsbyAaUlPUTqDHQHmF4U3hbfqC1PH8bQW2v03TOiJ
E18032f8KdiUzrAhdjpuJ9Nwd1VsFHZrPN7bH4K1aA92JSeYimO6YDO2wX+0YyfTM0rFMqx+uknm
kUUM5EEWmihpcEXWTrRsa/aqxlHJIla1Z18NwyO6GRLfzZ73I4vvFGUusTIR5mQuV2YmqLzemEeO
c/w7CUhCpJeN32sh3yiSo6dG5JGp17ZI6xWMhmfHr2Rp3Qt60+WPeHg7CsK9EwcXmuxYANrtjwxS
EDciterZiin8P474qRSAkSyBP1Ae/L3YpGgXPzglmVPQtNyUb8xYU+K2o/1FOR+29jxoHw7N3RvG
oef1Zcc7D2twaS5Swqh1Gdz1ieFQiYttleM12doewR8pX8wEPleIwxWsl8V5FjLE/Jk0ym4N4Ck/
FzCEUcFRHkLQpVu2dYmYkFhaOdiE07adxLNVYMOL3oHJl2i4iE/jwq7Du0/gQUs2ihNTACKrsNyF
ZJYP/D+lEF2SzA3JtyCHvyETep2cV1tmPaWlqTzo+XXxU1CySYTbOy+4HtfNT/lBUmTt8HpiXBNZ
RhEHEYDDNdHvArTcPwJK1kQKJn3sAULvaTbtyqOXnuvR4RJcpPi5Za9r/ZuM8vV4dnyBKXz/PG2W
s9IDB/hrS2aauj2aE7A4dLBBD79sHYrLALjyIQhLyBES7qW81IK9tRKzfhEJT527Pgh4iL41BWh3
nb9ilIemeGVuogcdQTt6gSFPEhXnBAB2P/e2heURy5MWNbNwnhEYda/wCSxJ7yI3bLt1kMi+NywT
ns+F4606Aw+/uSb3ZT8ki7HJzfHqryEoVue3MX/pqHOWWJj6cXdUwRt8BO+Xw3t0oHqpln3MF7Xo
rFqzlUkUhyz1oLV1yMbygniUZDEffMHYswcTEzf25YpHEvTUE4xPV0g6yIqMh/HnbSbScW7l1paQ
74xdZWDwG7+S6j3diwR+l9Dt6Ku5qbIe0C/FR4nTGQGVb+Wz/2dnod2Ks4NpPYCFYvD9Cvfn5BJY
tKGjJZGgRbCqBxYIZq/BIWHW+t2+JhhCvn8Pe6xcilOKue22TZUWLAXIZayMnkkxXZvoWZ52/+0n
qcmAuXOJkhFlfGybw54jm3Wrvl0qtPSj2FgBPnk3y9M26cZS3ijAcze2cPEQ6cUEFfWyjnmx+8Lf
0ZhXxOzGomoZlohJx4nhayw/6ssgIrRYb1J4E/GpynqKnOg99L5YEw1eICmAdSYbxbnZgXvFhcvk
HWR225TWgCLnXyudphlKQsqRJY6SyqunrvlvWhSLrgu4BCwlx94u2JH1llqkafwgvfdz8/RwNhib
7cm+fUoa4sEUzFazwyWXqVbIEq/udecTpiVgkrtihnN5jpsEQueBGEk3O2W5U5lwl5vi4v8M9/rF
H8AcWcuQFN0WiNaVbOotJzkV+mtXgIujodyZDDppSEe/UiNpC2b+XR5OFRxyXAnieSNADc8jIduy
TY9xUe3syZKoqOJ7Jl+hNMrvNH6Kfh2anVUdTWgHdkIxud19KYKNvvl7h3JlH8Www7aTtg874nFe
8ZSxJMt341mQVfgfmkqSjmMXZ2DIqMD6CGtZCATAhuD/0iK+VdTCL6TfUMmEl9E7SrzCqKU4eTLb
wFBPDnZDsawTxc5iWf8oPN5I7InSLODQyo4ovnVj3tfMyRN3XPwwEH4RSMucEyvBYMvvSTnvi8zp
95t9r0JMLnGvSCGbvmOaAvg1ZTetDW2bNen8Rot33LhDHob3NeRtAQdCxdNejH9Id1dbCNaUvzzQ
AyyJFgcL6h2gQuufu7uOLJ/fp7/1MUgPUscNkB/5OjeenoqN1YYG4cl+eYc0QWDSHoFy4N92niFY
yaiVgs+ZjIsKY0rtJenU76EGgGsRlxGFHKeiVztX0RFtyYTX+pss8oEfFC/UQH2n7wqaZAxcZits
nbUieLzkE2qCYa16FSDUckPO0lT4BXjpZuVquhVUV2v9G1r8kcdzJm27Kf5i79Yt59lx1iOPYeAh
4Rh9jIuTlI8JYWO3dnwzb7p0pJmIUHldOow4jIuCVHIkUJuMf25o6VEkw0VjasjMX6a/Vpqi1W/U
BtwBhRy6PzdF0UH2M61WTtTU/QLEWwDH82mCXIc2t/xDgU1YJzk7G+XaRn+/o59c+5Moy4DAeXnZ
miqnP05d9NEXUe124WVOIxIrgDaaDpzpsyMKHl+8HUqNe/glnvrcSMOi4Rc1A8xFP1kqvjE+P7Cn
yMltAOUdnfvGh3s6d+Obo1fNwyTykZ4vZy8tlA60Ti66SEhJ22C40BvRoJLs5eBaTdLUkavaz82u
bjoTXNS3bcBgBVyGy3xf5C8ScQj58cMiRpgCdhTRGP9W6SjJtHwGnho4Whjt+QZ0t8TZ+rYQX88N
ua62PSGECofOvD5bPzThcdLPU4ulfxIUyExF8omIAu2TimUcVXLXiSsm7cGym6qJK1Grih/FZdzI
eKqAyDF4qJahAg3cP085803OlZNtSutZtrVrCC/GV5waHzQdnQBo/s2JIKsdaIXB3ZGD6U3aT3lV
G6WtYlVc9rnfWdHMHD6Iaadr+edN69kizO2kkcpqJ6IxKICYmemvbiqGDbquK1J2zv24pF+45Bvh
AOOePjTBolB6kIWe2gehQnxRNoH20TZgyImh9GA0NEvGqODc3MlhOcZ+7LRQTFvUaSoBCpm7R3WO
dZDADXiAFxpJbP3SPGU1fPhAIF1/XMh3hTz4Kfw3lsrMPbfiR5Ru9DEwyp8TXYMMIfBJDyRi+2kg
a9DMKCyKiGa+TqUuCNHkf4b3VHPvDb9t7IQiIS3Inljn0/6b4dxjmCgNdODwkRoc8D3/YjgwtY1w
IRr1AAppuadubbrdRSVqzvNay86F3qaAHaeuWzRRc+IrqkxI7UEenRmMznCbnGRnCZf0E8fmWZCC
LbQPS5nk61kTces4vTSYZxoQX5l9vnwRO/EuQTVapdRNn/V3TxS7ENLn3BfxP4WRX5YFkzbP74hf
264PgHd2oxHOmPBP8wa/evYvwKTQQPdaePOcpBQ1tUdMoY1UR0YtoGAVMfE7sUD22Jbwd2o9f/rV
ZtRxkJI86HO4/iuZrvpUtN+RyL/u0a52uDyKEWtgAkTTJNnnVCOaCzGHsTvvTxghBlwZ7puOmkgA
NLQjb9AQCHAc/kt78KExv+bK2pYcoaxalmDGFEiNCihuwbl0QRK1m82vatUzFVEu3jcNYMxCUmmJ
KeMC0u/b9SYFIjM0wJxMkHrcHw/GLaSTsUXpbiehiovqG+Ut1ppjVFjIBQLq7G5cUddIX7Z84mtV
1SRjQJEcD0FzTBegp69YYwWx+KbI4YFuOh9CkS2KkF5iS7ESpl+ELPF9Ru2+TnhLyKhbF4H+bl28
E5ffCOir+I7smrkxa7734CxWMsCGRQDLtKGaCGf/DhH8GYi7cjulv15bSQW93qHDrk9TNtIKmkqg
2zWAuJ8Ni/kYsXqVpIAdEG9fycLBd/ECOjUQOfxZY+msygEgRWLdKoJoQ/lFGUC6VsRMM9JG5xmN
hoB14IdBZBZ8eP51AZzlAmvE4pPqDLb61dp5uFa/ludplLFAwbCj056GflGt+JiTila1/q8bhUbl
znaeBQATggr5qyD5gbiaJaTzmsijTiiNhzPLnggyltj6BdWdRxmgOkRxm82gHPqQUwn3w+DXBhIj
pJOSHeaXFg9eq2hXO5FaGAkO9nB3Qo16Xe07bM/iSvF6LmYIp9OzQmHddqrOKJcBXdZ9t/exA0d/
R71JdKTZQB+813+mrRLAnrMROmuY0XemRuwCkfcXbc7brSjaviVm0coOwLWQIxdYX8MWJhpBmfm+
uM3IhtH2wNIrVAoTWn/64ReXNyWaQngVZKdhrlHTDeguuEUFDCE6zWLQm/0r5HmntbfQl11q68Bb
XH8wk8MNvzLH8D6LZJf0twkFP2wJQUd36/+ta3l8jCZN/LwbvKYkc+7L6yAScvP7UJ/LdB52DxoR
TuI2/PQaKjSgwzgWiEGCqB7v/PQNIHB02cbY/CA9FsOePPxLa3yclQF3RjVkObOp0k8/g6QsMkWI
A/bOpeMfsr2T7RmvscJcnDd0vh2vKo+ArJU/2qvLZunLErylxdULZOKOtXBahYm0yRqQuy13DBnZ
VN6kFrpAVmiCbl4xvJBsknLy+cZ+c6GsxRLD5UBpgWbEhg1mpPx9QDQhtd5iun5JhAxZbNQEG8ay
BHsrpL+JTxKvPBor8iZ9C7uGV02rNLZEnEp+CsATy5QkKIUO72YewTR+ZAVA8lf7Mq6+yP1G+3ks
MWEU93qAdgorrNaQI4dSoW4300iDF4wmIwn/6xqQ0nRfZfvDHOBjqAmuvsoOgLV/+orUgxIi5f9G
Q2Xfz2W/4kY6Ts3HxxLxaO/O+8oYJxYPOkGGPWDW0vkFUAvGtLmOspthpnpGBz/cRfIaTBCg/RSv
UMRZtEwzB+pnm0dM/QAwzONCudpil1t/3fNt7WCjXtrSh4kygEGZlUffOY5rWr8m5DKjfNR70fba
9xgNIPOl69yP2HznAPdXPGxJtfcvyMVoePajNXNG6AUE4pf+ekvrJ2S5QLmxOE69soye7+RZU065
GLx5ZQq4iahjsVf08USXOUKbJ5lqiAOkRtsKVGK611XSUWC5PV+iU/zrhmOPuphFpF8JUrvf4frd
tivWIL4iZ1lWV8jTII65pYtrjfIy4tuT9cxKgGR4MvasSP3Oyom1ik8PkP0icAGc9b9wZTVZ7fEs
yietExfzHuYPjXWZzckihwjUNhsxE4VefzTNgSmVNqz72CD0UyRY4Tw0oJpAp0c6vuqtrOpuhWkP
5BdyF5j6bjN0qx9a/4pfDW21J+zEm6dOuLIBASt2Iqp4aC1iK9OUmKMv4TlqeWOwOrW2TsqW3oZL
mrTOInwgPL9MavUjHyDu/zO06cuJGquwB95WJob3OYhnWaQ1kpSs8mrD+1u2NaiFSJOmc7bpDnvZ
1gYbSa6UWTZaR+ap5L7Bjq+kuinnKComja+2IPNKwfxEhViouVxNE6X2S6k6qK+cyI4NA4RTYr54
L6QdnhmG8OA7Bn2786Dui+wXmfDQBUiT46ZW341uxZzfYLANSIle0E49gnNU14uWcNDHrDP7qslH
d1QePCB6GFjFImuwBK86aHLaMX/XrxLyh7B2GyA7XD/R8SyoShyFwDDZQKeHJ9u0TAxw9+/7u2eX
XK1bB1Fcm1Y4zRwJ3qYX6A1/URyrkb81xInXxhatQ3XxuonAoIAYNEkT1Gql0d5Xi/3A1xKhTNJs
U3LgRVaPlGgK9RxUC4z0arN5ga2mCZh2BlTBMtvXqvFKjWGFzZ3uo5nBxJlwrrnNOQM/X7LlqRpR
HdbkpNOCOP7vNhsw2Ak7qK2HTJZ/xsl9zoYU5rD61Ftra3m8Y4nv7w6NzIByMyi9xCvmulUXntrK
K0FVkDsL5yjia5jFpIHg9VqUjmR4V3LMYNv0YD87shDSHbFUdEo51+6PvWGfbZgV1ED8V+LTMqUh
aQLfm6tc1lahIvjp70ajaclphgOCPnTLpWrfDzNp96ecNfj2TvRHM+8yNYbfe2jKnBqRxqHzArW8
zsnEVEW+PobbEKncL5LHluAVzznjnr/JMGvIPCnA0OnqHjZMB2hxNRRWBVQ2djwQRHNTWbFt/REk
+Vyag3SJXVWClEDSrQv/SvjmAlXnAyqtWqJ+2W2n1/6MRgJpG1x+akvmcg/u6/dUgnk1hFa28UFf
drEAsc+d03wh15+rIAwTySAHWvdkmT4VIg7sZ5xeEeYg2P4kvPgsJXFw3nS5F6aTadz8Z7WPqMp8
E7nlAF057YuJAvLostOobvDODL5HKd5l1JaM7+6wB2f+ewn5zTgrVMkn7ARigpsMzMT8NAlgqxEa
Ji+X2yFykTH+lbwzWVAVG90suoxpdxTojeMtrOOp5B1wBO0ODFecKVxDXfefnYcUUdC/RJON/OJ5
CG56lJKoCD2W5uuaW9RHQs+GLCvPFq3KNBB93kNJRveXBvqwY5CNc0omfgl3rLNlZ/zbPtvgSEIp
f6BbzJ+2tJFLhjk5iG889h7eyKrY1MeknTJEn8HlOtMu1NaKGI/VXAkH6HXcoeaXXcbtQe+Yhl3J
+c9y0bK1Q4I7LT4FtEVm6vOmHvmi6rrYZJdhHhNTkvKI9cDOtmtijJyb5lHRTGoRBlHoetxoKER4
gab63XIGLDdHbn1vPkbPck+pXDeYydk92fZ9Gj60Y0cWcbBbz3qeEes6RokaJeOU8Wp+YHFiBPED
4dI34Sye35wD6LSt23qwTnF50HNBh38eYGlSAW5BYKviW1klBCyGnNe6YI48KwC00cEluJ8T6X0T
j0yLJUfTHbnX5MZHzFGdyFmGHIBP4639naVzjR+NDEMUEnP5EMsU650Q4j9A3ABCUP+sKOp2/487
xtL7lHbIteYP4UgRplpiOgkmhKwBVkDwWvFjxkGhDWCKb+SqjU7H26w2M22DFfskAtmopcNuInL9
bpV5Oiy7M9PVSb9Mueqpq0xUb/YRLbjH4jkrrje0bRhGyl70cs9Yn0OVfK9zpkEfNAYURf9MTJZI
wdvWIUEu5ppT6xJw1EuPnBeqaD0A58rEuwzw+adEMx48Lv1WctsFjaAO065U1Jr8pAOFdul4wyR3
nP1N6MUv6HBPglx8ssF4AyS2QWDOSX+XbusmQrAc4n2FE1/kjydtcSwKB0ONUfzGy6NQpB9D8O8W
VJyoduvWOR5C52wbP6jUbAcF+WnR51FleLduSyR9O7dSpMgXwjlAXjr0BpagrN+PxBmA+MREMsPX
g8Y26ubtCiQ0FaFcXFG1ckSiPhPBVt2MUnze7E3stQ/Le8eOHu/BKW1rVKR0ZCcRAUEmo3YwdKMG
5XxTFpZQjzsO5pZ0upmsZ7w0SHqNeizzI3XSeWWmUPYw1RIjsYEGZRvl6Ys3sge7z7LcZxFA8oFK
HDs1qPLF360R10uTwXfeMiSTAm2f8JLuGWRDVhxWop+X7HT03tWLFcLojq4rdCOAVMcXfS8HG6aT
v3wPcDUuL3sS2dmiJQGqsef7H/60QL6pnLF/zVYvmqqFAunCya1IlxsjftrfqDgntEoQq6tLFS3r
FjKOXbwgFT8wWb7lJxsUNqvqHBQR6e6gij3v0NLE/Kytu6asM+h4c7GK3uy+MNaxmA8am+WmrHaR
U0rwig8eVVA0+dLxUXrZ1j3TrqM9b1dyNbKhr03m8xRsuv+aXBL2J29WVabjvGjxjIQTOxxT/MVl
bI9Lid6kpfn3C+rRxlVm0otkHRPEwi9l4Mothcc1CNAngbdVSNplrfZ2pCfO86CkjLR9NgO4Ki/j
kHJFV61f1vlH57QIQEnGPl5N4MB1zoBpc/a3O4L3UN7aEOBeP9hX4+O2bYGgK2Jljy4XKryCakT2
IzK866oyTNuO+/3xUNcXtgW37DFlJaCYBJNM1QdxjiMTsHzyaqpm6VjeJY3rLsDpO5ixANWTz3J0
bRxo45ms50EmIexfbNN2iXjr9t2KPkBYeFY2MVnfU5C2wB1eA5jwoQ+6m7gNOojknNAN78MzHVTV
ohQqZhwM6cUT4dwAOPt9IXUJWvMvPnwb4dAIHMIuAfBsGKfgiiG2qgR5tZzRu2Tvm5zRTK90viYr
lxszZTFSys3uxHSP8wbcsLJeBQ4Au9RfU7iPEwlk2aS2Ce7dMYC7WaHad2Rs8ByqFt9HdimDmNzY
hHlh4xddIcCaM54hn5fjlqXd6FOaNzK3rFmX2SExCsh6UfegvS1fSVlVhnCX6TgY+DDeG0W3bAU8
zQTgrBgfGSoKNBffcV6OLP3EMcUnasJszqOZYF5Gt9YLkYbsNO0NyVPYoisyBIoYzDIU/QIXMiXQ
cXMfanu5a3fUZ5vsTY7Z1FmuZ5LlBi04oUcvSoB4rTAyiBFZ/46o58qJf3ZBj/toQKrnvNBwo6rx
T8CvrSpbWDIsY2n1Xy9adovTF9G5cHl8CVqe2gZ7t8l/3Lzx7P6X1l7RMCZHah3/TMKefkz6cDUH
lyq0Zw1O3ytFkb9WUvSFp7+ws+UQ6OtkAqqYSLXV97ODPBFTFGS6i50AESQufWTRdT+CnaIUognW
PhStOZdKrxvrkAwdKowZ4I6nrK1TEJzjv19a7w4hPOnVDcBL2krL67PM/O7K5lKXdRQ841LfWOf3
W7IWaGNnFp5kYjNqH520rj9LS66qo+XinH1xhOidM/sP4mQ6sLGEIkWz5k9jReqxDxXcbHOZ+MMm
jKsaniUSWXfyjXh9pvR3cIPY0d1AgGPoOCvvm8SxbTeVrz01m4BtZMcj/K5jmZR3es1L4rCOkenW
7oYBqCXB3HQGXWd4K2BeI66R/cXgQnn5jf7M7UZ41iXEsiUEupjQ7wJEZkaZmxHKoPZFAPyLNUDB
XmPNxdXwQdFOvRSvQEuocaCsFrs5qBklr2Kqkli6KfZ4d/uBgVwsMZldIYxMGbgyEqnU7w20bq2C
IqJp7fH2rz61Gg5nrRfxJ190Fy7F7yEaioTOyLvuLXmllW+6c3DlgVGZjLk6oHQlEj0ZUOREVEk9
LuP+wZQS9bBu40hR1bwvsSAHp/6aMlUDqTSwKfUZl+Lhy6Wr4c7aFiSc1moKuXMfsDi5VBNtXfCS
IvXcCjol4MgQ3pcq2V298vKHMtPMljBCRlTtIK7/1Msclb7UVE2+xzD03kOdKUuvXoS9GxGplQ7L
l1K19ZuinouHQInMoQhhUXIDOEGomm40V2S41PPYBUnMHVl9eJbkvM2T5eBuXR1DzPuXHE+uCn0V
t917g0+fyBf3CEkwnCSNYu764nZbISZEKz9abOKsfVe7VW7m9c1CSI9bd3qZkOUSdVIR/nx99d1r
qGiLVWUUq6EKOEwfCSrlpCdMFvchnHHg/3DDRoNWlq13xv/mpPgtb1L0BEOBhNnm2JEznFsCOjy0
Y/ku8l0yvakO/VxYQLWLz5ztDf5b+JO6JyzDFFuJuO9YiOZ4fT/odyrFbuMOld69mYQ+UJk8JRdR
4SXTbENq3kN/53PW5Y4R4ts1V+cm9upuGxmKs/c5Zkn4Kwf4mux+PyspTRTB2oghMs9Ar5JzWxBH
DNLg14XJqRG60ILQF+qWHEpsnrK5+dDVm/C+F5kObUaJw3u5Pm2gDDjTihmGW6g7CKwzThZKHXo5
CeZzC6TEyjsr8nOZGbn8MLuZqemgSz/0z+DVLPuUhP4Kh0X4appaH5QzEN5jPwvi4zI5Egdrkay4
rlIzDVHz3AltielPmahUXHhTdimSTAeljh/2cC0H+mVWEx4u4TAcxmHAhaZP5jHU5Le0YAqs0dne
7mMxJBrTdAhhksZLSAG/nCntT3D7HMbi+ppzmGXZF55uZgp8LOwK3X1tfTKOyqzuM8AR4X9Hgt27
Pvxv0c73au0QqdtwYkswyggX9rJbASFrzKO6rLF2CUi7fmb5lDSwLCxO3/RgEXgUf/bibpnik8jr
h7zI9tcUWYaoW4F3BpnJgNSdgIeMALRUDsqCxt1pGAWFcb0SFm+mt2wVp+heWw/Lf+v7zDLYpfGr
JrYQLXv+0b/xjwCxrK8WFK5VdfOdwiuzB2XJr/xBBhyI95tf/RQFBgVWGE3o2GRYSX+pSJcgko9o
oIKMzD8r/P9sVBFRq0Y7Oaj3iIsMOLdJRuGe4DZrpHGFm0glD0J9Q3yQkYDdFULps8NHbew3LeuS
L4AI2gEYx8lsmxGaM3i/zo6lmHAq4EzmWECGW58LWLlfIi3F1ajQZflitQwEjT+UsLSRolR31/km
UMjGkOhVT3/t/FkNhBjUuy4AS9gE4q1LLo+8jBLFld1HJYzRmFeX/4AWIhwT7kBfdfCQYOvWSGxt
vRUledmRZBhSQ0KrvbQ9Hu60u1p/t1mRPp5gXAnMWbJ99SjdpXcgHvq3vSUJVkka4IuN6birY4w+
Y7S79Zz0mL4N4zDM6NbWKbDNLfv2J3ld3lIR6sQH4LNT0N3LKkaU2QcqL+GTvcd3UE2BBeoxvOqm
NcLZsLbQhAx6CnCfkGlnPL72g/lc6try7+UamOHGrexTMkSoTY1CXgMJzDVfYUhN3ccDrx8TpbeV
dowktXQs4UdCPnCn/JCy7VRVxqZGVSmGVirrtT2nmBMkVlibX404fg4LrJ7TI0QKV/nPniXlHt1M
oNajffm7ugjQ4DIxyPwUl3IUJfgZXwRYL8AJeystmGDc2S4c+NMIf7w8o6M75ukq6PQssEvcym+d
nGoMh/fDUiV77hSxSKYPZlVCpS//GooTmCzxxEEKPRtXJDP+Fi1Mv0328TDGlGaLOoZOI9TIr9Mw
XII5mgYCQ06YKRoiZy1BpCY5XnuTmfANKLasuLCyUZ3JhtgHRa3VZS/FYgJn1Pqi/hms0C4q8QC0
NqvieaHrdklsPJn7mVFhj6reqIW5Es/DCVIUsxvyAGBn4qqCBbnPA1pF+gSnY+SIHIClnVXrCoJX
uHQ6/7ObhLggt61q+7sIAP70SUzF15s20qOI0Y6eAG4qRJV2rIBxf9v8c/mhC7PdHMSDM4mcRUeX
WxlpXYtv5FZ6Xco9jiM2vcbxO3N2d47tfiZDCd7pQNNPunny9niaL96Vi7dji7zl4j+IjTOwp5Pe
CWbdPXNBYaVwXf7KTnk0s0IF/DZZdTOxtRxcIsx5n2tinJhuFpTV8yg66zVUG9aj6BYY4o3ddJKJ
awv+dsHQngN2W97XfPgxvxVvXGEAu8b0Zfxi003DAuGvo1d084eWitO897isH2OzkHgx5tyxuOD/
L4bquXGFfzMWUB9MEH5LB2QAnrQ0kMlHd0bEpOQ4nQA9AMWvvd9+S5HQCrRwS2jcioY8kp7I3KoY
QdYXkYR3agsm0gusLysr2Qo8kDkX8Tqg4mVnbLhz3D7qNoZr8EueXxG2iEicaEnhBfQPyMkwcI/A
RDnMbGbgH/kPv8KziK5cbLHdCycTsC14QvK1r5xDjAV+Y55DxGTEErt4UIwRmAFOPT0P6liMzS6T
DPXYUW86MXWjNAofMxskiM0WhO1v4jDIjm/F45JCgMwoXvVcBxYY4oYIh7BQ54inESxwx0nXkX7o
gByEuFgOX0fFgZGe+rJZMELjd9yJtaMtkwMnTSiLpG29quYV+mgVv5asgvlF0ubE8ukuxGq/L4iz
0Ikkio9COP3dtEQmhdkZb3CDYuuaQ8s6zLy5Sco8yiGzT+sjdN0LMFXJnQnZ6L3cho2pKrgllVF3
EfDsWb6StbB4EiqjCBiECLAJ7bvgUpdHvH2yCYHto+FFbUUGOlUDw8gILdtE4U5X/uAwY7xq4sFt
yqvCtr8U6kfh5EYoFaG/XyNEZxO40NgeHtKb+9VsFB5TU7MyJ4DUWKhBpjfpqsXMlDqIAlP+8d5r
j+Okul0MVR5q8VyuK1bgZq/pj1VoDVNjV7MkaobinoGYO1jStKyf03s+B3VrYro5gVuWJIqs8iX2
OCF4bB5URqEYmPucoTny4Osy5hHHBkZ8pmMV7TgUGlqbzeTy6aIKl3AmqntwFcfXS1/K+jGExCMw
1W5wGBvFkajRmZhbbdgOA07+XVk8wSSFDBi4s94fKwb+bdxXHzTT2kQ7UCiX11YFPzdMT2zgDL/Y
FxtAjiUG/Sut1V8OIVXodMKxg4hgZl6/wyYAB9VRJjjrRH0XNiPmqrU8LZ71ZSzolRV4uPUfs8WZ
gSrlVPR2IJzVfjI/UVhsKvuDw9/0VEk7wLnPtnVzsDaB43dZQ504hq7jBq3oOhr295CstOIeGE+w
tWM3SrhnqSMtpqZojtHm4xIPUFYqb1ESzi2B0gg0xQ5isjXBO3flQlmexEckFx13j++mPI0oVfEW
63KNDJCovn3RYPfVnHkxYDcRmHFwVohW+BjRyYK8zREQ7/+JHE8pv426DgqXZ23rAMgeQ9MvOkBM
AAsrGMTT3JdWiu7y/gF5/AVOXzRLiqA80lkcck+Zx9watyJecSIlvNGUE3X2Msvogn0Cm+ZPtvKL
8EAYN3Hdqb3gDQQQpqA8afwK+ZNK1oEycqPD1d9N9CuzJQmYyfy4byhkuJ1kJeDZVxNuw0SOZEty
4RzDfjUBDD6dNfwqwjAjk63IofOqGg9GmIlhWgcZ/VZ69tJ2SkFE00Y7qYwOyN7aTroQ9nvQMxue
/T7eh10xljLz+0xe1gK98i3VR6F+irsRlrYk0US7KR9vdZsH1wQvyWrENSvMm5D1sHos0GPF66jW
GyRgWzKk0cvsX5MjQBIaBtg9KRk1KXSpkTu78U4NIeL/8NfsJWFsMO6Afo7Pit75EMm91Z/pHLPU
XW62yRYH7Ptt1/22P7XJ89cuw4Cb5MKV9ScOrXwXhKu4HaZeeHFXUdx3Lj2Wn6TfBdP+4FpmLbTB
x2WzvomBa5/5r0hvh4AVq1gkJozFZNubE+kqFH7BrWQAMAWgT3y8U6BwB6MsstNTqJ8uOaD3z9Ug
/5+ZC134Kdd2Svv1W0S4mEc9ZyzQxdj/l92bA4A1bJ41mk670hbuKWhgDeMszPyx5aNz1ceZdpBT
WsQiu0Y2P2qUrUBMo04TlXNWgl9QCt2/r0RAIwyYEEZAR3MoSPNK/oQQxyzCCiVk02wwlg2ztNHr
hYkKv6ja8KZo8TW3cVIC+Lss3nXVDOOj/bLwUkTu3floEwe2SOWOUBcXkIA6N+LEPbHbaRxNcfIc
39JL24kGJG0H/YY3jk0xawnG7flNme3e7fzCGnzqMOU54rO0LZ83Ae4oyEvg/+17kpULlGtic6vV
nOJCmyyqOfuEnA0I360YNwFpvt+kHumpTpNJXW9IQNTyHhonoJ64osUnu01wPJDArKRClXuxtFUi
RpsrfNQ51RdOTjY79yu6C2ckAQvqwI4RhbfHvMuw6hK3fr/YpPq0w5KxTuVOPuP7xGnVznyoCk1R
/QBOEVXGijohKBKfE0LY+UUl+p+WQ+nCJGAObWJ7swKJBtadfZa1OW6J24ZoOm2gkwtVFTVnrCup
5g4I8NLrqk2g/9bUfLP9KCCIEpKhu4oXxj3JeWHhvN0f8/uAyB/9PHfj/RF3qLmatoYYPbpDR4SL
fNsZsB9cBGIVpVTtt5fAaekZClRMOjin6F+dEdYcURk6UFqsj4ZNH1sVUtIrIoabADras9YKjqHL
5IMK94hwFzBMf2dbZQ/7W9mEuFALdQ3ynCa3hwPn2+72u2s+9+luoqBrU6PwUr7B8IkmNdkk+0WF
H/ToD5xWPiNzrnx0LfyPe++DupR+oyKUWDf/Wukv+IN7pu1xD9ZoagykNhyuMIzAFw9verZ4Tb6S
14jA/6WhqWA1mT51xh9Qec0kZXFCVoQZSK7y2TvgTu4gsOqAuyGXz2FFiJulPQ76XvwTehCwAJfT
IBZZk9812gk7VLLRAY4ovHkbIddC+jw41cOruUnJiWibpqDJFkOtNXK/yAnfz53Sb9ohtBewg1o0
knExngiQqOnjAKAp/F1YvCM15RHUEjd3Kn93O6LGczeLkfF9arSSFurFhgKnvX/o3xJ+aJWPUcT2
e3zfI/4c+9Jg46XhFYnLoWnRJC7eMBesjUIEhwrt32Os1lSDy5I1YXdV2Xw+FRDqgNSrTX8fVDqF
gPEPM4yL+ZZSPGGNHXdcCblLGrAoBOIHCSbNSxYU/doQObHKurapmGiq8HUIwIZZpggSJ5ioIL2b
6mT+x0hGri6vijB6lV0Pb3GqhRIsVqP0dLDjeY0rtLh/vREZadoDoPvJGPWngyu2X5bJ7iyHcz2J
PelUt+5Rw78QwfeU475JQ1TENjx32KNomGw/06fbnvGXPtKNdwFC2Dteai10pBZujGEBv4+NVIy0
PhsjKErnZP5wAQk1BlTwNrU0VATzr5mRe12Kduz/UpWkAshfYmIC6q+2ZbD6N5WfYDTC1Tq4l0p5
qi7RtPgE6M4AbSICt4R1DQM7UBLX+4uC0Il2UFwGnzhrWguTAI3VbfLGEpdzuOkNlOJmThn5Ybp+
dqFm9BcOMIDly0IVdt/HGMGQNxhP5lQfemjjFpvViMw2vTy3fxRLtSIyvxSkYNKpM+jIGeoEYXCG
rDKltHK9XmXD7j+6MCh68g0UCs2bXAJjYgyEIcXhA+1sd9dHvtOqSJdeMJkNS0qDU93bl8iGv6kW
2WOnFZjGMJVOrmryOF8jQ8a6cxGxTkHbYMqTX+4gUWwz/FzCEhv6m7ywSidvbdcLIZx/tjcwuh4I
Q3ToqpwNOpZGSqLWbpo9l9g5YXHwUHKpaLnsu0jq/RarN9n7Kg5B6tageHFeaOaZfLGJmFIrM4SI
v3JQ9cQd/OzFz3lJDDmmAPJ4T69TLAVIsOnGe2KoHa3lDVrsXqycaBp1Y9tYLjjtixpSatX6AbSK
U5hIsFaoDwvs6FPOC+UrpYe/P7sC4YH3IvNBFjaC5b6rxFY96XJTEcmIfT4DWd1I3S1tvW3jK7lO
Suo9Zm4ue3pn4SxWYDJw/PfPUaYZW8j83s4uRNDUPIkpRc1IQ98cIiGYYvBMUGjM5j4PhhkLH51n
CLvw+b61SAqm06fmQON++EFc3XHBODRTuVIBJwuM54/ZuISFCyGbzcuIsPKEj7y5XiWy1AscPBfz
itWOX9mHOB+V/n8EOc3MOnMqsjip4WfXTrd2hZabDsVyl+z3amdE30kWoLdn4aYDJN1buqNpGce1
6S8klRbyRoZLNvKQ86T56VoIl8R3DWPeyZS5AHnChG17OAkFHwzXcUU7xGo32GebNEnSUqUrQwCv
jKQD3yyfkl93bvUDrPoJMzBUva2WuKFjp+0V+rGhw4OhoiUgT/q8KV/XeeJAVSmuu7hXNdDwQaBC
lbvcQGz00jv472R7M7+Nnl2bAsrM1HVutkUJKfiJ4V38M1nmRJQ3hAQmFfRCQeAtO2vdCV679L6P
oN3cDzYyE9gcwTrArkjqZJ0+gx7Q+NRTp7ZVsZtiKL+mR+tzlQ6FVzK0hEI5JuUNjglIWTrNV1A8
Hb9I/NttfWd6QlDAq4YVgtqpsJCkMHXGB/OpWyFvcVTotGLoXBGKugXewaQWgVOvEjK7jjdzZuvO
pphH5NW2iXmkBaJLiuvqXiifuL9VeXzNe7gsxiIkf9ZU7Pw2Jrc7Ch1+pQ4FwbrdoLfMLUXBP3VX
c4G/kS5T0IJ6M03u4k/Cz6lOrIoPGZkvNrctOofdaaBy4TXloRSyl+i7ah6qoJTT3Ep1vUfwnFNw
zQYQX+7EVK73UwYY1330BUAvbjdA6SX7BECYuq3AFkJNQlCWApM0PXW5u4YnuLKTC9hCJUzj5SnX
H//ZKMXDhJZcntvR2mqVIxk7bwwSU4NNwY2tfojVVnldRZYmCTpsiLz9ldbg9pcYf+PxHOfNaXLC
QEl3d/fPdWv3YEhZiHDXBOERwzXwGpxQMJ0FxEbJD7HWdIs+3J/CiiA1CTF7UZxRKrZYbk/EfsqL
OrR2ZLvUt7njHWy6DkHf/mPQYjH7jn9xf6r2nxpNpSswzLfB5PyGENplOku69FhRzyC0DwDfAtI9
jzKsvPq6gxt8YVyhaVlaL7yAePRW8p6EwZbusrsbiR14cMuA1fVJb8oWzK7Hud1kBvsVZZuAf1Ew
KTLDQ/dmyESwFm/KENP8tKqMhrPnDNJlK55wcmtV7ZTsYdtrhgMIJH6Yw2xxkrxDzXu+AtFPicsn
GCHAYLnFkcsmTyRulqH8fqML6YMqKO0Wu2EwcS9GafDJs2uznGTV/5ihcanRrv4XPDGVrHQE3Aqs
odNvjYt3HK7oSkc62aTXMYVmApGLnI1Y5KQPJKhPjhLDhJTMfvg3zuriaDa5ivQNKIgd4lKWV3Lv
fMQlFjoi0dxsaZcdD0uL33yK1ndLO9XTmRGSjAXMk9Bk4T6LLy6bRDqYzeeweGW9UVZndrcqzZOJ
J6iU8nzOftepHqMo5/X2RnHGyaoGdGtmwR5q/3kPk+D7b94JLXr3Fbf4V21h8lYlRun03fS0+RNu
QaopvN2Y4AD7PKWg6etoo1wpVIn5S2rFE+mxPZydk7SKKuMGF/anIrnKN38aOKsp1vpJ2Xu/sdrg
LhjjABAnBnaI+95v+/azawJF9dWH79So9j/+qKyr3cUm1DYFeBrDWu2LdbhAXhLnIZ83o1Fjw0qM
8nuQcHKNUluLwzw74owX1qfJcinYeSeG8L6dQMr/0NsuMiFJYCpSx50XtPlRZOS4R/nxpBTynd41
XIauVwHNrDRiHsudTZ/tNIEQ7Js7KUyIduvIKlB9PdxCpJwHbnoLOmehEkmLYVFb6qEkRmOiK++Y
IaAR/cYObmGjDyyWjkPZsp3tfAvydH8mb0Wcx467ZVJDfiIZRjTlonocBPaqMrf4SQz5Z/CKBIO9
6vK5vBBaMZLgGBtmpsaH8g+j8TwXN4Qf/QD0zYuGrH+1GRDRvRt56mEqeC+Z0jc76UFvbnodYmxZ
POoFdgde0BhuxrAyuFqQQv56tgjxbf7ipxnxJYuDbijQTFtxiqYKHYJzLZIoRBmPwA2awfO314LX
lNyT+sbaoGFdqBNTdCXIwZn1KbVzy/ufiMJ/joWGhwqhxMY9YsU1emFgllC3zYsrREQuW6cOs7+9
3hjLYMFbPX71qXyzD9gaYcG1BZ41rjreEnVlwk1e36Sg1M9tpt//fnxabRT3/S4mDt83UJ5mFMAo
ruKT1NznRmqDpgIRg8+XrtBIANh4c2FbYkF6qcND/9F+dhQuYpdtxKrH1WdB4B76HEy+JN8AsTey
zxJ2tsLA3OnE5rqY3tjc4AZeLZXcs+U8THpR97RH7Q0MrBS+hpIToDe7ItLs5btN+XKsD75kSYRO
fK+Fs9Zo1JYkJdKkfLIKxmV59UbjFnRmjthhI4bGeJYaQ3M+1DKF4J1JRFFDCT65Un5DY7j4zL/l
yEB3aCQtAseL/YsQaRRGIHEdUoPy+Qn3HbKHf2bvhb7J0OQzy7QE7SxPuwUpbjOqrOoIalgG2qf5
oDpt8qEbdgJ15Nn/drH8giugfpea51lRWuGRPq2KZsUk9E9HS0GIPzmxhEjOfah5zGK5lMPv0Wsc
MgvD5Bpi0ylfL2Fy7uG9ycHTc63ffwDvCbve33lx6lTrKhsgg32gZoa/pvfiyDFJsiQ9r9KcbkNP
j1Yrxv7JNuR91AOLTbxZ3kZrWV6HoZEqGM68r9Gz6eidZNNiHBVeTHIZFZPFAdFH4WR9l+/oobb0
O8IIWd9IP8oWgXlgvpFr0QEv+orgbPGULxps/V36JX+68z4PqNaBCoTYUDESe4P7R9OE9Yj+Wk38
cS1rN16r7do4mSMhkpUXbJ51+lUYIsaS5Sf+2y5mh8SUPiHQbA+rbi3cHtdh/6zBSvq+RWHTkTR1
qXDvuDDEXcWpf4f8jLm5aVeR8CTugvCjk12WvYL9OwwYq6f+e2/ThOZ1I7Oz9zNnLC8G7ib/NRyJ
VWnSDGNDCBp1IKrXgFgM4SWoANvmVEUeZUablBnilIFjWyfiCxWaz34Z/DaLqKT3EAaLLpjFsTYZ
J4KMZRQcyZh9NZFwbcv654fNTqvN5KYUmssiQoo7Ro6ML58u7YAsSWtZruZIcDrFQaESugTTwOfR
JEbW0FqiaUojwe6gFItbH7nUI4/6Ib8RL7VTQGXHMB6Oz5HHqkEFaZ5siT5Xa3ZYAYdHAVPxUPLM
ti+5GBz2mfZ9sm0Kjn7gxq69lVBWibscWPCo0oq5eYwQMIHX7MHneKQD0hkJ8EtLqeH94Q6O9LlI
hhyRa2X+qp/6Fl00Jwdn3IY4xX8NtcgXB/imHoe3ySqN56zswI4+YH/OCTldgWXme1y1Wv/RayL3
Nu72IvimTTuGtxxyb6k9+1gQA0+6tkLJpl68SZqWl84YoahQVLIps7yu4JTUEngEzFJu25V5O8q4
5awKeYo3m96rXaurtZweutaAPVH7X1EJAvJfw4JjRkqVlifyeX+5/GQkEJdegO6Q7ZSA6tlkCe4q
EpkqTgYx3+/pyrBVTxXbayfOdnTLlwRBufeEw9cfAYyEScBMy7vAn6nEumqIMJo/R13Oain7U7IT
u7gbI1/QFaT9Zp5T5XRsvtu1yVDqCRjgn3xcUswYArRJcIkNhOoG/NKTW2eyog9o2x/mWsB+otBN
v7NgE1/g8aHY9GA3JOPywPQCzH1GEw44tjaC2RFMGO4v4XOp78+0BadJF5a+AmlceYWFyZPhs4vt
BVUJzGDg1G3lvLwtw3U0DdDDWMy1pALfA683H51cRry0vgZW0oNN6gX6oUiS/JYmJxKSOHZX8aWT
5GCt365NWrvRrrkdzsH/i7Jdc/3wQv3r/mwA92uyukfO1av9MRUr1wAzfC0Rnq8wICh3FBXIE2Y0
J2QVHEeElUhUVy3LAq94hcP6unPT1NrFAdiNSg188KbXmCS6VGwqJfC9hGvjHEYxPnCojEKbpgQS
HEurVKjuOTcbCM7noNkLtWcLVO1sxuirgM+Eu4JkcoXURLR95oVNa3p2hZSXZmMaST/SqGHyW8Nb
frv9dgruZv1jz0xOAVlW8Iruz4o7UNM0VI+RZS5j0FJdq2ftlHL7SAx4C8RaTZrEXoR9KahUQ3E3
wxtEVPtb2zTKLihkl6pnrRWvvyEjuiMDIL2bT6p0t+5exM1+XA1V8e0D+l7eBd4Ezqvy6UD3bzZh
94VkaMOOjRyxne0pK4Wzx9Jd7eaohmvaaEerChJOh94CPpFylPmilno/5TEALFCr5OAuN1Kg2FCb
KCgZc8XpIIcXMDD8nAYWBOLBF2qlMfbsqOItAqlcg5YUPWdjI20kwgsQ47ZXvihJxQq+NdofmShk
edD3gX+NyPag82OEJGOjaVtmn3FWoL5QmgjG2TJQrlCGpchRGPxZ9P+i0wsquyWkuKo/hdrYOT7H
eqmPf66xweV7XfB1kcrMllwFHemrlhUb7n6Fmso3x3m8BpXUW1/b/NQ3oymzVwkXg1htnN1SBGwt
gvfEwyFFLIfHVGe1S2YNiZFUMPnON1Roam/rwRTwQFEijDpII/XTLCu1JyNZf5tz+eo6LJ9A1RbA
/F8WCFw+/DPQFFWbPnKbtNu/sL5FuvNVlkMqzb3aP5RQ+EGQxGiQQBpninnNU+deOddDZ4cNswKn
asJtsB9IFDjSPA2p7PheSKeg60tnN5AlVKViQztnjHOXw03y3QB5YTbIdJh2wUkr6SjsB2vxPK/9
Jd43SSqHC0BTUngEDJVIbcWfY5z5x77LDoJKsbGgqJK60N5IPbMdrYCwT4Q8CqTtCMGUBvyQCq2w
JycFbIlAeDXgxJruCmRAqcmkhYyR/gFy9/5r0FHYVL0bqp2XTcEw2BCKIMkKPWDrluDZqN0OPZk2
b1wvrW8h1qaPLMjr9AgNkTa9zXLdweSyES/QwjZDNz0EL2UyEUDr0AFb6fz+LXBTnhzEaFxL9SBy
W/y5pwGNCKa2A5HiX/CbWjEz1LmgLYzjFw99lK8A6y5pnHNuIosjhAdboWy/wLXeo40+0iYhLu9v
IQzKal/5KuW9FJ4vk0Q7/qGMfnku3QJFPRAKdy5iRJdOXaId5Y6Px5uL2PRpS0l6b5ULgWEV/tzb
gU2f6cyhFNrOvFHVca0dafxShJDrwMkGvCkpDhIroyEKZNQOHftEyrkep2a0o73uxLhO/iDWjw5o
o3FdcYgcAJBdZvXNVymz8xUwn2/lYq6CGpPTcJoWxr8V5TWQiaysmPfnd9jA/j3lkojzMFGFhWS2
qQ2pCIfuFXnn86CQxgAMsiTI1MHjTWOSs8HRS5E8OSe9Xiy6fiYOjSfkOVb0tpripeU3X9CI64hx
6S6FLOG67r7Zmru3nGTiQiNc303G2VZd/Mt8LPbwU3xBgq2h87NT83wbevBXgdZesH08Ae5x8wIp
QULE6726MIjZLZzT+to8BfluH/YeSdcdQp7Fh9AUJoM7wKYag6wiq6DvEL0t3ccfqNUz5sWA7ikQ
bkwEw8zS/1HXouFWeqYBS9Qpu+j3dzOIJ21Nt+YRjI55KvGGIbf7WhRKthxL6GBuzPgaZ0SkQl3+
EksQBTx9ro1snbkZxHtjlPDGdyhHOjtcUqaNl4bbtf8JiaHynSFOVwCTM8FI7rRGi2gxbcdcZQ51
lXP5HD7ojc8ua+GSJ6P8PSQCFyk9Tc8cU+yEBOY+fmuqlSI4fqXhoKxa7aaHnNrBxxWhi7wJQX+4
/MK8AVSgujeZ2+89cRF3S/0f8z6Z8UWsFHwaoBAZr666PzyGpYpi3X+qpt2/XA6dOneWvtZ9hUIk
kAG4k6R2v18rfMK0JfY/C/nCKu78h2ZwTI2AGxi42JgA6shoCwQabfcfu2pHjZ1QeFVX49++sL4h
7w+dVpM2q/kHTewrD9/94KRtc57VYIT2CjlhlNmV8qLO4YqeqYlxv2R6/P33W5md+FbXA/rHmEya
xcKWDnpYnY5PNCzdbeuMsMR/kNoTdvrZscO8XO9SstY1zFFgXO3NS6aRYhKkUoED58c666LLISIM
YUPJh13xLWqE3GdLydr6oZlinMUOFJC0cELYiTFZcQr/YX02RqJFKqLbR+NhtUJPizcgQseWYCrf
1gwtQp7pxRX6SmS6F9+g+O6s7e3k97Ik1Vhi6tFmF0E3Jaav666JeobYMEuVNO9og+t30eDGI+TK
vjuvC7WDfhVp0OUstH/80+UGBj7RyX1JuAVrYAu4LBSCOcuKeGPHu8fez0srdDiCuV3nTU6HR2k1
n2FwDflb1LeNwjV14rbm4SzupTTW3RJfCS25ThY0p7YlqY/m51ME8DfdNPYIV/nOb2JdC+gE1djm
Of/MYfTSPFgd6ZwvCzUr5DE6/ZZG1MPFw9R7vmY1RWLijO0c/68/tOSRieAb05JSkbFVJ9PSXLgq
5YKWi8/fd6lqq8Qxge4Ry4Xo1aGnA+RCTzEAT5Lxqi0MeOmlKsZAJxPsgLC78ETjmUg3nydZV9/D
mFHt0t0u8hgfsSAgzoba05zTiYEK4vPpM4QWrD8M7dUFwqFmESmnMU1ZYCiJ0iziq/XTSTigzGXI
qX3alMwPDy1RpLBBKaEqb+V4WCNkksZT2aENy9+zga/Kn2xtZloTw44qoEBGmBRZD2VHMgwwHI/3
GWcJic2JlN+wNDVu5pW1z85vzuCnBmw/mqOZ3KsV6p7RB7F5DhqL3fyd3NXG13SOauqY6EOEqUwB
AwrMprwvfxjAFbS/uXUiXpFpD6G/CwHA4GIZ2MJEvbfZb0202QgXnq0xtBo9yBlUVacMEzSURVpH
pn2mVFxd7aovW821MgUIAtYzDTOkf4eZtibKREh+iA9Z5SMSishJ6pkyPLaAmcR+S1R6KfxMmQoj
Eufp5eJFC4KUZY6Rcy1WAxiyGamOa/roiAGcRpFdhvxOcs/xqSkLdf12ogw0aZz7S5klzeABbTm/
p81RZ5AFPyk1F4Dj7lSlnMeUReZSkPewuxunqFtvqqfV+bvVeo/9P62vOOhc4Do7ziNCXVJYD0rH
KDCq3boFhTlJ8bjNZM3asEXCKNj7ntSj/M62JXo4xTJqYuzR4J5f3CaZs+PaRbzZF9HU49or15jW
xI+/C805wyf786fVyfsWoncqqqHAXh4OsI0/unBFeFXkc87kMuhjldG8+dnb3Ee6v/iO9oqz8AZn
CEEJ2XZ9OAyeGkfOOCICRSPdcASZhduPyiE8AcLg3X47I0Igo17qX9eBaanBC8ZalJsEdoNVIBOq
a8QMHiH5ZO+lx09vyHRfl/GeaTlJgusD7M/5hM89u+eJ7CyRMWA6exSZYX1uxNEmylx/xfrRzFwR
YDoezzFLUpQeL7WhvyOUKwDUhuZ32vC0z2jAQdXTAuu90uykcfAUsY7CviSde0nfvUom//0x0l+A
G+GES7ZnXOcvEPYQ8t07VV1VIcRUm1lOe4EhEgMMppAh5iRDD5lwq7gs64gdiVdcSyq2XGLJQcRD
ZCoQYAjkb0bDToNSMaVLRqxiRKaBd4fAXNr1Jg0+b0IDMNfzaCS+TNhnfccG+amRrHRhSoqIjZe+
Rx57UW/gTpb0XMNmPz4bU8R4I9619oW3yeiUPzl/Wq0/gD1Uqwfuw7kq/dLc3hx08AzeY0q2p7sG
f+1BTrDv59wWG2gwuy/f7Qyvk5vCPAsm0oMnQKCtz1OgdpZRRaCQwUAEVw9TzaLtE0YuUwkpGzUN
/Gwxu6xZabDpPjfPmhQ81DwV4CffyaPywORJJya13AoRazZIBpvxPLoiPfp3L+A0HMEr0iO1bnz7
+vzX2Q3YjKf2DpChMiC4Q6sWxAGRwNIdGlYxvktziv9JMduJYgaAh+45YbLpUttcDm7brSXM2Gsk
5A0u719Zyq/E34ZDXnvoqQNYsE3/C03SSp4Iw7MTsWLn7gHTako2rl5erC14bDVmT3uktwT7lHtn
EI9/iH9U3knH9gdVMKBezJExRbIp42DtaLDHPmcLWWRhmFy5OKGK7gmh1IlsvEOhlOneM9M7bT0a
GX7UknU3Hj7Mbrfo9Zi8DR/RSVVBDg8kLyqmRxn9qsBK8s3cptep86AUqGGz8h/HaCILK71moCwY
5SY8k3hWkDjkdJ+xi/7au7bV+OcqD1HtAX25rHYfcUH+LoQlvDi9+WResixgEgsImm0MkXFqrsp0
BBJGmJxtyaAAXs39EPw87lwJ7JUNpOyOJwbU3I9UXXzQwlOlfm5ltnV/km45Zw32G/zFwP/zP2g1
xH6GokI2G2PLOyFMmUV87wSHdweXECmD2/PupqpuD5EgkO1MutLUMCnpHaDgxyNz1I2xj+ZkWaRo
lw1K+ygCehxT2BT2kM23eIM+rl98Pan7QFxL2gJAHVuxuvOG+kDQM78+PRtX8EiWtlVy2y3ezwwi
kJ+XJGJ5kjeAygLIrZW1hzInId76jIbotYV/v6YbBXyqon5l7GwC+c+vZmdtJ3CYDtAO3KqxndeX
BKS3eFC/3vikOC/FZWGtv9LdFHniyYCCN9Ybk168Nms/Y3wkl9UaHLHorjPRxdkMjB+8eqtKp5Io
oXFhXii+GPIgkfKZkT5Z0H9Lg7KnkrgVC+KVhWAZiVB3CeexqbHDdhqqGPHsun8EQtpXSS39wwYL
KCyqIfB3sg50aBqy2ACmEAnZIT8B3f7AQrAXirMki5e4J1zeSkKVjNG3wlyaCPn6x51lpr2EwOBb
6XJGq9uhvvwNmMZfFEEjnu//UTviBSYRiBsB/PSl0WVuzkYw71XXZzekwsp+TMYXoqRV+wExlXcG
EBsXSQ3JJtizhwOTx0j5Dm6hwUf5f1kai6vF+apzPgi6Ch0mznq0pjGZyVF9IHCJaPpuwN9+LC0+
Mqy9sp4Pvbn+DP8hHDJLnpGtJA+0N1GhGjJYDU9+jzlFWdswDThk4hyDz+7SflULnGDe4jQHhWKp
WtD09j4OZ0NjwzhY1+F8Gr5jRiT7pdJx0gGxUipPPaztDlQ4m5TqZ4XJySDfUhz+sD4WXEBG6W+X
t+wE5Ljl1jsq87NPiLx+ZMvpssdO7bdL0ENtAsNa1WqlHYqzwTDJrS1PfCjOepsuFVgjItF16YxA
o6ZYcncEmn4z8VU34iLE61V9f4coN4S43afzXlxuXXvPLSJIn9eKdXctq0fGUq53UIh5AQAjSwP5
RSY+anYp0W7DMzoPIMgTD5lJfa9UqJuSRfmWAMhylbiNphdaithOcPAch1O882YGtEoS/5ft5Ah0
6p9k/nExBBiHVihT/mF3EKlxSDO/T2bROUzxG4i6mWmR3ASKplpe/7EJ/tKEYEZLsco7NWBbtQHO
a2+vZx7rVhL5d7DnDKAV1zHMNmHp0yRlr5jlkNMLTmmEXlNmLG+jZAqJqTtPy4B3W2eM6C3mGS2E
v+n3a4v1j0n1xeuAH34oHL8/BIMeBvLb3tlc0X6Cu7BgqzThzcEWo0D5SQHIvOyjqmFGcJndaLs5
P0IPsVWvr1GtduhA7dAM1Ese/XKdrAOAvptJtnVOkrMS9BW+KH1tekfF9EF24BseyvVMnMGwTQ7F
MdmtHZ+OVRHXgZvfcqCMxbIVOXkIzlHGNPcQWT3tmVZ254UE8DRX1m5sYQ9Juguah6hR4uMCK58a
9/4GR0uZO+wNDHdxmohlovTZ8g5MMRlFHfT1764Q57aCNXyEi8ukf8J9jzahoJzhb1h4Ad8mlgfq
6SfrYRZkRJs/Pf4Xu/b29j5mfA8FWVmMuFsg6g8592gGyWmm6L4wVl+nogaiSe2XLaL4S1ibItIN
XGcbvh9T/8iiZcqQEzCYiVYD8gtjujhcKEWVuin/1ubi8if1qNELZSwV16dzHEqgfULE3oFkMB4l
nLjr+keN/lIvORmAkkVBUoJ+FbjdtKFyDBdFdqZFHYDWrzXahKfOZ7knMDM2Il7tzczK3ozbqdC5
pve7DCrVBBgI6EO0lyi6ASKEDYwS2wKf0BwFnWjXA7QUqMUS+ra2U+mKPryBvshW2GU37X4hYtQg
Jcx6DGDX0C6/qTtrfb2C15WcHDtzD5lJaTZZLqYgRPkkb/mJigVfE3V2PQzXErAQ8xXeOmybYQ/k
coucehxXFJuqZQ6YS/18kuGNk8RFNCqeZ8TBLsfSZKZf25ll0kBXwuz7S935yK/84kVE2N2aBCPI
gN3ruohe4bYl1FiSFXM0GVv9IwG/Sj9eG2ohrJRj/VKFAyHQR21WziW8h0BLsQ1pUn/lIhzYSn+R
wWHsbQ/3kfuuqiBTPtFJL/odgC474PZkvWlPv21TKlJEDIOzpdwHGrK1eZ96IN5D1nuXW8GBwgzr
Lpz9w05iYYXNyaELcDXyaoej/0WyT844DfsKFQu275hT1PNeXdTk4kMbGnoS1I1g6bd7+toa8m4p
v00YOsYgmkAii9FXlmY/nTp6aYpyQgoJhXONpj1uD9whp89VPNjYp5F7wwEpOp924D9XLcrwcfQr
y5NKD891WR+wM7cP7nmS7uLdj9C0k82MHDcqMoZmX8TcG4GiEiQ9NaD/vw7q2QQOGN1kdGN8GSZb
pqRSreRzj8PYXgMr+QcJ8KYt0cjMNQcm6em18o5iJQzi8aVBzPBcfIvkNREub4+hrbRBlwVf5uxb
qdh+Y7ugiczmkxa3xsO9DJyIbgV8/KhwI4TaNGuOl4rq7jlJiwVynAeLu/9Qo1riFpHPXRBY4QKh
5U8Xan3Z2VtwUIl8v2LC+tYvhdtAMCYEQaMkj3q//aMDPHCyDOkgFMkuHAfA6U06jeJGNY7ofP0T
FvPuKM5VdMeoPWtpojf2P9FTljml8NsdslgIJR1VpR9L7frkxr/nI8RHsUObNvtn9TTHDtPb9zaZ
ibJIguQaKz7hrUK6qyqLN36sjYy240oP0dtu8bWCFzzxRcfiwLuXPi2bYHb5WetiymqMQJhaopmW
hwEvaSWBRAasUj5wNM/yrOWqSUgq5aph5PcVAQQt/ryAQLT1ChJi25iZQ61u4cqS9jT9D71UKgVg
wZesLOrxxctMQ0Jn211IKRRRfJODr4gwXDYtjhIt0aGTFCJjaDNAnvpxczHqJUosCi5QDz/lfVg5
TN04gSAiHcbVSehRhIY29kUlFva1Vxs4mGw7SXV4rgmsjJEx+ZXZmsm3OLSZ5YNxja52v4+8/Clh
Ehl8Zn9q2QSh93eW3ONePbG+z+LPABS15F4ahSNaTfgVCJfLn3FiY0FkfFQInYRxA2yn7vM90iM1
G+ICmaTOFLxVWOzopn4UB2WJVWWdjPxGjpDCkALI9KE2X8iSJqBRIqzwrwbKvzO0zDhVLVpaUYYn
FHu5UrAaVytVIpiL9pS1gafJiAeZ+ddasJ+KAw39zHiI6mxDnqMiWRI5+8fHMeS8XJCBFtlDfLka
FA1d1bJwqhKJOX+1SaYskTp/Y60qrP/GRPi2jtGYtt5CdNvSwe95dShWgvj1iGeUqbd/WslMYtZV
6WNhjJzQr6MrfDIWB3FudblK+tjF2nGypr2pH4Q9g5LQHJCgcAFIgdTlyLw3KWlHghs6aGUZuo/N
J4U6ATO7YVfp5XQrSOtwUvcZhxfipcfefRruyqLpuPAe9gSzi6ORKjKkOHA69CtPDdgCm4G4Fr3f
ngbnL20sj9mqkNFZsP/iCpFxeR0NgmMAl4OhCLUcCZs2tc6C7qFQmf0WMHpB/BeKkdrAjjt4031A
YafKv/BlW2g5DGjKarZi1/Y/jRrxV15zLoT6j7P0Si0bkScyO2VqXXR0DXaUXsrP6Z2UZEbD0I0R
gEY7T/0Co1xANt4+b4f/8JpRquci6sN8pUeD+UYnaWougHcnEXOuZ/XJ6t9mevTkmO6C1OIZCQjr
sg2puxcN+Mu8jNfvbqvBYFQItNCF/EPDI7+tHPzw3QsEiNGdE/ozHsB91hZ1UFC6Qw5tQKHLcsOd
jvKjENClLz64Ky7URyDj12eN0+5/MwgDvmnb3n6SfMRJTRoLKQVu25+u1jsDvGitxdbWwnZDQwnX
4UN41UTuB3bA7cKCbl060YB0gm0MLx9b5/nYWToa7P5lprV87xY6QcgOwMKPUSWd+GEPqHfHPQYQ
KJKYbejubxgTSqOJLrOHCL9uAg34du0QUeI2lMrwGd4F1e+TGiv/EjPfT/cd458gs+jlUIht/0Y1
lYtjT1PjgF22gYS332VvXn2NGgN5eUx8sPHww0LT3otHGBmqevoOUf5rjTemhhHPCxVchgD+0+Gb
nIjrCBDeIrO8W3ikXd/AmLqIxfq6hKVBq/cu5fitItOAuqcPcoAYMtzP7T9ettKqDdSgjXU3IGh8
A1WJiuSOgHB85yYuNXep8PHv7Rnn5QqYFVx1cXw3nBiAzKcnq0k2Upyfw0rz9OLjItq+ZfAer3K4
gzlyXmJBl8jb0MvGwdO2sw0b5dMMumh/MUjJ+1md0vG7Uzjvv8JLozkgn3AIyvZkb4TBKs159N+4
GM29FD2TFLme2TeFtWRB+a1SztgB/LQ0u2MohURcHPpkpVsMJR3tDqSV680imkxXqp7K9oCwltqN
c6yWkkztgTHz1gC8V5bJEEI6P7raJ8UArGZYNcmEB3thALPkt9nZ7FkyX44Om7Qng2D3I8ZIs5mm
+Wws17fNuUDqIZj8/ZhDTMgWTlbh88Sv8o/5Jm6IcTXQaS9/49CNdGRmK21itvL4yN2mcdS7B0uz
sWoaYy9EmazqHN13eGTizl1TMW06/iNODUl0xfKoP3vFIiPPKj8+4c3xLkDwF4hTpxwkBzPBob0t
F8hFfXrCqefkmYK351F4zSso1jr/vCwfheNS5Eoh6lQMSjmMuwhV3A5BJjUfLhbSz1ofMJHSzHBY
MML87++I5vj4vLNE48bSnP66a9flWPlt6v6BYWV4ZcAwyBklOuHgJhjhTVJDs69sVr3bNANEfZx+
MiHYGGM3TfnUzp3UqA7sowWv++qbp3PBUOu77RP0a04sGQnWuptXzGSljBmaW5Bj2soHW80LNHOZ
VqZSswoG7y9Y41j8yQM6sa41TWLGu+OKrrOZmT5wijIqWqWHW2pYT00KCbKFZfOTkUBmZPcZ8+9M
IHfScP+Alp6KyfjAGACWWM06gdzBCl3nySZZG81LCN0emZr1WaMk45rnS+4KbhFn5sc7x6e1SgCu
+gyjRdDSqMY7eaQhdfDY6qIB1uaIus9V0WSh1j8jZPKy52YwBylVDOHOIJmfPFYVRjmkBNjC7taq
4OZUjMVouOEEZJ81OqoyauvRnOJ1NV/I80EaD9CVnXGgi/b7VrhbppbulnJaTw7sWH12pOi8DoZe
NxxGLH7xW1gwxdOb8QaNloxk2eRiIuYIWOuZjfI2U4wKOIe5Y+1NTtxqfNFvrPRqlfPagW/znP4F
+JyeCy7T5Fjiws70ehRB6QN5E9zV5Ugu+iol7AEzChuteYKZ/JPd7VPSy5zUoi61m5SKnhP3QQji
vr7bxkLhJNMAGgBjWTklDXy6FCEENE+Yq8mjwNJCoPjpVaFLJtR0sReQKfIcamAI4uG5isH8lDzp
pfitP0Lc+jgp5dlldzrcg+oTEkD9ElOYuU7RfCTh3bC0gToyb8MZ+zS/WrUtn72zgta7LhRbhyyd
5oStl6B0kQ82rmZ4tb0FhgbvIL6T6fgDVr139UQxvmzo1iE4cZu0sqOF4wVx24hXD1JKjtUlQujc
RnZrkIHonnhkTLrvaHZXhXLSp5HJFxMbBQl0toQ9gR0L98xed6Y5JwkEhYbucWp6wD2/1kAUNGrI
uBHMqGY/EWJqjmsdmn/m2RUxfjnVYntNAj8kKlFb76L7WNmQV8iCl1iL8J/6Fs3UmIXMSRev8RFr
L4KqhVo06CSynKoCL3MlMXed98igyJsQzh/tu1IqK0mRO2FY4zWd84xzxNYY6UYOzbJjHxEAIDKZ
6LHg1hCSYM39JC7DF/j6jTxGJTreNdtCLKAPgvY/T7w2ifqESgbRWqI7+eId+V2Odt5aUb3tI1EX
GIzS5wtocoU/pu/DwDS5KJHNvnunwVOJxU7VSET7b/p1UdlI1d4VCwQkt6YrxGIhnMAzF/7K8j4W
jkxApfWpiKF3yz+djuzMb6oU7M3bValbVLnsqNK7t/xb2RxZ+NMdmUGHJ6TjHUpUFIUXvI/zc1wl
MZtCKYX0SML4M3bYerl39Iv7awDux7F60moZOuHoK8gG2US99Qn3iyQflzY5W6auEM9d0YYafeKd
S/xJby6unsYHH9IJRvuhTblOs3JJiadP8EurOAvTgYotGuVeauFuenQE1wkBVQjqU2JLGQif0xsS
92CCxLRmjsZJZJLb9VhdBn8OxQq6rC/b2A7w55J1L226RfaJr9CnmGkcAIdjREA79h6AE9FQYio6
UspfjlgG8fKmHGhloewbkKCDqqGLDAwioGY2pQkf0nHLXAbaNZJmO5SkLAU4brrfCCQNZ2E22Tgx
UAtF3K9g53rEPdth/vAmNsXd6OKfm77SrADjILGLVsXjA9Q1IBfltf0tkW/fe7DCKerOETrMaNkX
MF/hBGMsFZ1gnHHiqqOT2wfDgvyhDKysm0gi9GgVXFZLsxM3aLMS/oo1R0HKpkBz3ceFIZNyrTpt
vMXMm++ko57jrgx+P2c3lHju+qHoiL5BwZfr8PsJdoXKdF2GYUaFXEbCb/BfdwNV07wcAlKah5E/
C6/MQzrny552woF2fKFKSG8jKtBtU9AULQTn0zwFXL3AgijuMkNdthBx82Na2euuIZdkgGQEoILl
bbt3NXWDCfdjgd1ISR0KwJbcwbne6ct7z3ne+pHYopTAA+DkIYQ6ihd14elChSRlHJw6Vs2arD+5
YoqMw2zOKqOZGdUASRJZfKYKrZaO0ww8CYh8wYeh0Y6t3i5tyUMcMBf5M92WH2MmLy7NTtBig0DB
+t3V5UWsbKNpEHsiIZLidvppRtaLI1aIAWH8dy88SbhRlmo2esxobAQ3rRTlw7B0+8gjUfIe5LRC
YRCrPzF8Oqf52X4WAcXqFLbEgxHhLeGtJCakWERwrG+60/9upmKfQ8GJ3D50HeK1oOGc3qhwlWQQ
uhRwmjmTCkPodEnDwYyMMJgwtcSA0WlfLB9nLpqQr85QnDI9j2FEojdjrznqasLWv8J5L65xG2sz
6qd6OgD2hegNK/bZ5eRYePsU8DeVmBYPrTlnnWfHaTZolaA6yRuLKkTdZtZ/neMn/GO1uyPnHFub
eiHDhvV80HZJlccixMfmGatJqK7Jn7H9M93oGveGSV9rRgqgHwVWMNEnEm4ovvqwZ7eFaLVHTZ2+
IHDD6zMjDa99y+YBL8sWnse4+M4/6bxVYQmXsduSnoS5PPt+IttkSdIBDIpNg+qJss0j1j1uLAIQ
y2GyCwarqMZfEA9fF/4kKgTX1XuebrQbPCLWuL6V87LRyrAfU16EXks5Azy9Z5yJ2e45r5tZ4IXv
U56UzAoS884sc1Gmu6Y5RVR/PRB3VrjSFvehCeZ+ruZjWVU2u4W/Sbk8NftkZnBUNmYyHC0YrSUo
TdQmhuQMb0M3U6QEfB021P3VJalJ/ISmNoCQF9LevXDC4NqjKKGddCdoWWl6aJC7WKAxabdI5Le5
wOzc3a7ld/osi68zg7F6DqEundHfyhHgzjctyNqkIsJk49Znlep3NSlIyKMyOxEURQb5woiN5LSc
W835nHopc8MkLNRePGu3VJXU4kr6Nrj+Br05k1KZbmwpfooR7qUjJ2QHJ4sKvbf26zT3BcKz5Ulx
JeljFRceMxaUUmIIPtZBxKfCdadqtFCAtnAQ9PZcYWrmLrL+kv9RFX/Ml7ueShCrBcejOf2jZY0B
Empr8Q4qvKCyabMpvUhQqZ1CAy/Q2nEWOPcU/PXbidgYxhUf8xGYBtpFrNRNb71i/HD8V9Gsw6hH
TSKaUt1lipa68v04a0DofX3vR7u11Z60lwPSBIvuOca4O4Z23O0g59FjUujYa/wyPIJRW3t2JJn+
pjGF1Y6Db1fJOKHMpsWo4zYBpECx7c3nqTIasIGzQXrrFWviC+84hkZLjg2g8Ot4y1aDY0wxu05k
QJ4h4hpK0WfMgWWxCJeRuPOhgteb/GcLg6QT4RlF+rK6YIkBnfjb3/VO8H76IEfI4jKRBuBniNse
2mA6SfPr1zzuVok/LdU+mCVPv9jgwZSnUdnZFMoJ+WIIf7U3Oui2oIrI/Jv+iru8zoRMuGqjOtgU
dEKySSTvZIEealK+nVDfk6JA9cryGJy7UFX9mKghUFreYVQS8paICB6TIXQkYwHfCCjNgZLBV7Qe
NeRlhypvh1KQS1l71Fj/nh1a+UWA0MTjFpAT5an+IUnZ9Z2ePDVOV7nhd7i1oiyQX4tg6Z2p66to
P7grYzGD71PL7eYE0ecPVwDjfIgY1e9q9/kzUD2I/U7oy0KyHWnE1Ijm4jkUiTpjz0f8D5TGdyBE
IztQ7gBdaYhNsV2zWEaQCEltl02Wr6hhXqxTonMIQ9CsuN6X97xz9mE1l+OKUG+EKPT+EDyP4D6U
c/KcP8YGNMuw87XgfR5CefMZfq+JeER7fQ7M6teIOW0KhtOcSqKKi7vWRiBMasmZTvPDORDsG4kj
B4budwOKKLC+JWxlYRh2unzG6lkCYaPtga0zsFtOANjJEgkxHnySKCF6+8NS387To9PLfdk740Ej
OfKPiFU/qEwpNm9tzH91gMpxI4PZrXzaa4Xx4+pEY2q9AXJRWz3QUItFJDAiYPPC49ZFMnmf2V8J
wYkWNaUpF1Z8NAaE4kkH+sjojEf1loX2fIPwLo3x3Gz0OCdaJiTC5zjdiIAUAIgGlYd+o/czciBs
vOCuXUun0yfOqYSvhONXbDD/utngSNHvlEVLTERvBHm2lylCuuEfhKBOaQv7tpO7ATgQcZs609eK
RDnTZqVkPxoLcLALWgtLSo+V9VuibpIwdElJz5siCg8cjhlnQ4rNyTAqx8hDWIq5mW4nvj9Ebpp5
JMPeq7EmdS2DsijJmq8yZ/bB+r5rgZprAne6B5AcK40R1T68N8es5+bzP4dFgIroa2fH7K4h4Xwc
KpFoPQG+KjuP9ens8kxnpYT+20zJQDjewGeWUagQ5S21uBgLXVOUA8E/ERYhcsIlkKS6gqRFih6T
nsN90x7sJQNQ1uXKQ8FlzFlGbSXjVI+NSDU5MvZW/gc+Uyr0zJJwzybQv4cNWsX0ShuZ1El+FlZF
lOzVH7R7JbonOiWcKb7EVcB0BI86GooHPTelQwRojgSaN24LGYop8jr7ryCnOSGVAc7KkkOmE90b
DqlSMFVRPy2oESNCBRci6DbaiUBI731wT5gzPo9OswtUwkVgKsTuXRJ2HGR58ZY1n8hrNDnTjZOF
Bb5k1ad4A8VLZbd0PxjI4fbrN4191VKr+cfxUnk07J0/ptZnocDz8vAnWlGw0gGD7Q2LU3PyEmtK
9lV1sqUTpGAGF1l+RudHbyAma4fiPq5/KaLIW71RwlPPbFyMPqPLTHwS5CPMXwtSW5ybMdCtQMGt
XfKn4oDn73JObKk6rP6IjLHo2N8iEq1424YZRiJP8uZ+KNANDsjDyXFqqikNH7GuQxB65XR8h0Dj
8pIa/IjMfZq1X5NUsI1nVMGpoS1usLvEe8HT1lqV/3tlY76UXvklA1gQC1dgfhj459p/dvhdafoE
JI4h04pApF2SiJlNA1OCza6yYGGJA3lqwWmz00elHRO7Gj+7Uny+qlUXI4Ubm4XpwheXVC+iavSl
z72oXSwenH2dSVmiBUMgS5kDbFQ5LUdZH3RP4WzdPrvENtntw2HYgXsAZVavruVQ0aVcNfrz4XdI
O6JZWwEk0H4U/6O9wfKQskikEr41/W70hgkxxFv2nrZ1+O8YJ/bPxNxkkrcy969Ap+r2VnK0rXYC
cqtFdeoQRgXAD9GBJtKKeGZ/G8VLVLSX0qe+39fMnWYQ4w6nW+NUI/L415FC5QlcaOBbIl0hQoxy
S3v8i5uw8x1aeCNjolLQdMVhJs7KzQX4ufQGS67xD+FMoTgy9K7cuJN/+kY46gPiyIqMtJ29sDzI
WF0Inxh67Xha39PwxXYZfWDFIzspCRit5LV3zQdo33J4tBtwg4iQI/LYl/smRKcG0gMXOV3KkOhz
b57y6Yk20bNtlUTkrOidSJS35Z+nHTqfCxapQq2qt3mkw4zvS/XqyW9plxkCn0ybMafMWu2APCzp
TCEa8GAfXhiZFENtR94fwsFwrLxciujPncLU57OI3YymfKfsntfPnm9FhLMHYrbmtii2auxghFLX
vCgtZjfG5MtYxF01YHqOilb8s+TcgFuXDE/RQUV2fP6RRhDiyBpeO8GziAsBWCmPOKl3xiDWa1RI
D8h8fsDhivhfCXWcOoK/bAZWSYWRfOkrZDGk46ekA40GgMD/+LUD9/wFoasksaxyIshGCjkihWGH
cVkSUUQ6yyGRwsqxiUQREdthP7xPHK6pRLFqqh70EasxD64slysNHLo1N25uVjxl12qA6A3MBMoc
2ICvN0w1uilmOmt+0T9Tis8d3RPJiCchYBaOmGZJdePO8UTWS88Y0v48HKy0nXy+tX2woWpg/VQd
hD9O0aheYCcz6kd66I0YWKWPy2lj1rhH9GwhHYy3gxahB5mirwa+qFEUO9BfVxAjgBcuwCgbzftv
UTGzvHGf71ImOwUysMUVDIN0xPbEadQJ/Om4KP9lYbT31kuA7sWy2ipFtuDbcwZak/JFrHZu57uH
eT084y0fcYwek47ieYF9kC4zPJB8rS5YYSgZisrwGZv8EyuzkzTF1CTBVpgJFow6Gv1b2PCd6ypN
gFhtbEVArJGcycTSXESDy/02zz+A2sDNmO4xGL3dqZf0dCc1/gIA8exN0LJqw6lyuw+z1Z5SuhUs
E9HHBmAM1OrkKhfPpp/btS0boWeh6mos8sxN6AiX0+PyETOFbqz2vOYjUcPk2CrL9LfkBykTVvWR
JHTXXTw5MU8i9zdzrdgaWolcK9F2WagZ+/7By+DhIgnPkEPPg37FN5Cfwn3YUydN2hNJogAeWEds
AUa7Y2aMt0Q6Sln4wsGyMcQe3NkjW3HUjQb46dCoHsw3AlvBGMjFgZKX32hMr5RaADmIsbsg1sGX
uaM3HJP3EnKmC6GAn5BFcevV2Hv+ddIOhJumlLBvFDSUR6IaZ00CdeIOk3k3+m7Xs5/fl0tuMRuK
feeOep763aseoECU18CXxYFlyfKrrO2T9QBB8wDWBtKq7a9mWcrqdO3iFEwVkfijMILVgg6+nnvv
Td8aZlFF1VgrRACKa8TakvrHd/Lvg+hjpcjRfHrnGILKIKvHkfTs6+sN3UqE1ksDmmQXySy6gN2v
wb7CJf4mhMiBY1VDahzLoZqzFwiHpN0pjeFv5GB8dPhB3eENu8xz7FWE0TY59OeVH7qatY44nAbx
jZ6stQpzmK7ryn/BMoMuQhU+aoWgizdQsme+kd3wRlyFw3sz7eYE1d53S1wPj4d4pmeqF3Rzi/GF
pyuEj5gbEx57tGpFmYHuMVxC/qWYg2DlTkrV/B17/PVy8pOR9i81dZSChiJORpMONsUrfKHImgXn
rgGoWnObTNJXZymzy+2H9qMYkcNYPGHfrlEG4DxEgHlMSbkJ6xd+TWEtKfd1s5t9c6LTkUAVXAhP
WA53mtIhaqGRlAJR46hHd0s+q5mn8WCv1pS41oso2ucxRxUU6YmfcvEEz4YC6cBOaIPdDCNuYNkI
JAm/rFWq8Tx4pjLC+0iT8y7WQujg6QzF0EKnwbducuY/cj6pI58hA04sMtBLi7j6VE9M1ulhXJFA
ftmKohoAgjlIspUiXpuMa2zWikZ5q/dE9lhbEhKX/Tt7uy2O1Wa2B+LclslWLxI4Q8q/ZtrUzK6T
wnnIpYnNEkkiFgZ/nDXeRFtrhVVr7vKBEHBuASql1vVgHrvl1MGF7Z9nH1SSbdO2xNqRQvru4vX4
Dd23i6weimTK9uPDA1p3/J1T0+xL6w1FLKMNI+kYYKewNKImyJdCz5hlRldHZqF4Kcp+NJeBge8+
y1cU2ZdGkTJffhJlqYoSFfa/Xv1/TMkoid5k5Esijsj14QKJDdZQoN1SM37cx1jX7qqZvMScOAEM
qoncVgZpTgwyga2gZX4UkOC8nqSTpswtYwSl0Mpa4gZRb26UPlinOLYGzzauSImlN0EAWh32Q37u
FkWw8IzkiVVJCAv+y3oMMoQtYfNmNizD+y2uGLxaO2kkt3LRhkyiq5yU3d5dMiJwFEW2pzddhJcm
MnIPbHZOU9MO0i6eduazZTqD0KBBr/YMhyuldh80tf/XmGox8A+8nWVoNpkbHhYoWDp7Opokbj8y
aEYb0AgA4Y/o1VDrbCZQCIrvRG3iMadrFzEYmeFlfeaswujQfi2QFavPVDIT1FfhvxYzupYr26cZ
pke4NMFzfGc3Bv7pMiy7aw3nzslItL96P8zfKCfydScdReiugak2ZNLftyiDncbzH5DQhVIIxwre
tSD2MOIdPegvuiTF1KL2Er61wgqGwHl85qKwbJMT0harYVCRiur+8eVSWQBoDk60bE5GTQybPGvL
C/SgP9+JG0liUEGW7xXuCoehWO9bXQpmVUY7gpb/3+nn6Ui+a3pv8mTD4bOBnar1M+gH+A/imQMP
IfKQzN4LX/nuUHr+H6MLiWjbSTj70PJGuueX/8S8Fljw1Wf2UPqP5jr5l5IDKTJ+C3/yWkDn6Tia
LNBBMN35QomdCsenmwq0rROFyOwRu/JdI5Et5jf0BHMOgAPp7+yJbd/R75xYyR00CfkLqDTemzuC
2hwoZASDWurYVhUD85ISmm+z1viu868wc2Aik8nFMOVvritE3y8BW5sU5e/iwUeKo+/yOBGfs+wv
pWIL8loG9ZXZDE1pdqVl1fXAkvfiZzZMOOGiZ0rrd/kTQNf/a6wBtlYbLMIpd12vKUtlgn5nl5K+
D0dFLI1c1drnL12U5WWSyc4VT+tvJlNa/N1aVdSCF0xahaSkq9DaBBwQ8URwiO9UwsP7fvHd7rdl
bGFvbnfefWd5gGc8AZ6I3IlSUk9I22MyQ0I9LtLxyKYe7ELfkVbwHxRHhaf2VrZTdUI5KFww+4k0
W8wuTOx3wssM7jee4ZjxZ9j2apDSpW1qrPey36YCqfZ5JbcQHNQAxpcANb+2OhLNyXlqATYacXve
1Oa/1zW2+2NzXWoa46F2DzOFPUlGZTbHVyNP7OqRaluRs1bMaDbm/mPC/3GbeRIVjtGz74iab/Fx
0woA7xJZeswKGLfhkZiPKbQsJ9gY9nhfRAQzZYuIZvWjl7O81Yl3fNx3DWfv88ENjijXlUAN8S5d
K0MCSCDPvIs2APIGcnHjxjcp0Wsj7hGyz9qBN85Ewgjs1YCpR36IP2eussAtTKmi4zyOyYA9+6WC
LAztnlp301Uy3escPiYoI/goJNp+C/a2sYxDZulckAsYDswDJLowKYOpexoUWmHkbC0A263Cj2UJ
yQ+v6eruJcNRoPpiC5PvdmNQ6ixOs6STVOPC8us4vUDWz+OgFMTAU5sHZrAXPP/EEQcf87zuaW7V
2zBKgxk6u44ixu8o6wSDvHSa4j8ukbasEtl3n180n3IcaXM/6IAUruc+RH7Zn/ob0Hf1dWM30S7Q
nNnHYrM5fV7qFL1XRDEQlhQam2RJMR8xBJOgm8Yq+5sKXLh4iKa56N2Kus2GclN7IaIVfssN1mty
eZvHX1VjfYMCm/RzZLyTAc2OLw4sWXEtL9r5AKH2Koqy0YEt49q91mE+UEFKy74JIPK8EJAXoB3V
vAtS7AHb2Npb+m01pkm7OvbUulnReBWUBBiHkStzA2ty3ku0H0s1sF40u9fZLbEzg7Eq7CC7JjSl
10zQUVWE2OOVIF9ormo3s5dKzB8wkLiV0TxbEpY1u028qbvu0vzTgu6agXdqCP3PMNnbvgIOjko2
alyou2vYDKxX51uV9mZtJsQh2ss3KH2OTKnEWDWAMVttJKuAMi/2jV7KNTijU0HUst+sHKiR1Vad
7s1rlFyS+rm+AdCNougklyKSwM0KKf7d2TZca0mrB35Z9rUKBBJPcV7m2pA50jPHYDhjv/Lm5chs
qcgfO9WCSSf2ahjhPvAz9sVLE2nnx4+K+mD1r8zCz52sDqLS8hQb8+yC1Atrc2gptr6trtRaNXHJ
NR4wJX6HaxOv1cprRDI+VvqJJgQ2VXBhiJhtCnI7hWteiGokCPOtVNhI1J4aWrh1zdXp0dCIFcFJ
khNahl3f57htc6+f7xH0j9K8ZJP4l9l0ED/Gmz7NdXHJfRe7MQUvJMqrDUXUj7skdYA0biabIC+E
X1CMfyA95lII8+dxUSmUq2SXlnUbKTvJDkh0+3LxjpObG7Xfzfw7eVLexI1/nv8sOXyf9Z/3GxED
FlmEIGTjBT6/aHEXZ6Codo9dTYx3aAO4A9wNsKXjmwW8z1ZhAIRzGkwTq3tkIUGvS4KoVFUdgqkR
wTrS94bVDs6h2E1Fx589H78iHbsUHTLC7mDgYOgelU2JnQ22LRpw+yi7LmE0vey9+2zmBjg7q689
xWrfxHNyOZViSb5vyA1Zj0scKQkhw3pstHDDzRjLLa85A/H3EDq4pMZ+NQbcwhPCWwACgPLGraot
eyve7CUvy9zFWSB2NPVb8rIT82cPzEzk53AOPZ605urExZl67gKhCFFhD7K9Qo2eTKUVark9abQD
rL7NM4nYnUSuE23Stbx+f8eIQYomnGse7N+bA0Kdz4dKqPJngN2hWcmQf9n/bAvzLFjCt3MjRIF7
uixAYUvA7Byu0O2vjy2Zc9MhDefVtVirbcddo9KC7FXaoSScEyCOguSE+tH4SFqhXIHAlh5OlLo/
EGGcck0iRaDLaRD6UuUoCDC6l+AE1yy2zanJS0l+2qWHh57facONSxdF3epHay06gWzuTmCYSY+T
ExO9ylEAG2BkVKSkSOe15J1tLMQ9eTZBkBvOrPxhscRbJQwTXZjX0nqyqnVXFkFyHjb9xO+72fNc
zyAQj8HJYfE2gKmHhvGGcOkRP0N01vFLOB/u2IcpeWFZkgMfPWemv1tYNmGgvUwYpgADDzpth6Ja
N+77M0pM37j7yJdAt/dM9kcVgYWOujBSWDPDV3X0Iqgoj+qr20P0/pTHg7WtQ7anTNjoPJT2AvD1
GvkgpyAtnEoKbTQdXRZGUAxB4cxE/s6C/4ys7vyFKQ1ikrxltqsWcm3LiJKTFTyAoMu3VMgDDb9d
uhgil4DdIXSIbTDA8Bcib/wzLMq9h6uAaD4/DUYQUcm531YAVZpgEQg7/Gfakk6SVDv7Eo1pxtpB
wYUJBNF/bPGG8iwmqrpdNIXg0cTO5JeU4WtZBviUDMWFmsTkItr0O8p0swBEFwLdFejoQw1dzn0m
glzfhf4jx6gLmsND1u/mkeMeH7xYKO8zj5kRGtDDMc7oRB4e5D9qRHOL+fx3VnvZ0fWiP5ERXAEI
yMNAlhcen+DKCGkP5nFoLVLeTUg9nFiaGUs0rj+kCmTXXaR97CKC7O/lNJK7rlrt4RXX112IOWGc
FLIcvi2spj9Ik2Zu1TMeGbn7KyeqbFqhkVrIeUR6U0OQc8rH3G7fkXlvibV6cd1NiY0v7CAlQeLa
HNedryVJXCKrZ39oVg6jiazZEv34MYnv/4QCFbAWJgOtF8ue0j6ds5lYOLukqofJUqp+iCWgZRqz
gPXsLbfpMmLUS281zjXgCpfWphwkzmpa3UuvIcLYP+VphPwzmI/GWce666yDZ31/SLb9IwsAscnq
isOywDUXPY2tRdeqqUzY9Wt1y2lPEbuhfpBJdIH7wBwV4TnmrmljyCTkN+zOtR+aTgVvgULiU9LR
OTJ/h1iO8r3SZ9Xs7sRQ7ICkX3O+rU5wdykd1Y4OesNvsJSb2882rmF8hsjAimIeUmozDCw7fSN7
9Q3RsdWgNmTWT5/1+Jfc4Egja5hX9Fv6CQsLz4UnyALbh18wM1t3Gm0M1ETWdsrS6v5BVX4VrpM1
HfmIVG2et5PIcDpnplNbNw7JNXfhMn9CRFjiOUfpAQoM8p1nx5mZ7oULo5yY05/GJsVlM1N3Cy3i
OZXWkK+TR+r5nowYLXASFopK7Noq2kkQXIhVOLNOp6gaIs//jd1zz7Ha/tavEsQ25GzT8lB1KyZM
mL0b24+Hd46QhTGqcPYxyxHWsS5igGxX9vx3qpwn9WDRX5lawE7RNIH4HaVQL7OeGt2JnDSOr4fT
bnj6dKFE7VXn/HrVYZXGPDNvjLeEZgGXIZ1XFznqMZkNysEUaJJYPAD5v5bFE2SekT/ZMgGyI1z4
nfBz3ddSNBnoYQ6tYKDhmTnY6ONBonv32OtpWSpgOhoLQ6ja3a7TKhOlzBFLNfzpB43lEcZBgP5z
3+HINchXttaynu4d5n1aV9W+W04QC6Bl9b/h415yPe5C4Fd61s3gSPAmy5hh6jLg9MRC4ydxoWne
YRJwKuCYWGFGeKCY8S4NMPUx+atN1yVdkjGGCk5vRolEL7YMlEO78sG2kNohRQWZ3ySidIV9kkZ/
B/KEoY6c/yDs3rYR+sk5rWxViqCVSiiZZQNodDbeKEFdFwM4ADgMxdxz0YBl8forBqt4xVMrqbDN
8ejaruRgZu/dk4pKn9uJGAFVhODPFJ59ooP/04DebgkHMG6NxdiWREaLsfjY/UA0z4OF+5SvEaAT
eNiX9grnATRzvPBiCVLGyZzfCwv6/FUbTsFzX0NbHKk7z4s7wIJ8nXGGriQOVgrCQFcVdSB7j8lK
z8A3TnSw+j/y6rzHhaO9B4o0jvzhfvKd6yuekuVOhT/P25VDXf4epXqzKdO+FZN/pAQrzggMyDCk
CnX04aceoJcyCVa3QzqSsUEuB9UNKzypss6fk5xqFDGZ20THnC2E94HmLS1x/yVhp/xGmzQ87z2m
VopDKLWlTUurzga4zz+Ue58zFiotDmyrxRxD4efmMuedVWJRPgVfHfmW7u7RrVLGul90DkA5DXZY
7Ux+5c7+GeCGUlAvQ2A2kDOxPtw0U7le2LnJja7kH1nfqbze6I2eGBZE2acUqcMQ4pxldqFxBbdD
MCdT5nIyHIN1DVFHVK11VWw3YauhByQOKXOfFZlcb9EyByEG7+gciCE+RWCxxYKg3a6sHrk0FUru
ZScW/ahEYiHp6HPt/gVRYeGcaVMGhffhE9qiHFX84WfLWfe6gljiLYQqp9faSd9DzXt5dRpXYurf
VlkT4rDehRpso0m40/ngjSi90vlIs/LoproPRZF01kKQNciPetDWonTLVMfMRDbpJWy2A1MTP6B2
9Ho5t9A41+fT1+LwWHvWz6CR+hTZvVnlTSdIvHwGdlTUD0l7r7IvBkt90t3dUbFlmWYaghgjOlm9
qZbEeEbbziXdd9SduH8MhE2T/S8spzAfsXTXxwuexBQJNo+6Zs3QV/HAxnfTzwvutSxqycs6Mq6k
7/dev9Iephct/wOrPPklJOgRVU0EafUvPMdrJee5jIHSgwHxUj5ljviRffS8uSvTm036h+rZZiCH
cSiWZEP3WYcgFXYjXcuC93bs0943x2U+ceeatAuac89fjrg0hqkTyWn0YYX7poQH2fkUsLoD8YwU
Nqe98GlCyMw++Ap7GCGXSxE7DJ0RBvDEajw++R5sF+kBkDfXacOUMpgW8NQvnc7dBQH7P+o7gHZM
Ew9Am1EZY5/nLK6scKSzvskeTj5E0vX0G1EAD3Sibq2LCppReIk6soPaw9CQdAYeIwjvTltX6eyr
DEDu+5W3g30U21QtI6hryOU7A1DTclxxgJaZy7g5YDRUJg5vm08I7iTc8Zyc7+Akz18STaEJr5ME
C00wmEHZVIW0cz7o0nGwVs3/xWlBvVGmZsznhczyeIINXjvCwXkfF+KjzSZ6IwXkROZcvTOKdRUw
qdb2gBgI4LG7bmfxfImFFnvIv7Bo7Ee8dUVj7HiyjG4HA3gBI2DoeShGxgDy7r20eUR0hVQH4h3o
XFkThg+WY7oIk0Gor3dBXZipwPvH8EEv8vixBEQYMHNcJu9GWFpzcIc2GdL1TTT3Pmlh6eWqkXRv
XRx4DpbdYUjhld03gS5MJQbJdwaztYZ3UhxV/b0w1tDmvcXcW2DbOP3gjgJAaL9nvf3n3XGd6Z4v
lUUxtRdwH5hlTGaz/xYrzjVbJ7i6Muuli8t2K8IDpd/D2DCN3gnU3yLoAybtZTVNsb1EowPR8Z0P
r70Hjm+vegHLKKeXDcPO+zC5QbEKlEe5rgJLTsuGEYc8hz9Ie15+VNeAnevUqIPj+j8Qt2+mQIy3
Q88BOxjBO5dsURcAQ9v9RaGz6d3GcPVTxO/H0ypBcPrWIGzAOu92B8sCDcKNr+8UjRvb+xWHmS6T
oYWVAiUhC/zjnci9krwTbNJNsUC0WgU6cGPshy/wrziOP3EzHH/Sb20d4rDIyMpmOY+ZuJczM/Ir
Mw3emCK1U7HMH+Tub+/XqSdR8UG5WkL+7M6yBxyUq0C8kpQgBfXRkua8MYgXu6drarTNZ7pCD66D
ZhtnldNGm8poHDCwxqjfCyjxx740uHPSbo0kJ6icJ6tDTr3rncEEseR46iETQq1DwBcNAH1MD9f2
kesYvf/37XHw7y6QKOHfjqPI+BbSeLE9IkX36tKbaT6+OZSDsPEagXTeXD4Lufj5FUdLKSFgC6kT
uE83/ydTuZXNJr1dNT1fZozU2l86CD5kljKJPBZ943fWeBS+fmijo+oJcL5LkqWKbD0a/+dpANzi
Odc4MWfFLIQb9faIT1w4oMWDQkynHGkxbsXHRmwa4QQIBMGD3/HzUEeMP2/qlVi+n/j0K/jk/NVq
EtKaWhX/GlzQqK3RYj+193KigcdfC9u3XxCuq6is3vXzSinDiCZhNOJvpWqJXOp8D3PukD4jXKSO
H6Al5gZcLYtKd7l+kvgpsSuVVRObozHYkD8Qm0Doz7QbIZhl/dKGoxnXDjkgH3dOtrn3PpcnxJTC
Cp4Qwv1Qkpo8DTLo793F1yLojbkB8JEwVKdH8Ik44xMxyJ1XX54axZij5k2iWZaUkb662xGc88fy
z/CGbIoQuFdQkDVf/mYHthslEFOnoVNxI4L7RcORvv+jV8M1kAXWTmcHPqfVzGEkhfF56AvdvdnR
EjFeuqBvJmd6F0Zk0w/KUdJYWF2VfYiZ1F60SEg4H20Up+YIJlc9lVMxfpF2qEsb/FQe74N11BKs
xFSWyHv63O+bX5mhSzmMtfTOy4PReMhBn2gddi0yZ2tqMzHZVfL4ud26p0X0j5CIsIZVJzYcVPbA
UGwCtARF1X5cccBo47Dq/QnRCB4HWgJKvY6bbVMk0iCvLiFQRsU1ndV3xmD7fbWHty5qCEIAMs3F
B6Z/MfqXvD+68BoiZmDG5taiyiJfu5kj+4H2FxYIhd9A2/HQa2ss5GqxBvV9sPIMCo3ZjwgJqAMy
XQFIqFv9bb7jXo+AWd2OhkVPOsHUSj6+xfuP9blh2VvxygZDodoAEa9U/ySxuh+FCCjgKQjYI9o4
vhRtE5w6I7P8dam6GOqUXtGKRgGq3R9/VLEKZV+MEdC7MpnuWn51LUyetnXl/ggMWO2KqvSc4jaW
ynMnWNAP18Nxez7Kw+0JWtwFuKK1gw4SOkVxEBks8FFMrFFq5TKnejSBavYatET51Qij/9LV9inX
ei6XTbFO1PmcWIjLQpD7lW/ZGCy1lzdxVJ0BAZN8BjBzcfVZ7B6/o5BTpaD+SH1KaDzRp7liGTF7
iWcJ0a5ztLiyyOAXwpt30vYWjCYfJSdd5W7WuQ/BOYUTeCU2qsgxaHgdS+1QZVRLzJ+9AvztRMYZ
0XaQY2kehG+wDVsgR1N50yqDaXcVrzzsRDdWeDNr5rtZyHL7ExbbZplfXuBQmALYZ22DhXS3a6qb
Mt6r00gwx8WzszF5sZTeUvfOCF5EVNEPjDTJie1ej0R6rMO83dQCscaQs0Jhcrdw9pvwgiyi5Efg
Do7mDaJLf9mwXPrEN1CcSN9SjAxPaqVxv8pkTdBongH7fGSUdsUpzxRl0l/g7z7GsaZFVZ/DhE/V
14Gc+eq0R62izEbQCLKK4MmquaSg4FilOeBpcGwbOe+V6PAxeDvDcJI2QaSDB7/8gxl7u5QmNPvA
QQw7ZjV1xuBQY0j7eY3ayi5wZzqAxgEjeelAzqcxGiCfxFdYBM1ja0zzrR8CnqCa5HwMKzftV9Fi
Eg3lW/xePjSZ+QnaK7dGZ2MAY52TZMm03ZX7SYxc3hq5uYrOVRSC3Ash8QYXNIlZDnZfVVIkLMxx
fgTOjQ2K8Ost9MJCzZiy0Azs0BAwQgzI8XvPFf1v/ToubX6XSaktJXijYE3Cy2qmhc4TFIplJXqd
+v+VeLbtsMTJZ3A2cYZQAr8kWP7ipdA8Tt7gW7V5+r42qcTuQdfrepitDm0kInrujoSnayn0EXI2
77U1QNZNLiCFn59D0GzwuyrEvRdfskm1KH285LYnCdOR6NSMmQPv60J4FpAa0DJGDksMbMfoDg2R
vtm4blNC55Dk1qBNb5j+ytolZRMIDGUTfwmpqhmEpS2hfuO6B4iNzZOWe0wdkJsKfBcXQUSiaf50
hyzFiPdOAJaM8LvounUeYl+8XY7NiPvK6yDijPaLuYZMlybkJho0Z1vgzIWFfrvYjWzmpRRHv1bL
zSNSPgA3hujDs77bjB/YGAX4DaXNOn/pfFfdF678/Auoj7tLkpCfs2dY1c/p4duE6BLlMQY3cEbO
5Bka95V/XjW7dwcMbRnz7FD2dIDihP3FKV7LVet4UM1js4m940rGvJgwlE/OM9RcOGGH3RDQXb6o
aZ8IoRrGYHyFsr97/GbxmsNCddtmmtrd0X14twRD4HJj9GwVMwz6Yl9zYwYAfOLYbiqIRMAzBTfL
Nz78p4Pew+MTtwBHEyfw3Hm42T12m5gcveW4zTrkksjyQ4IN/okaaFc/3YE35+nScvRwVjuiObg+
TJIStMi3Kha/Hggpm0/UVitLZ6M7xJLpbwcbMrBWFs5Qr7gW6/P5oL8e1CSrERpmvAyc4cTDNKWB
vtxqG8kfhJxcHmc4qIGazLvPq1fAkNEWFfTpwRln6cjDJSCFuR4CDOMuYAA/Vda5CAYZzoDRZlng
ZSWy3fWn8SbJEPrsuaZKeRjSW4oBIGyJRCbM+D9o0NPk4FcKPlrJQMYV0DkVaQiZlvjqeD6CeKmb
h308c/EARCwBAzl78qNBYQorM6zVwm+iJjicQvRBm9mivQ89E5uI2j6JcAKzMQ8btXMbmoiSjUKT
Sk3kJncY8/KFo+4X6aPNKXXfUh9CGpTfGcwL7hJ/s9IAGjXA9g8Lj4BDLbUNaM2kyxmM95RTmSPy
sNu5Vue9+e9WvQllVfgRSWA7Bd9/wMyCbc4C2Y/emLq62c9LpBgLEkfod5gBcA/pWqjRcn+vd2mm
NDXIZKPqcRdMc9qW40sxAZLCED4sfxyUEEgOMZeTABvuH9jNTTiv89U57tK7lnsFoPbG8ll6CkN6
hIYezST98T3bAMqUx6FLUjzZshg8JW8dRwOePaelhtxXhPcs3d40hFewv8aBvIQq9Q/DEcwwUnHg
WqoGuog8V8S+KJOTQ2CVpB24Hu7a4nqSXsmZBL/Sueympy2SO+9BzyCqRXr2KbZPXr9wjQBDpj73
fVxR0y7e7bCejxR8/N7FGL1Rqj4uEyANViXAZ3xq0mq+ka9hg9r6ZV46xBT5Q7wgo5HQFsCNSX1H
zC6Gou0V9yn2vDXyjyis9r2CpLAZ6oNacHtsK9Yu9cKjUu+QRElzDJNqruvq5lVrgiFrVBWdlqcs
RnSsRnuzwz0bd4xF3Q3jkEK2YYgsy2CUYKGSLxDMiVAZqUz/+5/n7OjLor42rnNALRem8+tSvn0z
XY3Su5rE563skENVgKFK/zEAWEfr9Nn7bmPMCyHbRD1LU7AfqJRQFLfA/NFVycOyx6jsCtswSnJW
IEHfIDUQMs7V2lC8Ii5uOfpALqBLVvEzrIhWJq9bEjd4mj6D8X4/Lg4eERiaI5vyqILqpwKZxLUK
IcErmI/T73ucGh7RTcxhMGaD/eObdWohEGqvJeNJJe+uDffTPh3BwPq1KEg1mlhJoKWywap8PADy
WHdRivYbs4s3lPH6nZtsvVUiqBsYar5gGFqVOq1Q/XKbGU5fnlDqRCVcju/RgU0TGrM/dgfqRLVr
PGm20XNV+jzy18L1ELrrcBWnx7wBsgAGZyv5Y/un03yuIGLj3WWzZTxVCMPXiTzCgg45Zv/tI9qM
eOudtAskpSlg6anXnDB1CHLIJkpxJ/MyGhwNPg9ERVbr1DUTGrg87wkZvJ3imT5DX+RG6Kr8yxy1
o9B6LBxWfRJ3d127vNoQWdQ5MtcpU3o5xIG/WXvMnD+UbEpA+uIdekskXANQmlH+ZJKwsoRFBTYQ
wlezTb6zR7LQuXf4pqCUyep/JaCJ4475cAchjNVr6AtT72XdtMVRCKN/QaVn+oOaWFWhgJDLeiSF
qlssJm34bNBGH0XokALeTn1kx9TyHZCjYZ2wsI4CIWMx0qAMdTczTGVoNEe1/5FJw3KzzsJ5UlAP
IRbv49myUPApnSu7BJGzwfK3hyO+vqDcStnqRZRONmnUgjW2f9WMh21KNCDRJY6gt8xqUfnwrPp+
XB37YUfmWFWn6WKKID0+8KioYTiwoHcomu8JN4PfKnGsvR1qwg3u0wqFP5vZwkLz9C6ubip+NDTg
ALna+qJ32rPkLp+JZm7le3qe3lC6lLEiEQzjUt3HCc4Zi7E5htRYueqOcgiPFipYRMtMhnSVNjjL
jmRbgjL2R+slvLKNQOypAguiCdx7X8RyMynvHRSovmUAxzULRBBuw3TifJBrZ+EBioqUbfpfHKSD
HA+gfhOhqo/APRNpCn+GT/KP1p9Sl9t01Suv1uU9OjUC9Cpmh+MaDDudc2j4/J6goadfDCbH67t/
0lVNatafev/bAx6knkaa/0Urd/17cZ/ake0FguYcxnngNYbcPkpBDTv4ZV6/lnIATjg7Edsli8T1
rFl+IwHv1jBbfMb8BWba78h4gUYXcnZo6DXWzHXrk2UKK9A45Y295LbDOwJtg4pcHtw8M/Cnmx7E
Bf2flQamImSRIHpe+IpKhmfXo+tEfMAIqZ2zLjOq724Fxrug8ao57sAZ3RUj7iYXttr0k1Pb9YO4
3khXajT3ryKGmKg6WJ2Bvv3nGh5CZUd5zYWXS71q1+C7epNYF+wmt8ZKLyKLmrWHS2lP/sKOFaho
67aWOu2IjvrXLylm0ARLmLv3DZcDb0Ocskm6QENgKyU34miaoZ9tPHf7X0rNFw2Gg1Mti/DsHta1
JoTbnpmhffDVebhxojvIgvdWH6+o3ZqYHVZXspYonRbUXEccnHVmSOimJm7MBCF5FkTNZB19foWi
HMxRqJx/Slxvaf8uozCWmD8saqdyJyEENcn78FJ3GzCrj6sxC/szY01PupEN9b3hQx359SKBQ+m1
HXzVKAnNgOTOgkSo1UGuYFuJ56oExlftU3ohi/fi7wxRaM/fXnLuQ+l6mfihw6/4QRb7fnN5oqbX
obiBFC0SVtdUzqj1f7MPeGpfyoKpPuHnzLN01MdLgCZmryp04MlgCtNRx+W7uXL4iFIlihbukpPQ
m+z33JnJgEcwMH3vStzzzAdH2r/eXl2fx0n2Fkzn9KbuROkEQ/3zEVBNmUUyglF4w/NKV+RHZ/a0
AQzcz/vBgBfzzGozlnh+KHntCU74M6sn16rKs7GnDjUo/ahm1t240CPvTPxJ8uvM4vqAEFQjHGBj
mwA+bTGQ/2dSt0VAGmZM7BQ8S/tINYA3waYZgcmdgZymqv1TOzhxb4hxfBJBfKlGwKasLmmNDlgs
jZtL5MhGo7XmVzGEqN2o3AYlF3fBsrxVzNSA3t48946DmEN+YPlzFmqX7aIGwIY+egvyN5iBYUNn
jTwwin8tBQVXMEMATz8ZQZbQpqV7B4H5cD83XIzg+jweoJCdt6heCQ40Y7E7V7OTFV2DukT58YN8
1zbwm/OIrsCG6pHjkKE5is04+RfK1iCygtoVr3P8PHzS4+pY9vcYQ1eOS8yk8Xab6xcX34S1QdDG
9J11iPc6kMaPMLZIQQDFBIxOmHlce54cayDrOx6qIt0Oe6rVt3CrKaIut9fUvO5KDCNtEHDbenKr
SolvD6PWF07HqBhTtkHpR4ZqN2p9pamSqc1UjgmucBrM6JnaMRHiV1qbc1DCBbftRnDxgwMBB+23
+OwvhvBqEtHaWv9+Oc/5mBFXaYHDehn8PeGhBfkmx3K8EFOi5XqtQoHneqo0pYZv402+kyEhKc0/
pAmqMTSwr9RoqnfF/LAgwFA++vQ+6IfDKdkaBbXvRFUaBlrlT9na0UEByQxKyHoW60WBJjimdHQJ
IsdjCMIb+ueyPOlUnxtFPyfTxX0mka5j7UNt2bKlnNa0L09Tiqd6u8N189cCoUCIlP+pF/kMU7dZ
rZ5E1chnI/irA+hRXnBZ/J35Oemc8+BCg+kOy/FQmYzMszeU/TiixcOZi44wi2R+GaMQRhJrNOSM
BQkSQYza1Jr3d1b+eOux0ppk44ZKQELlayhvH0GAPT0BR9a4Khl7+aqjRDBrUEM5oDjrMNi5qgeM
8Kd6hyAETm2JNnOE8cGJUbtxOL94oFDUFJzyoqkpTCgY7nWzIX7cFhVuwGzh3lrI6deOeBdX7x4A
yfIqNUOcrYRgTgGopKor1IoJdAYTewzaI6YY+gx6S6EUaUuP0htuqwxA9bkIWuStJ2fszvHW+emu
c8jsBZVaxjgYpq/m/k8k11Iw2waiGwG11Z9uyP0RytpVYrZrtHTPY8QlXNn8qecgSkBzASXMrwpU
2BQmQtuT1bhuKMgFwWEES0LraB7WzpRcNwa/JntuKO/8zQtvjFSVQg0IaLCMuue9kPfZktNIyklQ
kbuI+RrDKno5ZvluHdWORM/ig4XQnxRFXq0CZ1wQJ1/J8Xf+p9a36bikMz8iBey6gqh0wps02z7n
u9/6qR5OS0I1RC9FfBJ1+7DO7WF9DqTurs7rQH5fsQEZemMm98Fpwv3IUgKnbh1xhgFWtvKNMZ1Z
XIGp7Ukgwla6JbPXPwUuInbJYeaF/jL3TEkzNVxaWQIQ8DPlAJ7V64K2Er3aBPmTBiJvbmHfKH0Z
lJS0ruccHta+De+Zza0HtPE1bl1VePGivV1t2fgAkMb5IWKBLBVSCDXrG0ZO4f5qqgnw0Q7xbsSK
1naMhUmztEqc67PF8KhQn2i5zD7D2DnoUmye4zkk1M/dfKyW49j67h5GfBXM8fUgKxQ6tFsEeRen
upmbPt1uTUV9tVvhxCki81JmgxeInz1GtjmJGP9HBWF0Ev2u7aPOjLtb7j5EeOoamPj4i1MaYQzj
VfKOM8lRBeUdjL7NZh3Dvi47J1mFwRaHVEEXRjvTuXIJO1mVGZF4wbeLE7tRM4mF5nc2z9EMZmEr
N0W8d/K+Qc1ck6jD5RHhk+gjjtcv7LFoFvkUL6CHgaIQTKJT/B4u5GY6v8NS3tTRh0dP47LrLHiH
fsDYQCklPWXz8Jr7KF+WumX536RtD3BJG+ySY7itfGyW9zN547bM0k/OGnLGm8QCTOhlwRn516Sj
aJfJq72lvkflzjdbRHBHJxDsx1AuOvrfBbIdU3GY7EzSdagUfjmDiY3l8CFjJo/dvqo9wQi4H8Te
rS0fSZlHR6bJs8WL8Hssi2TwE4kDlfWaLN03zx8puh1MhoTBYaCI60PFXdYCgRBEag1hmmcHp8zG
ejv66+tYnNHB1ZT5dyFbwwxs0yxvYhR/gI6TxCEXVTSjF3jiKQPydVY78S0Dc0LgqUhSj/kPDOo+
18u8RtINZo7/udmZa8jDCXPNXvuRzzUwStNeDYb1sl3S+nXHIBNRnv6LWvsNOHecdtNQ9AyOHR6n
yIfuDW+Lv3ig6cXSjtqdAjYQmFfSnjnvNJJkH+uFdzP5iAiRvL7GutRDGD7fKLdpzvIu3pNS3Pb7
DophzwZXvaWqAhq/WCpWRJmdQJPZo91Kjuay8J5BKOylXaGsjziRabGErWI1FlfV4nkjooMxa22R
RYTq3UcD3gJccjack0lxQtYetr/khpZOLzqc1elootgBL6RNVMZtRGGBZZANYEzYQGlnyf20waBY
dvBZI8H/zCdWNVGw30Yrrbjs5PWVPsQ4twz4RBz8ZcVClVoFje+wIOJjfFkpX1jmTkmDDM7Xgas9
q5xv+cLZ9F0R6nATqpIm89krD9VX1DPv16WfM8r0e7cjP2ONx8KiMg1lXrm4mMMDCKxAh8rVaxQ8
5k+938m6T4vOykYo7Ci4kFiKdoDUhWDgwqbHq2BOOVaEw2TYrX2bELDotQHHDzAkH45aL3lXGBp6
etWGB0L7V8P9tC4XX0YlKioBmfDiIznX1M3ERIXwyIJPUB/J6L6avgRbUL5AKscvJZVZ9HNFnSP+
M6F4r/WtcA/dpemuwFHGPB/TYyK5mhJcQ/5BBcTALAiGz9PH/EA+Rl+vCThzKLA83Zac5EwpgT1D
4ucEA/JjrEeQ0CYQ4w/IeTqiWpav2r419GSduvfCsVbv+B/wcOttZaClcBv4lW60Qhmo223beQCA
xxsQKnS6eaoGbErTIULxsym5BNR687J8+ZRJOZn2OkcdeVP4GEw2uZUl7GQtKhLMqffXhVS6ym90
THke+fax+Byf9Fyo613t7jFwwQKfjsH9QmZU8RLcoM3OJpbybyq6lktZBpalug+FnEbsfTPanhcf
7FcCpXwbmr4agVJfcLtxIViQlHUMiyj880FYF8pF3sUUo5WEMORdm+ptKLJGxh/rIS9rnMVtEmiK
hfLnDW5uHRLuIWcFdzqyz/VXcZMOLKUoKPb6BRdrSQAyiAycvM7b2nMB8GIxIA2vpXXhQvMdg1cw
YSmHez7jyNi3x90VMYh47k7I+4xKYN8YPwSiReypypfwhHXNuvTWqWRtESd2QR6iVa+9ZPp7SMof
f6HTfxQ1reirWR3W0pGcmi16cnCkHVXNwTjOujUzwixFLbxvyUrenoKnSUkyBmyeNaUQrqOw27co
yXN8cObTDHyIz3LSwopk8ywx4P2/TYEt/fPLf+AaUjLT1MBhRt9HpRUtF4Slc0FENnerMzBaaWqI
R+GH/E08S63P11ePlphlBMo5lQjD2IAz4fX46qu7L1BmcM+R6rBcRF7pbROjri3xVOMy7QwJU5iu
J60SWMruABXOp0cfND/V5kN/9YltXQ3KgKIa9w2mFa8gvNS6YN9afuRd96OLNCs51vn8ST9p+0DG
hKVz9nhrJLlpZyxPhI6iLAZWj6+eM4bb8sstJM7uC0w5q2tccyryEDwzkOcOPUmzdCt0AZeD79WE
J0Z+0id3Yosuqy7UX3908Lk31mz2mGroeBCYH0I/wwyBhbFYlRH6pqTcXdCSiOJdS086kEN2vi2K
sFqrlHauN33XGDu4y/aPNqGu5df1iDU6eNpfKQWtZqjCsL9T//I3peFOSA9ONJG46TpC2i0mlJ1+
NfXbhkLZaMjSSct1FtdLyUgGozb9T3IoXyVi6Zhkn+NwV5PPcfjIVg8fJirhlB0EeTOXPRm45wt+
JO7+9gdCW9nk/PNqyPHslH02NeY8waxLLvqZIi+Um1Fl3+zRLGxzSAQUJ690rVxPzEcFcZD+dCOC
M5nIkYZILHpONQgXA8fHDB0QxUhoC8wfCPP6b9HC0V9CyOtFpC7XZ/ivSA7SSl/N/9oGcCtAkjrq
MoGbCD4UlnBDhhPfgYD1fwTPAWPI9lJ3Q7Jr4QUWlsYnjj94r1tdKNbWNUpR98QHEZcG0LVEPKE4
ceufaQZCjMRNuyXFr5jtGmpbq9sIXXDt4rTEiNM7y7zgOXPFn/A2zI11VneTr1+6itbNbdaf5hih
eSHH/SKLAGIx6tKZbgyKNp3wb0+iwbw1dchKsMQWw2Y/flXj6duWIhoqqVvChB0pU70ul9Q2oaPY
mdFf6c7TA4Pp//E7+bPCg0qjbjA0LdIb/1919oUNZJy7WXGXhA8r7lxBXv8A4uXkgZvqyAuVJaKU
CaW/eNtrE3G1fBPlaJafaM1R/pqcDp8rFoCF2uaKFiVj6teTSmBYK6Pz5fCJF5EGGcSV20bxW/IN
G+OU/rN+5mBGF1VAI4pfDF+l5bVntqFBMXib/NDt7pdAz6NNbUcKmP9STeqsDDopzzQtXsN+5by9
C0Yz0/hX9PYBU0a5QQjYcp5dm6jpdTHFTI6eZrM8AksN8UTbejYjC9KUyXCJ3GdF1aiApBiX0Whp
y6RsPAI56WVTqVG2Zm2tglNmRTLOk4hlOHS8L84vTSEosOZqRx8pB+vT8Q68nHUNvYWnsSfWlqeE
gYHme1ehVdzEZ1RwBUdlLLxKI00qK3EN4m4RO+uViCLY6xrNtvnsT7mbr8gCe2qiW/hq5T1b3wL3
G4NqR+TZ6wvovV7W3Jpq5i8jNG/5nLD3wqeofpVzndI7INaksOh3TdNXjtGgbuJ3+xHB6UD0jAsi
pQXJn/7xNDuNHZv8Qwsmoqzs062cu5ahV8CKaqu9YKbDM3lklSfuK/760IVZ3YIKLcFG49i10A7S
S06ll5LXWUEbT4YnWSntlf9W1QtiyTjW7gvkj37klKqjxrw26edzR+VjkeqXqooLiacdzX+9K9O7
F5rD2OaGk2hXWfTFu0B72CyyjTk2iCRgI4kMaS8kS6BAoDFtofjq34Ty71+BqscIU2e9zH6Qbk+j
vZhJ2gxAZgZtNTXlpMVyYSxZcK6sjfmf3rvpxbRgGTqAL8Q2Iex112MCMWmyj+w+pkoneIVxlCXI
mjQyvwP9vtSsCkRNFXoszzRsv/Ls631Bdv8iI1iXA+W1hq8EV+lfIyQULIElGoJABa9puD2MVWYU
npCaNwbYoPeeyNkQedEN2J4R7AOHymDuLFw6GovdirIIzfp/RCUrnfqHNjTVxmcwYEN5s1ssTbyn
6Vfpq/UhJX2Sc0FQQAlC2m6CmvIGmDuG6b3LnDr31KmeccyGxeg5u6tziClZ3UWeNDtbIOosgUrE
1zgYDexKKf1/zAmp3ytgOsDWMpIX4n79/6Yn+XKzl07sEmwnyvh0ONfbGFH5dK44k/w++iBpGD92
Ah56gka7p2aER8DeViULqZtoJH5/c7hv0ZQf8Eg9oFvVspqOq8XSQ2kc+EtbZSm7baXMV9TNiHPH
E7XV25yjq1Jpj4fzkJS5sd1vZd6hXlQz1yCdti07sDGaZUwwJExgdWNrwpZSmsmiueggtQUrk1dJ
TBIXVxzB13hUilREOW9ch6qNxtu4MbtpimtBUyBgsjNMGEDgcxTEv6Zhq6OYFagmmxK+NJMOje4q
TiwNibGCntASOoN7uhHx/oz6NurZpyivkcbnOebOs7KJXRApV/v6uIZWzOrcYRztZTVbAsSbHO8K
2kFCa/M+806XDj+QKXOkNTcVfZeE0cJ3f958JYMXo7antWWgn9OR+Py8qv9lxY6SevObHz4fYXqK
qsROlPcvKyqR0Xxv0KlfNWyUE4q/J9dIHLHx1gXI81C7PoY5kMaDsySXhqD8rsGe2NGQ615WK2IU
2/o7bsOp5k6bzBzG78FHZzbme6oN94Qi44LEM8+lTnh/94TWG7Qz8qJ4j1UgnpFOXYklAb2ujhoK
ft2TsrNc5ESF7Mc7ASdyJq8X+a4f+nKd6o6x+B14Bzdrua29pK9dYyVb8KZZI57EWAn0Pu+AUd2L
MSXg15EKNBOr8zPv9g+4OOrgDUGwxKjzHIhEgS4f2k/syMLfBCfjPiZLrr62iRPd+dKHEn39e/N5
Pkb8x/RDUPpuredOAdbpmrOhBIwOMN5jHHbDGQq3vVDBHsJBQD9qQ69CV88QjgNx8rpsPu5IqPoX
1IBCf71wCCLA6Rg9X24siaQpVUO6llOU87JCtsEyQVHnE0QOW2r164kkajAuu28ZlnSPsiEfr7n7
u1tCQgSdS+V02bn1RiWMoy8r71bzfJEfb3/8dFLcwh4Vs9FH+AAakPcSKaV4jOWZtoySW4FtHhng
T3ERF+mfVoZxAC/f0K0rhgj2jXy8vXIhoBbfH8aPQfG5g3N7tPvo1sbzOtow4HcdBZ2y1ctbr2vz
CNfEojNRONtpokARbOj27fCnwVcTr78aCL0x+tBbdPfDhh7be14C5K/H2yuXcQseeZgRbAysvDeM
CesxJKIl3HcdGKyNfCY0IEwWk1JkYBv4E9oCESMqbx9CbqCbhccUvGdGwg8Wo8/7yPauDsbRRdFM
R8E+skfyK43c1rGHli/S05SaxcVw2k0vKzATLyWK5m0Rci1LWJUu+aLV3T7HJAFXOv8Dt7y6Y/fe
3JRbw24q15jTL1d+5kxv5tJehzMex627Y0fcdpsifVNzl9wJHrfL0PR5r+I7Z39GKtLP2o93ANS2
SedNUDo54e0rMeFVfyrPnLNBCRKA/efsaKhAR1sUZ3oGKA7kEZDcuv1tF6/GhC5wZ3ZW9baxgDge
gVSIYQjX11MWLuseXdLVQZ9R3UEwaAvvZD7cS+2gGURR3QnT5zz8wYXfgLjTy2Kh+zV5VdFW9QSE
Y8uUUyCnyWdpotNCNsPnkcMLLwPSIj+tmECGHQVfN4qN4gNBDHNzk3C1TqMXEe43WVd/xS+tOUpr
nemNOrZWHlsvNSCwudyu6/dLAdheXQain8mrS90jiurKFJB5FMii/meZL5DNpjilV/91EQAEh//+
Ds1WhCzU5V8tKwWE17314L8Xk5g8NbYRC/PJPmmdC+hD/65ofCv1bquT/r0VqabovoQmLFHu1Uf9
VeH+GrgBryXNuJXKnPSI7RmtdBOQGqbGA/DC1YQVofSEgksOAShqCtD9Xu2IyATRGJLFh5vBLLqB
h1ehqOzVAE1R9Bx2b362MYAiKhjEy8Sw8W1CNP8FbVRBZ5zVyaZQr414vY3VO0ISmQnnbgEKkMaR
v++BIwK47zBDvafiFzb4CNX//NhGTPHH6gGmI9V5lT8fDqqhc3JXOlPZYigIQ7sJ/LF0Zg6uNDbm
gB4s63jU4RUdCuooGPKiUeUBnqW9jj2gLqJo7yGW06hbPuzVcePmhteaEE+OMvJ1FDLmUMZVD/Uf
bgo88UlulKj2xg56XWme30kwJiDPsSoaxuUUJbPDXZ9TcgvEVjh5dTTmE9LQAaN6lB0FNfs/1dHL
isqdmAX8gKL4OSRmQ4hOrImB80Zg9IM7PfuH1XN62iNvZX9FwoCyH3okSdrV1/f/1Q84olKWfi2D
gnZk8eoXQjLwUPcXGkPK5O1qTgfu3343Ht2t3TlR254M18IpkJCS0nQHY+D9hGy/nxFwFo9RsgZX
EtHc3RV6CivGMxhAzmW0RexAHWjOlWVbcsoD+Mj8ShC+SqnUhwij20AX3U4nLnuiAO/+7Dfh3pCN
uu3GuzH9OVzIebapVEBxAWEqrEB0oe6WRn2W0zPP/LlrjfSx5idF7ejWepBFhNhJVGcGhOtccrps
hJvz/TDYNFWhBVwafW0CxEZyM4fzpqXREeAQ9QG7iuSkoxC9SsD0NVYTUrAed3RCrZcTo49xKBd5
a297EwK1htUNcvyyVjMWmakMI4Wvw9Uzgh6NNXJQuNBXvAHanta0n4cDhzsuQVnM0qu93sfo0dZG
y6maLvrv+23QJJa/1A9GocpDQqPFcWsrjCTRN9eFe1Dbf+rgcZNBdwrrS7U8fxHmEn3cdCcbg19P
l23gQFPFFY9QLVfpSRpc33Tg9KVaCr3k8JaA9iucx8rrdITYmSbqLqnAoMwfPzk6zWPy1OvrwM53
HJBauvnqfr3kvDR/1rSkeYn6I0YmZmEoWjtE5eNLMWW4NRBx06nWtuGIf2As+30esHXbjcE10tnk
BtW42W3u0rB/FNZhCjDYiqw3XPnZn2fGnRUxFiuNob1iM/Gh5PlhMZGvIBFH2l3iWvAVnh/2u1ZQ
MfGVj4dzTIWpDrNnDOs+KBSgJBjVbUaouzMWBdkFcys36C8Gt4Z4Xptcc7uWIMgOe0kxCVCvZlLU
EoRCb/T8ZMKoXiugfhkEYjZ9A7wJE6hP2jGlnl+5/ldP50tReirErd4iPFkMBa4CjLr+O3c9RMsy
RrkN79qQPnmBrpPU9A363h8mncttX4Dr+gFOtVetwChkA54oQfDVEbJc1qq/4Cw4U9KTvD2yYtzY
vuc4Q3McR98Kjke/H2tbNe1zbpX0UJNiWkauTQ0+yVWTjELzL0bRsqu97fn4MTvCcd0Qg/vfCEbr
cNhOoFBcuMleW/EllAT4HkhNJ+7Dp1jktrEzxX2q7aZU6p5Ni1TJ45wqsEpbD8Ha5JbYZM+9FcFR
nndh5YYkWvXJvPnzZKmbfCQ2KVmC5qQf/TOVLo8B5GCB6CFg/oNaJvc0VGwh5K0umVA4HZgLTctV
4VNxOUSqwuPosLXPH07LnodnvaRDOLs0XF398dY2q2Vdd8ZAqJTActKVcInbSIh7gZ5QZ6anasdx
JlKVNWnWqRCtdRfe36hzK2jG5c+aFGiVfSiKjE+Rzn6zIwTl37VpXq0N4SEV6PGEmOnuZ+rY2l66
4uQrLXBBXFvUnglpbsWD+lcSvEtBYruGx5y1c+kxfJU/o5kVn2kp+jphJ/e/Suo3nre14EmNj8Se
xN2MhtcsP7+1YQln3RNi9Wv9AZqH+O58pC8B2hZEnxGvvZiRzHke/I9W6yIujmyABs/oSnRp6l3A
5kscERSjlpb+eMX0F8kI9/A8O91dPFUZ++qqwjQMaDc1ktOiKcXq4C4Rl9JS2aoyZJeGoREHU2Mg
xSvVudUpaBaKhRznMANEvMSDNX9cWzQc0QDc/vJKRbYRG0dRo/h9Hd0a2s/zwh89GCYqJlDc8nID
GY8Icwqsr3z9aYTtu7HEordmI5pkD6HM4jKjmzzFB8aWGPggI4FQxfrC7GFjQuJe1s04PFjEcv67
g3/OCW0BYgGKmTgQDhwk1bsQTJEaL84ZL4af6LWcTdFMrmYptfme/+s0hbvzvbZVEGxJErkP4+hc
EyL8boZTzuB66jySuCPEUiDJgqragH/a5DebX/QV8zi2gzCS+H6HS74jVRL3dIOgEgw+Ibs3hgli
Zq+36QVW7AqXxAQdvyjVOt56wcbRYykU0y0YSlr+1qlnzNMVZJeF6xy1uFNqO0L29zhZ0+GZSlJO
dcMfyRIkEMMdnAlh6WMJgQ/KhXgLGSIqc3jBUYDMzLnpwUf6TjBC5T1kRyMcdUUoof0yfIrZxr5z
eNhhKntJIq/YWGd7EsdjqtbHiusRVfUUbZOZ3VUSGw0m3xWREz37XuS5AwvXSuZ6awF7vREEko2K
nXD5dziUKB7I9hB9zHaf5PcRcd5YwckBemFe2Rb0vEgyupMvnnrC/+c9NTHmC/MCn8ASZoHOjQS8
rVLmMqIPh4i+H3UVJuiyLM/yYRchNa/hW+fhQwrr3hKjV1aZ8hxraZiWO+Qovux08BRtvs2HKTNg
jGlMlm2YnqRdSpg4y+dkOP0tSuUpJReZuQd/Ne5ZxONvabCdGxOWSRdrXTR7P1Twk6q+e8xQWsRL
cUHmivxDtvKnY2+QDBeSRIWTG/LqZeFNf4m6HDe5vGhui7VtgDSPZ57YqgiLTwRkPYnhdSLMNB40
4FH9jKtg51CUczS3vmMKQRNzVVzmemv4a46Bbx4nE4AIcf/OEW8+jlG8qMU3UJRvliEw2rrjAv4P
XXhTfYUGgErJO41C9OsXaOSqboFvXwerC93iYyZ6p5izT7jwhJMksApF+WlVFPOKbSqLmPwbGtbp
UTWKgHu6akddfpP7qvsViaEpLuhSVejgZBSqE+CksxNl7Nu/3xEmJPT5lZuoJJh/h6bHODwgWxw8
RZz8I3opZUTBaD2ptItTQKcQwDSqapX5X7gR21C1k9fbNKAvhC6fIipE0QiAY2Rwh2MxmDT5B+Xy
tAk0+fNx8T7FtH81VBUkpfHkmIsriu3loOYjGhv1r7uxkqqnzX66B3qqO4TAfwpcDv4cDXaKiKXD
Vur6SSur9HKsfQ0QSHyIIk8jyqoSfMdpbb7zNTzXgf1Rd03aWZODoaVTTrtryk1y80iN1UWY1/i2
0LqAukcBhhMh5xEpyNwP4w1bHKdqwEnNc/PTKpv6+N5L0iMH2VS36ykfevCZ1xwHSYS71tVHe2oA
0FhmQEkNapila60kQ7cBoY0399nUBOqd5HvPdqRE1f2NYOc75Mz11ZZhJOZfkUiqcHvql/xD7yDy
SKdPF98WuWtvMsGQCIYWDQh7LZUm26Yj7r9d5PQbK+G3FNtZ0xUlImqiU8k/B/xdxM6611ZGfQS5
Gl7h2fO0bG5s4jEo+x37wjI1DFExNiGH2vKpgZJFmmaf775mGeXOowkwNVBxhPI0OvQYGgRWH+ip
c2YljYtz09iENJEbyIWDJajw0S0stdcFXtE/UxdTq0volqZYAGkdx9hlCuJe05HPhAfFHpA97Lu4
Ok7Zx/HjEExkPcQ+D5b0Xz3PXG6b+KElNGfIDQX+WtQq1F5ouVlg+X6fSddcI8gJt8OZ2QPHB+NB
mEUDwZHs23JJ4tRjPGVlHL9KBK106nVTnBP8npLdEfWrTCd0M9VVbQVaUkQHDgAc2VAtZgb3apYn
j5rEpyKVvqQjJtrs3rHgcpcGAd6DSUuU/yy3u/nE7cwBTc0EYLcxMps/HYlaUnCjfgI7jF+mLaaf
kP2XO96OU0mutDThi0tzgyZaLMvkc3CM2aDzN9+8VkUbkbY3F6PSln+VKPqcfY/TTauZ0bEcZDa9
KZ+6HTa7AHP1hF5zbs6vRxCsxrNIyX7t2cXXaa7RUN4rgH+Evt6D1oVZ3XaflKN7abM3I0sMICiw
sBVNheALoI9TDwTj+QHtQX5wqACmMQV52cRi/tdB8L7S41HzPYhxGOUImaggdYhxj1JUH9zcLLJ8
eoDSv5kxA82Oo9SAUQjmSngaO58D84/m/AYQfKZI4Zx/A393NPfpoycMpBE9FAkc6pRfcbMVe+TP
2XlraRtY9U4H9tQlc8sfhrgF43d1vp4LtwuW8oSoB/d6JDSsb9epBGO+o7eLNAGI06RknkOHk08f
a+vDnBD/BYw5X4EG5++Q47uZ36wIVA56G7CaOveK1Hz+PT0gwkOdL/yR1LgQ4koDOwXLV7gdEYVx
4m2Y+LN5LpjrrF+7IFxJ3jaaJ4fG/kh2tqrv+ukYQl88/Wtsk0GaZHNgyKHjzKzgNk3a9emBiVag
h40Iqp6gMshX3w5rpBOMHtldh9EvBRdc7BKR/xmiL5jSiIP9jJH25X1Mb1jcSPtEgIQaXoKc+8vT
Ey4Rnxuder9n9uPbjrnSAVjK2YNLTI47biDyVBGvzZZRCI6DChft0xX19zGtu4wfnXRcBM4bk7zz
gxN4lFHCBmZkorewKUJ/kFjCTSW4Ofi3nBOEzfm+UR+9/rU4wbiv6MiLFjUCdgwsxESZqQVDaqZT
YxJXpL3VXsIlhUAx3hmY29DLv8FgECm5AKAGER4UMcteDxFh1FHH+zud9ITU
`protect end_protected
